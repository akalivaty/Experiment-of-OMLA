//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n208), .B2(KEYINPUT2), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT76), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT76), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT77), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(G148gat), .ZN(new_n216));
  INV_X1    g015(.A(G148gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT78), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G148gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n220), .A3(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT76), .B(G141gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n215), .B1(new_n223), .B2(G148gat), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT79), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n212), .A2(new_n214), .A3(G148gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT77), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT79), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n227), .A2(new_n228), .A3(new_n221), .A4(new_n216), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n210), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT2), .B1(new_n211), .B2(new_n217), .ZN(new_n232));
  AOI211_X1 g031(.A(new_n207), .B(new_n205), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(G113gat), .B(G120gat), .Z(new_n237));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n238));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  NOR3_X1   g040(.A1(new_n230), .A2(new_n233), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n202), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n229), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n209), .ZN(new_n246));
  INV_X1    g045(.A(new_n233), .ZN(new_n247));
  INV_X1    g046(.A(new_n241), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n246), .A2(new_n243), .A3(new_n247), .A4(new_n248), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n242), .A2(KEYINPUT82), .A3(new_n243), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n244), .A2(new_n250), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G225gat), .A2(G233gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n236), .A2(new_n240), .A3(KEYINPUT80), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT80), .B1(new_n236), .B2(new_n240), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n246), .A2(new_n247), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n263), .A3(new_n247), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n257), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n255), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n260), .B1(new_n246), .B2(new_n247), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n257), .B1(new_n267), .B2(new_n242), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n249), .A2(KEYINPUT4), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n251), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n265), .A2(new_n269), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT0), .ZN(new_n279));
  XNOR2_X1  g078(.A(G57gat), .B(G85gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n273), .A2(new_n274), .A3(new_n277), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(KEYINPUT6), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n274), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n271), .B1(new_n255), .B2(new_n265), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n275), .A2(new_n251), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n233), .B1(new_n245), .B2(new_n209), .ZN(new_n288));
  OAI22_X1  g087(.A1(new_n288), .A2(new_n263), .B1(new_n258), .B2(new_n259), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n230), .A2(KEYINPUT3), .A3(new_n233), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n256), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n287), .A2(new_n291), .A3(new_n270), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n284), .B(new_n285), .C1(new_n286), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT27), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G183gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT27), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT65), .B(new_n300), .C1(new_n296), .C2(G183gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n303), .B1(new_n302), .B2(new_n304), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n301), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(new_n304), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT66), .ZN(new_n309));
  INV_X1    g108(.A(new_n301), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT26), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n307), .A2(new_n312), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n314), .A2(KEYINPUT23), .ZN(new_n321));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT25), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT24), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT64), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n298), .A2(new_n300), .ZN(new_n332));
  NAND3_X1  g131(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n313), .A2(KEYINPUT64), .A3(new_n328), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n327), .A2(new_n335), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n329), .A2(new_n332), .A3(new_n333), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n326), .B1(new_n337), .B2(new_n325), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT29), .B1(new_n320), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G226gat), .A2(G233gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n295), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n320), .B2(new_n339), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n320), .A2(new_n339), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n344), .B1(new_n347), .B2(new_n341), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n343), .B1(new_n348), .B2(new_n295), .ZN(new_n349));
  INV_X1    g148(.A(G197gat), .ZN(new_n350));
  INV_X1    g149(.A(G204gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G197gat), .A2(G204gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT22), .ZN(new_n354));
  NAND2_X1  g153(.A1(G211gat), .A2(G218gat), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n352), .A2(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT70), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n356), .A2(new_n357), .ZN(new_n359));
  INV_X1    g158(.A(new_n355), .ZN(new_n360));
  NOR2_X1   g159(.A1(G211gat), .A2(G218gat), .ZN(new_n361));
  OAI22_X1  g160(.A1(new_n358), .A2(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n356), .A2(new_n357), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n360), .A2(new_n361), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n366), .A2(KEYINPUT71), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(KEYINPUT71), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n345), .A2(new_n342), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(new_n342), .B2(new_n340), .ZN(new_n372));
  INV_X1    g171(.A(new_n366), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G8gat), .B(G36gat), .Z(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT73), .ZN(new_n377));
  XOR2_X1   g176(.A(G64gat), .B(G92gat), .Z(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n370), .A2(KEYINPUT30), .A3(new_n375), .A4(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT74), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n374), .B1(new_n349), .B2(new_n369), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n384), .A2(KEYINPUT74), .A3(KEYINPUT30), .A4(new_n380), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(KEYINPUT75), .B(KEYINPUT30), .Z(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n384), .B2(new_n380), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n380), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n294), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n392));
  INV_X1    g191(.A(G22gat), .ZN(new_n393));
  INV_X1    g192(.A(G228gat), .ZN(new_n394));
  INV_X1    g193(.A(G233gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n366), .B1(new_n264), .B2(new_n346), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT29), .B1(new_n362), .B2(new_n365), .ZN(new_n399));
  OAI22_X1  g198(.A1(new_n399), .A2(KEYINPUT3), .B1(new_n230), .B2(new_n233), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n397), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT86), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT29), .B1(new_n288), .B2(new_n263), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n400), .B1(new_n405), .B2(new_n366), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(KEYINPUT86), .A3(new_n397), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n400), .A2(new_n396), .ZN(new_n409));
  INV_X1    g208(.A(new_n405), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n369), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n393), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  AOI211_X1 g212(.A(G22gat), .B(new_n411), .C1(new_n404), .C2(new_n407), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n392), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G78gat), .B(G106gat), .ZN(new_n416));
  INV_X1    g215(.A(G50gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  NAND2_X1  g219(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n373), .B1(new_n290), .B2(KEYINPUT29), .ZN(new_n422));
  AOI211_X1 g221(.A(new_n403), .B(new_n396), .C1(new_n422), .C2(new_n400), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT86), .B1(new_n406), .B2(new_n397), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n412), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G22gat), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n412), .B(new_n393), .C1(new_n423), .C2(new_n424), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n420), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n392), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G227gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(new_n395), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n320), .A2(new_n248), .A3(new_n339), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n248), .B1(new_n320), .B2(new_n339), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT32), .ZN(new_n436));
  XNOR2_X1  g235(.A(G15gat), .B(G43gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n436), .B1(KEYINPUT33), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT34), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n433), .A2(new_n434), .A3(new_n432), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT68), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n434), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n320), .A2(new_n248), .A3(new_n339), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(KEYINPUT68), .B(KEYINPUT34), .C1(new_n448), .C2(new_n432), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n441), .B1(new_n450), .B2(KEYINPUT69), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT33), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n439), .B1(new_n435), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n436), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT67), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(KEYINPUT67), .A3(new_n436), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n450), .A2(KEYINPUT69), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n451), .A3(new_n458), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n391), .A2(new_n421), .A3(new_n430), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT35), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n429), .B1(new_n428), .B2(new_n392), .ZN(new_n467));
  AOI211_X1 g266(.A(KEYINPUT85), .B(new_n420), .C1(new_n426), .C2(new_n427), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n391), .A4(new_n464), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT72), .B1(new_n347), .B2(new_n341), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n372), .B2(KEYINPUT72), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n367), .A2(new_n368), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n375), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n380), .B1(new_n477), .B2(KEYINPUT37), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT37), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT88), .B1(new_n384), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n340), .A2(new_n342), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT72), .B1(new_n481), .B2(new_n344), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n476), .B1(new_n482), .B2(new_n343), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n484));
  NOR4_X1   g283(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT37), .A4(new_n374), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n478), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT38), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n283), .A2(new_n293), .A3(new_n389), .ZN(new_n488));
  OAI22_X1  g287(.A1(new_n349), .A2(new_n369), .B1(new_n348), .B2(new_n366), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT37), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n380), .A2(KEYINPUT38), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n490), .B(new_n491), .C1(new_n480), .C2(new_n485), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n487), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n281), .B1(new_n273), .B2(new_n277), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n262), .A2(new_n264), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n256), .B1(new_n495), .B2(new_n276), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n249), .B(new_n256), .C1(new_n288), .C2(new_n260), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT39), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n497), .B2(KEYINPUT39), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n496), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT39), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n289), .A2(new_n290), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n502), .B(new_n257), .C1(new_n287), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n281), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT40), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n282), .B1(new_n496), .B2(new_n502), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n257), .B1(new_n287), .B2(new_n503), .ZN(new_n509));
  INV_X1    g308(.A(new_n500), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n507), .B(new_n508), .C1(new_n511), .C2(new_n499), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n494), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n386), .A2(new_n390), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n493), .A2(new_n515), .A3(new_n430), .A4(new_n421), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n294), .A2(new_n386), .A3(new_n390), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(new_n467), .B2(new_n468), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT36), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n460), .A2(new_n451), .A3(new_n458), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n460), .B1(new_n451), .B2(new_n458), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n462), .A2(KEYINPUT36), .A3(new_n463), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n472), .A2(new_n473), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n472), .A2(new_n525), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT89), .ZN(new_n528));
  XOR2_X1   g327(.A(G15gat), .B(G22gat), .Z(new_n529));
  INV_X1    g328(.A(G1gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT94), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT16), .B1(KEYINPUT92), .B2(G1gat), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(KEYINPUT92), .B2(G1gat), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n534), .A2(new_n529), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT95), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n536), .B1(new_n529), .B2(new_n530), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n537), .B2(KEYINPUT93), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n532), .B(new_n538), .C1(KEYINPUT93), .C2(new_n535), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G8gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(KEYINPUT95), .A2(G8gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n535), .A2(new_n531), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(G29gat), .A2(G36gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n417), .A2(G43gat), .ZN(new_n547));
  INV_X1    g346(.A(G43gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G50gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n549), .A3(KEYINPUT15), .ZN(new_n550));
  INV_X1    g349(.A(G29gat), .ZN(new_n551));
  INV_X1    g350(.A(G36gat), .ZN(new_n552));
  OR3_X1    g351(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT91), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT91), .B1(new_n551), .B2(new_n552), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n546), .A2(new_n550), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT90), .B1(new_n548), .B2(G50gat), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(G43gat), .B2(new_n417), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n548), .A2(KEYINPUT90), .A3(G50gat), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT15), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n546), .B1(new_n551), .B2(new_n552), .ZN(new_n561));
  INV_X1    g360(.A(new_n550), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n543), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT98), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n540), .A2(new_n563), .A3(new_n560), .A4(new_n542), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT97), .B(KEYINPUT13), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n569), .B(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n543), .A2(KEYINPUT98), .A3(new_n564), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT99), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n540), .A2(new_n542), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n564), .B(KEYINPUT17), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n565), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT18), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n581), .A2(KEYINPUT96), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n580), .A2(new_n571), .A3(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n579), .A2(new_n565), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(KEYINPUT96), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n570), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n583), .B1(new_n586), .B2(new_n582), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n576), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(G197gat), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT11), .B(G169gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT12), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT100), .ZN(new_n595));
  INV_X1    g394(.A(new_n593), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n576), .A2(new_n587), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n588), .A2(KEYINPUT100), .A3(new_n593), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT105), .B(KEYINPUT7), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(G85gat), .A3(G92gat), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G99gat), .A2(G106gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n608), .B1(new_n605), .B2(new_n606), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n604), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G99gat), .B(G106gat), .Z(new_n611));
  OR2_X1    g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n578), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n614), .ZN(new_n616));
  AND2_X1   g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n616), .A2(new_n564), .B1(KEYINPUT41), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT103), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT106), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  OR3_X1    g429(.A1(new_n619), .A2(new_n629), .A3(new_n620), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n622), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n626), .B(KEYINPUT104), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n628), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G57gat), .B(G64gat), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G71gat), .B(G78gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT21), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(G127gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n540), .B(new_n542), .C1(new_n641), .C2(new_n640), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n647), .A2(KEYINPUT101), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(KEYINPUT101), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n644), .B(G127gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G183gat), .B(G211gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT102), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n203), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n656), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n650), .A2(new_n653), .A3(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n616), .A2(new_n639), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT10), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n614), .A2(new_n640), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n616), .A2(KEYINPUT10), .A3(new_n639), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n667), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n670), .B1(new_n671), .B2(new_n664), .ZN(new_n672));
  XNOR2_X1  g471(.A(G120gat), .B(G148gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(G176gat), .B(G204gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n673), .B(new_n674), .Z(new_n675));
  AND2_X1   g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n672), .A2(new_n675), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n634), .A2(new_n663), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  AND4_X1   g479(.A1(new_n526), .A2(new_n528), .A3(new_n601), .A4(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n681), .A2(KEYINPUT107), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(KEYINPUT107), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n294), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g486(.A(KEYINPUT16), .B(G8gat), .Z(new_n688));
  NAND4_X1  g487(.A1(new_n684), .A2(KEYINPUT42), .A3(new_n514), .A4(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n514), .B1(new_n682), .B2(new_n683), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g491(.A(KEYINPUT108), .B(new_n514), .C1(new_n682), .C2(new_n683), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(G8gat), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n688), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n692), .B2(new_n693), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n689), .B(new_n694), .C1(new_n696), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g496(.A(G15gat), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n684), .A2(new_n698), .A3(new_n464), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n522), .A2(new_n523), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n684), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n701), .B2(new_n698), .ZN(G1326gat));
  NAND2_X1  g501(.A1(new_n421), .A2(new_n430), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n684), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  AND3_X1   g505(.A1(new_n528), .A2(new_n526), .A3(new_n601), .ZN(new_n707));
  INV_X1    g506(.A(new_n663), .ZN(new_n708));
  INV_X1    g507(.A(new_n634), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n709), .A3(new_n678), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n707), .A2(new_n551), .A3(new_n685), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n516), .A2(new_n714), .A3(new_n518), .A4(new_n524), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n472), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n700), .B1(new_n703), .B2(new_n517), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n714), .B1(new_n717), .B2(new_n516), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n709), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n634), .A2(new_n720), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n528), .A2(new_n526), .A3(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n678), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n600), .A2(new_n663), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G29gat), .B1(new_n727), .B2(new_n294), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n728), .ZN(G1328gat));
  NAND3_X1  g528(.A1(new_n724), .A2(new_n514), .A3(new_n726), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n730), .A2(G36gat), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n707), .A2(new_n552), .A3(new_n514), .A4(new_n711), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT46), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT110), .ZN(G1329gat));
  OAI21_X1  g534(.A(G43gat), .B1(new_n727), .B2(new_n524), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n707), .A2(new_n548), .A3(new_n464), .A4(new_n711), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT47), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n738), .B(new_n740), .ZN(G1330gat));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n724), .A2(new_n703), .A3(new_n726), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(G50gat), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n703), .A2(new_n417), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n711), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n745), .B2(new_n746), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n707), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n742), .B1(new_n744), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n417), .B1(new_n743), .B2(KEYINPUT113), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n724), .A2(new_n752), .A3(new_n703), .A4(new_n726), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n749), .A2(new_n742), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT114), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758));
  AOI211_X1 g557(.A(new_n758), .B(new_n755), .C1(new_n751), .C2(new_n753), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n750), .B1(new_n757), .B2(new_n759), .ZN(G1331gat));
  OR2_X1    g559(.A1(new_n716), .A2(new_n718), .ZN(new_n761));
  NOR4_X1   g560(.A1(new_n601), .A2(new_n708), .A3(new_n709), .A4(new_n678), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n685), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n514), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT49), .B(G64gat), .Z(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n763), .B2(new_n524), .ZN(new_n771));
  INV_X1    g570(.A(G71gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n464), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n763), .B2(new_n773), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g574(.A1(new_n764), .A2(new_n703), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n601), .B2(new_n663), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n600), .A2(KEYINPUT115), .A3(new_n708), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n678), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n721), .A2(new_n723), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n721), .A2(new_n723), .A3(KEYINPUT116), .A4(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786), .B2(new_n294), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n779), .A2(new_n780), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT51), .B1(new_n789), .B2(new_n719), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n761), .A2(new_n791), .A3(new_n709), .A4(new_n788), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n790), .A2(new_n792), .A3(new_n725), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(new_n605), .A3(new_n685), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n787), .A2(new_n794), .ZN(G1336gat));
  INV_X1    g594(.A(new_n514), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(G92gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  OAI21_X1  g598(.A(G92gat), .B1(new_n782), .B2(new_n796), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n798), .A2(KEYINPUT118), .A3(new_n799), .A4(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n784), .A2(new_n514), .A3(new_n785), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G92gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n798), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n806), .B1(new_n809), .B2(KEYINPUT52), .ZN(new_n810));
  AND4_X1   g609(.A1(new_n725), .A2(new_n790), .A3(new_n792), .A4(new_n797), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n807), .B2(G92gat), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n812), .A2(KEYINPUT117), .A3(new_n799), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n805), .B1(new_n810), .B2(new_n813), .ZN(G1337gat));
  INV_X1    g613(.A(G99gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n786), .A2(new_n815), .A3(new_n524), .ZN(new_n816));
  AOI21_X1  g615(.A(G99gat), .B1(new_n793), .B2(new_n464), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(G1338gat));
  INV_X1    g617(.A(G106gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n793), .A2(new_n819), .A3(new_n703), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  OAI21_X1  g620(.A(G106gat), .B1(new_n782), .B2(new_n469), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G106gat), .B1(new_n786), .B2(new_n469), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n820), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n825), .B2(new_n821), .ZN(G1339gat));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n670), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n668), .A2(new_n669), .A3(new_n664), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n675), .B1(new_n670), .B2(new_n827), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT55), .B1(new_n830), .B2(new_n831), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n832), .A2(new_n833), .A3(new_n676), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n598), .A2(new_n599), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n584), .A2(new_n570), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n572), .B1(new_n568), .B2(new_n573), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n592), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n725), .A2(new_n597), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n709), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  AND4_X1   g639(.A1(new_n597), .A2(new_n709), .A3(new_n834), .A4(new_n838), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n708), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n600), .A2(new_n680), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n703), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n844), .A2(new_n685), .A3(new_n796), .A4(new_n464), .ZN(new_n845));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n600), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n294), .B1(new_n842), .B2(new_n843), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n469), .A2(new_n464), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n796), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT119), .Z(new_n851));
  NOR2_X1   g650(.A1(new_n600), .A2(G113gat), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n852), .B(KEYINPUT120), .Z(new_n853));
  OAI21_X1  g652(.A(new_n846), .B1(new_n851), .B2(new_n853), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n845), .B2(new_n678), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n678), .A2(G120gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n851), .B2(new_n856), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n845), .B2(new_n708), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n663), .A2(new_n645), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n850), .B2(new_n859), .ZN(G1342gat));
  NOR3_X1   g659(.A1(new_n634), .A2(G134gat), .A3(new_n514), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n849), .A2(new_n861), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n863));
  OAI21_X1  g662(.A(G134gat), .B1(new_n845), .B2(new_n634), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(G1343gat));
  INV_X1    g665(.A(new_n223), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n700), .A2(new_n294), .A3(new_n514), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n842), .A2(new_n843), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n869), .A2(KEYINPUT57), .A3(new_n703), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n869), .B2(new_n703), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n867), .B1(new_n872), .B2(new_n600), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n847), .A2(new_n703), .A3(new_n524), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n514), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n211), .A3(new_n601), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT58), .ZN(G1344gat));
  AND2_X1   g677(.A1(new_n218), .A2(new_n220), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n875), .A2(new_n879), .A3(new_n725), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n600), .A2(KEYINPUT121), .A3(new_n680), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT121), .B1(new_n600), .B2(new_n680), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n842), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n469), .B1(new_n885), .B2(KEYINPUT122), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n842), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n725), .B(new_n868), .C1(new_n889), .C2(new_n870), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n881), .B1(new_n890), .B2(G148gat), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n725), .B(new_n868), .C1(new_n870), .C2(new_n871), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(KEYINPUT59), .A3(new_n879), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n880), .B1(new_n891), .B2(new_n894), .ZN(G1345gat));
  OAI21_X1  g694(.A(G155gat), .B1(new_n872), .B2(new_n708), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n875), .A2(new_n203), .A3(new_n663), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n872), .B2(new_n634), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n709), .A2(new_n204), .A3(new_n796), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n874), .B2(new_n900), .ZN(G1347gat));
  NAND3_X1  g700(.A1(new_n464), .A2(new_n294), .A3(new_n514), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n902), .B(KEYINPUT123), .Z(new_n903));
  NAND2_X1  g702(.A1(new_n844), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(G169gat), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n904), .A2(new_n905), .A3(new_n600), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n685), .B1(new_n842), .B2(new_n843), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n907), .A2(new_n514), .A3(new_n848), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n601), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n906), .B1(new_n909), .B2(new_n905), .ZN(G1348gat));
  INV_X1    g709(.A(G176gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(new_n911), .A3(new_n725), .ZN(new_n912));
  OAI21_X1  g711(.A(G176gat), .B1(new_n904), .B2(new_n678), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1349gat));
  NAND4_X1  g713(.A1(new_n908), .A2(new_n297), .A3(new_n299), .A4(new_n663), .ZN(new_n915));
  OAI21_X1  g714(.A(G183gat), .B1(new_n904), .B2(new_n708), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n908), .A2(new_n300), .A3(new_n709), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n844), .A2(new_n709), .A3(new_n903), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n920), .A2(new_n921), .A3(G190gat), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n920), .B2(G190gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT124), .Z(G1351gat));
  NOR3_X1   g724(.A1(new_n700), .A2(new_n685), .A3(new_n796), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n889), .B2(new_n870), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(new_n350), .A3(new_n600), .ZN(new_n928));
  AND4_X1   g727(.A1(new_n514), .A2(new_n907), .A3(new_n703), .A4(new_n524), .ZN(new_n929));
  AOI21_X1  g728(.A(G197gat), .B1(new_n929), .B2(new_n601), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n928), .A2(new_n930), .ZN(G1352gat));
  OAI21_X1  g730(.A(G204gat), .B1(new_n927), .B2(new_n678), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n929), .A2(new_n351), .A3(new_n725), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(KEYINPUT125), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n932), .B(new_n935), .C1(new_n933), .C2(new_n936), .ZN(G1353gat));
  OAI211_X1 g736(.A(new_n663), .B(new_n926), .C1(new_n889), .C2(new_n870), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT63), .B1(new_n938), .B2(G211gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(G211gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n929), .A2(new_n942), .A3(new_n663), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT126), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n938), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT127), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n941), .B(new_n944), .C1(new_n946), .C2(new_n939), .ZN(G1354gat));
  OAI21_X1  g746(.A(G218gat), .B1(new_n927), .B2(new_n634), .ZN(new_n948));
  INV_X1    g747(.A(G218gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n929), .A2(new_n949), .A3(new_n709), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1355gat));
endmodule


