//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  INV_X1    g000(.A(G230gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT99), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT7), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n205), .B(KEYINPUT99), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT7), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212));
  INV_X1    g011(.A(G85gat), .ZN(new_n213));
  INV_X1    g012(.A(G92gat), .ZN(new_n214));
  AOI22_X1  g013(.A1(KEYINPUT8), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n208), .A2(new_n211), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G99gat), .B(G106gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n208), .A2(new_n211), .A3(new_n217), .A4(new_n215), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G71gat), .A2(G78gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(G57gat), .B(G64gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT9), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(G71gat), .A2(G78gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT97), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(KEYINPUT9), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n223), .B1(new_n222), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n221), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT10), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n220), .A3(new_n231), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n235), .A2(new_n234), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n204), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n204), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(new_n233), .B2(new_n235), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G120gat), .B(G148gat), .ZN(new_n242));
  INV_X1    g041(.A(G176gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G204gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n241), .B(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G29gat), .ZN(new_n249));
  INV_X1    g048(.A(G36gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT14), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT14), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(G29gat), .B2(G36gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(G29gat), .A2(G36gat), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT93), .ZN(new_n256));
  INV_X1    g055(.A(G43gat), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT15), .B1(new_n257), .B2(G50gat), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n257), .B2(G50gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n256), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT94), .B(G50gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n257), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(new_n257), .B2(G50gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT15), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n255), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT17), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT17), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n260), .A2(new_n269), .A3(new_n266), .ZN(new_n270));
  XNOR2_X1  g069(.A(G15gat), .B(G22gat), .ZN(new_n271));
  INV_X1    g070(.A(G1gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(KEYINPUT16), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G8gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT95), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n273), .B(new_n275), .C1(new_n272), .C2(new_n271), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n274), .A2(KEYINPUT95), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n268), .A2(new_n270), .A3(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n267), .A2(new_n278), .ZN(new_n280));
  NAND2_X1  g079(.A1(G229gat), .A2(G233gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT18), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n267), .B(new_n278), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n281), .B(KEYINPUT96), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT13), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT18), .A4(new_n281), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT11), .B(G169gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(G197gat), .ZN(new_n292));
  XOR2_X1   g091(.A(G113gat), .B(G141gat), .Z(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT12), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n284), .A2(new_n295), .A3(new_n288), .A4(new_n289), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G228gat), .A2(G233gat), .ZN(new_n301));
  INV_X1    g100(.A(G148gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G141gat), .ZN(new_n303));
  INV_X1    g102(.A(G141gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G148gat), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT2), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT73), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n309), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(new_n307), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n314));
  XNOR2_X1  g113(.A(G141gat), .B(G148gat), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n313), .B(new_n314), .C1(new_n315), .C2(KEYINPUT2), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n305), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n304), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n303), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n309), .B1(new_n308), .B2(KEYINPUT2), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n311), .A2(new_n316), .B1(new_n322), .B2(new_n321), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT75), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G197gat), .B(G204gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT22), .ZN(new_n331));
  NAND2_X1  g130(.A1(G211gat), .A2(G218gat), .ZN(new_n332));
  INV_X1    g131(.A(G211gat), .ZN(new_n333));
  INV_X1    g132(.A(G218gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT22), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n332), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(KEYINPUT70), .A3(new_n330), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT70), .B1(new_n338), .B2(new_n330), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n336), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n341), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n335), .A2(new_n332), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n348), .A2(new_n339), .B1(new_n331), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n351), .B2(KEYINPUT29), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n301), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n327), .B1(new_n344), .B2(new_n345), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n327), .A2(new_n345), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n342), .B1(new_n355), .B2(new_n343), .ZN(new_n356));
  INV_X1    g155(.A(new_n301), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(G22gat), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n346), .A2(new_n324), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(new_n301), .A3(new_n352), .ZN(new_n361));
  INV_X1    g160(.A(G22gat), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n356), .B1(new_n329), .B2(new_n346), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n361), .B(new_n362), .C1(new_n363), .C2(new_n301), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n359), .A2(new_n364), .A3(KEYINPUT81), .ZN(new_n365));
  XNOR2_X1  g164(.A(G78gat), .B(G106gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT31), .B(G50gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n359), .A2(new_n364), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n371), .B2(new_n372), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n369), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n371), .A2(new_n372), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT82), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n379), .A2(new_n365), .A3(new_n368), .A4(new_n374), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT85), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(KEYINPUT40), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  AOI221_X4 g186(.A(new_n325), .B1(new_n321), .B2(new_n322), .C1(new_n311), .C2(new_n316), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT75), .B1(new_n317), .B2(new_n323), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT3), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT76), .ZN(new_n391));
  INV_X1    g190(.A(G134gat), .ZN(new_n392));
  INV_X1    g191(.A(G127gat), .ZN(new_n393));
  INV_X1    g192(.A(G120gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G113gat), .ZN(new_n395));
  INV_X1    g194(.A(G113gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G120gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT1), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n393), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI211_X1 g199(.A(KEYINPUT1), .B(G127gat), .C1(new_n395), .C2(new_n397), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n392), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G113gat), .B(G120gat), .ZN(new_n403));
  OAI21_X1  g202(.A(G127gat), .B1(new_n403), .B2(KEYINPUT1), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n396), .A2(G120gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n394), .A2(G113gat), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n399), .B(new_n393), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(G134gat), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT76), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n410), .B(KEYINPUT3), .C1(new_n388), .C2(new_n389), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n391), .A2(new_n409), .A3(new_n411), .A4(new_n355), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n404), .A2(G134gat), .A3(new_n407), .ZN(new_n413));
  AOI21_X1  g212(.A(G134gat), .B1(new_n404), .B2(new_n407), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT68), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT68), .B1(new_n402), .B2(new_n408), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n418), .A2(KEYINPUT78), .A3(new_n419), .A4(new_n327), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n415), .B1(new_n413), .B2(new_n414), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n402), .A2(KEYINPUT68), .A3(new_n408), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n421), .A2(new_n422), .A3(new_n419), .A4(new_n327), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n413), .A2(new_n414), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n419), .B1(new_n424), .B2(new_n327), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n387), .B1(new_n412), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT39), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n409), .B1(new_n388), .B2(new_n389), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT77), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n424), .A2(new_n327), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT77), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(new_n409), .C1(new_n388), .C2(new_n389), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n387), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n429), .A2(new_n430), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT0), .B(G57gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G85gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(G1gat), .B(G29gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  AOI211_X1 g244(.A(KEYINPUT84), .B(new_n445), .C1(new_n429), .C2(new_n430), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n412), .A2(new_n428), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(new_n430), .A3(new_n437), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n449), .B2(new_n444), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n386), .B(new_n440), .C1(new_n446), .C2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G64gat), .B(G92gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(G36gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(KEYINPUT72), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(G8gat), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT71), .ZN(new_n456));
  NAND2_X1  g255(.A1(G183gat), .A2(G190gat), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(G169gat), .A2(G176gat), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(KEYINPUT26), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G169gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(new_n243), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n459), .A2(KEYINPUT26), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT27), .B(G183gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(KEYINPUT66), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT27), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G183gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT66), .ZN(new_n469));
  INV_X1    g268(.A(G190gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT67), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT28), .ZN(new_n473));
  AOI21_X1  g272(.A(G190gat), .B1(new_n468), .B2(KEYINPUT66), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT67), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n474), .B(new_n475), .C1(KEYINPUT66), .C2(new_n465), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n465), .A2(KEYINPUT28), .A3(new_n470), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n464), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(KEYINPUT64), .ZN(new_n481));
  NOR2_X1   g280(.A1(G183gat), .A2(G190gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT24), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(new_n457), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT25), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n462), .B1(KEYINPUT23), .B2(new_n459), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT65), .B1(new_n459), .B2(KEYINPUT23), .ZN(new_n489));
  OR3_X1    g288(.A1(new_n459), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n485), .A2(new_n480), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT25), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n343), .B1(new_n479), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G226gat), .A2(G233gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(G226gat), .B(G233gat), .C1(new_n479), .C2(new_n496), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n456), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT71), .B1(new_n497), .B2(new_n498), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n350), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n499), .A2(new_n500), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n342), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n455), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n503), .A2(new_n505), .A3(new_n455), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(KEYINPUT30), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n503), .A2(new_n505), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(new_n455), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n451), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT86), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT5), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n436), .B2(new_n437), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n437), .B1(new_n433), .B2(new_n419), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n418), .A2(KEYINPUT4), .A3(new_n327), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n345), .B1(new_n326), .B2(new_n328), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n355), .B1(new_n520), .B2(new_n410), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n411), .A2(new_n409), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n518), .B(new_n519), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n424), .B1(new_n520), .B2(new_n410), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n351), .B1(new_n390), .B2(KEYINPUT76), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n524), .A2(new_n525), .B1(new_n420), .B2(new_n427), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n437), .A2(KEYINPUT5), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n517), .A2(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n515), .B1(new_n528), .B2(new_n444), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n517), .A2(new_n523), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n526), .A2(new_n527), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(KEYINPUT86), .A3(new_n445), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  AOI211_X1 g333(.A(KEYINPUT39), .B(new_n387), .C1(new_n412), .C2(new_n428), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT84), .B1(new_n535), .B2(new_n445), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n449), .A2(new_n447), .A3(new_n444), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n439), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n534), .B1(new_n538), .B2(new_n386), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n383), .B1(new_n514), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n440), .B1(new_n446), .B2(new_n450), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n541), .A2(new_n385), .B1(new_n529), .B2(new_n533), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n503), .A2(new_n505), .A3(new_n455), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n543), .A2(new_n506), .A3(new_n512), .ZN(new_n544));
  INV_X1    g343(.A(new_n455), .ZN(new_n545));
  NOR3_X1   g344(.A1(new_n510), .A2(KEYINPUT30), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n542), .A2(KEYINPUT87), .A3(new_n547), .A4(new_n451), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n382), .B1(new_n540), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT6), .B1(new_n528), .B2(new_n444), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT86), .B1(new_n532), .B2(new_n445), .ZN(new_n552));
  AOI211_X1 g351(.A(new_n515), .B(new_n444), .C1(new_n530), .C2(new_n531), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n550), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n550), .B1(new_n534), .B2(new_n551), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n504), .A2(new_n342), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT89), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n501), .A2(new_n502), .A3(new_n350), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT37), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT37), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n455), .B1(new_n511), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT38), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n528), .A2(new_n444), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT6), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n563), .B1(new_n562), .B2(new_n511), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n543), .B1(new_n568), .B2(KEYINPUT38), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n557), .A2(new_n565), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n549), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT90), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n509), .A2(new_n513), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT6), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(new_n532), .B2(new_n445), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n567), .B1(new_n566), .B2(new_n576), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n574), .A2(new_n577), .A3(KEYINPUT79), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT79), .B1(new_n574), .B2(new_n577), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n377), .A2(new_n380), .A3(KEYINPUT83), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT83), .B1(new_n377), .B2(new_n380), .ZN(new_n581));
  OAI22_X1  g380(.A1(new_n578), .A2(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(G227gat), .A2(G233gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n477), .A2(new_n478), .ZN(new_n585));
  INV_X1    g384(.A(new_n464), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n496), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n418), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OAI22_X1  g388(.A1(new_n479), .A2(new_n496), .B1(new_n416), .B2(new_n417), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n584), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT32), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n591), .B1(new_n592), .B2(KEYINPUT33), .ZN(new_n593));
  XNOR2_X1  g392(.A(G15gat), .B(G43gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G71gat), .ZN(new_n595));
  INV_X1    g394(.A(G99gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT33), .B1(new_n597), .B2(KEYINPUT69), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n601), .B1(KEYINPUT69), .B2(new_n597), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n591), .A2(new_n592), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n589), .A2(new_n584), .A3(new_n590), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n605), .B(KEYINPUT34), .Z(new_n606));
  AND3_X1   g405(.A1(new_n600), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n600), .B2(new_n604), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT36), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n582), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n549), .A2(KEYINPUT90), .A3(new_n570), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n573), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n534), .A2(new_n551), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT88), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(new_n567), .A3(new_n554), .ZN(new_n618));
  AND4_X1   g417(.A1(new_n615), .A2(new_n618), .A3(new_n574), .A4(new_n381), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n609), .B(KEYINPUT91), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n381), .A2(new_n609), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n574), .A2(new_n577), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT79), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n574), .A2(new_n577), .A3(KEYINPUT79), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n628), .A2(KEYINPUT92), .A3(KEYINPUT35), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT92), .B1(new_n628), .B2(KEYINPUT35), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n621), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI211_X1 g430(.A(new_n248), .B(new_n300), .C1(new_n614), .C2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT21), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n278), .B1(new_n633), .B2(new_n232), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT98), .ZN(new_n635));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n231), .A2(KEYINPUT21), .ZN(new_n638));
  XNOR2_X1  g437(.A(G127gat), .B(G155gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n642));
  XNOR2_X1  g441(.A(G183gat), .B(G211gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n637), .A2(new_n640), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n637), .A2(new_n640), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n268), .A2(new_n221), .A3(new_n270), .ZN(new_n652));
  NAND3_X1  g451(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n652), .B(new_n653), .C1(new_n221), .C2(new_n267), .ZN(new_n654));
  XOR2_X1   g453(.A(G190gat), .B(G218gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n657));
  INV_X1    g456(.A(new_n655), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n657), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G134gat), .B(G162gat), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n654), .B(new_n658), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n659), .A2(new_n662), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n632), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n577), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(new_n272), .ZN(G1324gat));
  INV_X1    g470(.A(new_n669), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(new_n547), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n674), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  AOI211_X1 g478(.A(KEYINPUT102), .B(new_n274), .C1(new_n672), .C2(new_n547), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n672), .A2(new_n547), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(G8gat), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n677), .B(new_n679), .C1(new_n680), .C2(new_n683), .ZN(G1325gat));
  INV_X1    g483(.A(new_n610), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n672), .A2(G15gat), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(G15gat), .B1(new_n672), .B2(new_n620), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n687), .A2(KEYINPUT103), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(KEYINPUT103), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n580), .A2(new_n581), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n669), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(new_n362), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n692), .B(new_n694), .ZN(G1327gat));
  INV_X1    g494(.A(new_n667), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n614), .B2(new_n631), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n650), .A2(new_n248), .A3(new_n300), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n577), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n249), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT45), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n549), .A2(KEYINPUT90), .A3(new_n570), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT90), .B1(new_n549), .B2(new_n570), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n703), .A2(new_n704), .A3(new_n611), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT92), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n578), .A2(new_n579), .A3(new_n622), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(new_n615), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n628), .A2(KEYINPUT92), .A3(KEYINPUT35), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n708), .A2(new_n709), .B1(new_n620), .B2(new_n619), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n667), .B1(new_n705), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n614), .A2(new_n631), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(KEYINPUT44), .A3(new_n667), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n698), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n577), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n718), .ZN(G1328gat));
  NAND3_X1  g518(.A1(new_n699), .A2(new_n250), .A3(new_n547), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT46), .Z(new_n721));
  OAI21_X1  g520(.A(G36gat), .B1(new_n717), .B2(new_n574), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1329gat));
  NAND2_X1  g522(.A1(new_n699), .A2(new_n620), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n257), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n685), .A2(G43gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n717), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT47), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n729), .B(new_n725), .C1(new_n717), .C2(new_n726), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1330gat));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n382), .A3(new_n698), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n262), .ZN(new_n733));
  INV_X1    g532(.A(new_n691), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n699), .A2(new_n261), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(KEYINPUT48), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n735), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n716), .A2(new_n734), .A3(new_n698), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(new_n262), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n736), .B1(KEYINPUT48), .B2(new_n739), .ZN(G1331gat));
  NAND2_X1  g539(.A1(new_n668), .A2(new_n300), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n614), .B2(new_n631), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n742), .A2(new_n248), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n577), .B(KEYINPUT105), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n742), .A2(new_n248), .A3(new_n547), .A4(new_n747), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n748), .A2(KEYINPUT106), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(KEYINPUT106), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n751), .B(new_n752), .Z(G1333gat));
  NAND2_X1  g552(.A1(new_n743), .A2(new_n620), .ZN(new_n754));
  INV_X1    g553(.A(G71gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n743), .A2(G71gat), .A3(new_n685), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n734), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g560(.A1(new_n650), .A2(new_n299), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n667), .B(new_n762), .C1(new_n705), .C2(new_n710), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT51), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n697), .A2(new_n765), .A3(new_n762), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n764), .A2(new_n766), .A3(new_n248), .ZN(new_n767));
  AOI21_X1  g566(.A(G85gat), .B1(new_n767), .B2(new_n700), .ZN(new_n768));
  INV_X1    g567(.A(new_n248), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n650), .A2(new_n769), .A3(new_n299), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n716), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n213), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n768), .B1(new_n772), .B2(new_n700), .ZN(G1336gat));
  NOR2_X1   g572(.A1(new_n574), .A2(G92gat), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n764), .A2(new_n766), .A3(new_n248), .A4(new_n774), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n775), .A2(KEYINPUT108), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n713), .A2(new_n547), .A3(new_n715), .A4(new_n770), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G92gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n775), .A2(KEYINPUT108), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n776), .A2(new_n777), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n778), .A2(new_n782), .A3(G92gat), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n778), .B2(G92gat), .ZN(new_n784));
  INV_X1    g583(.A(new_n775), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n781), .B1(new_n786), .B2(new_n777), .ZN(G1337gat));
  OAI21_X1  g586(.A(G99gat), .B1(new_n771), .B2(new_n610), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n767), .A2(new_n596), .A3(new_n620), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1338gat));
  NAND4_X1  g589(.A1(new_n713), .A2(new_n734), .A3(new_n715), .A4(new_n770), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G106gat), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n381), .A2(G106gat), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n764), .A2(new_n766), .A3(new_n248), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT53), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n713), .A2(new_n382), .A3(new_n715), .A4(new_n770), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G106gat), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n797), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  AND4_X1   g601(.A1(new_n797), .A2(new_n801), .A3(new_n798), .A4(new_n794), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n796), .B1(new_n802), .B2(new_n803), .ZN(G1339gat));
  NAND2_X1  g603(.A1(new_n236), .A2(new_n237), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n239), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n236), .A2(new_n237), .A3(new_n204), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(KEYINPUT54), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n247), .B1(new_n238), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n810), .A3(KEYINPUT55), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n241), .A2(new_n247), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT110), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT110), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n811), .A2(new_n815), .A3(new_n812), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n808), .A2(new_n810), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n814), .A2(new_n299), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n285), .A2(new_n287), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n281), .B1(new_n279), .B2(new_n280), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n294), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n298), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n248), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n820), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n696), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n813), .A2(KEYINPUT110), .B1(new_n818), .B2(new_n817), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n828), .A2(new_n667), .A3(new_n824), .A4(new_n816), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(KEYINPUT111), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n667), .B1(new_n820), .B2(new_n825), .ZN(new_n832));
  AND4_X1   g631(.A1(new_n667), .A2(new_n828), .A3(new_n824), .A4(new_n816), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n830), .A2(new_n834), .A3(new_n651), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n650), .A2(new_n696), .A3(new_n769), .A4(new_n300), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(KEYINPUT112), .A3(new_n836), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n839), .A2(new_n744), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n574), .A3(new_n623), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n396), .A3(new_n299), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n620), .A2(new_n691), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n839), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n547), .A2(new_n577), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G113gat), .B1(new_n848), .B2(new_n300), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT113), .Z(G1340gat));
  NAND3_X1  g650(.A1(new_n843), .A2(new_n394), .A3(new_n248), .ZN(new_n852));
  OAI21_X1  g651(.A(G120gat), .B1(new_n848), .B2(new_n769), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1341gat));
  NOR3_X1   g653(.A1(new_n848), .A2(new_n393), .A3(new_n651), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n842), .A2(KEYINPUT114), .A3(new_n651), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT114), .B1(new_n842), .B2(new_n651), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n855), .B1(new_n858), .B2(new_n393), .ZN(G1342gat));
  NAND2_X1  g658(.A1(new_n574), .A2(new_n667), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT115), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AND4_X1   g661(.A1(new_n392), .A2(new_n841), .A3(new_n623), .A4(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n864));
  OR3_X1    g663(.A1(new_n863), .A2(KEYINPUT116), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n848), .B2(new_n696), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT116), .B1(new_n863), .B2(new_n864), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n868), .ZN(G1343gat));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n610), .A2(new_n847), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n839), .A2(new_n382), .A3(new_n840), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n836), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n299), .A2(new_n819), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n825), .B1(new_n876), .B2(new_n813), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n696), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n650), .B1(new_n878), .B2(new_n829), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n734), .B(KEYINPUT57), .C1(new_n875), .C2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AOI211_X1 g682(.A(new_n300), .B(new_n871), .C1(new_n874), .C2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n870), .B1(new_n884), .B2(new_n304), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n871), .B1(new_n874), .B2(new_n883), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n299), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(KEYINPUT118), .A3(G141gat), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n685), .A2(new_n381), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n841), .A2(new_n574), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n304), .A3(new_n299), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n885), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT58), .ZN(new_n893));
  XNOR2_X1  g692(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n891), .B(new_n894), .C1(new_n884), .C2(new_n304), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(G1344gat));
  AOI21_X1  g695(.A(KEYINPUT59), .B1(new_n886), .B2(new_n248), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n878), .A2(new_n829), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n836), .B1(new_n898), .B2(new_n650), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n734), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n873), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n903), .B1(new_n872), .B2(new_n873), .ZN(new_n904));
  INV_X1    g703(.A(new_n871), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n248), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G148gat), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n897), .A2(G148gat), .B1(new_n907), .B2(KEYINPUT59), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n890), .A2(KEYINPUT120), .A3(new_n302), .A4(new_n248), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n841), .A2(new_n302), .A3(new_n574), .A4(new_n889), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n769), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT122), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n907), .A2(KEYINPUT59), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n886), .A2(new_n248), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n917), .A3(G148gat), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n909), .A2(new_n912), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n914), .A2(new_n922), .ZN(G1345gat));
  AOI21_X1  g722(.A(G155gat), .B1(new_n890), .B2(new_n650), .ZN(new_n924));
  INV_X1    g723(.A(new_n886), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(new_n651), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n924), .B1(new_n926), .B2(G155gat), .ZN(G1346gat));
  OAI21_X1  g726(.A(G162gat), .B1(new_n925), .B2(new_n696), .ZN(new_n928));
  INV_X1    g727(.A(G162gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n841), .A2(new_n929), .A3(new_n889), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n928), .B1(new_n861), .B2(new_n930), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n744), .A2(new_n574), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n839), .A2(new_n840), .A3(new_n845), .A4(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G169gat), .B1(new_n933), .B2(new_n300), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n839), .A2(new_n577), .A3(new_n840), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n622), .A2(new_n574), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(new_n461), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n937), .B2(new_n300), .ZN(G1348gat));
  NOR3_X1   g737(.A1(new_n933), .A2(new_n243), .A3(new_n769), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n935), .A2(new_n248), .A3(new_n936), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n243), .B2(new_n940), .ZN(G1349gat));
  NAND4_X1  g740(.A1(new_n935), .A2(new_n650), .A3(new_n465), .A4(new_n936), .ZN(new_n942));
  OAI21_X1  g741(.A(G183gat), .B1(new_n933), .B2(new_n651), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT124), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT60), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n945), .B(new_n947), .ZN(G1350gat));
  OAI21_X1  g747(.A(G190gat), .B1(new_n933), .B2(new_n696), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n949), .A2(KEYINPUT125), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n949), .A2(KEYINPUT125), .ZN(new_n953));
  OR3_X1    g752(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n935), .A2(new_n470), .A3(new_n667), .A4(new_n936), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n951), .B2(new_n953), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(G1351gat));
  NOR3_X1   g756(.A1(new_n685), .A2(new_n574), .A3(new_n744), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT127), .Z(new_n959));
  NAND2_X1  g758(.A1(new_n904), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n300), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n935), .A2(new_n547), .A3(new_n889), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n963));
  INV_X1    g762(.A(G197gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n961), .B1(new_n966), .B2(new_n300), .ZN(G1352gat));
  NAND3_X1  g766(.A1(new_n962), .A2(new_n245), .A3(new_n248), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n969));
  OAI21_X1  g768(.A(G204gat), .B1(new_n960), .B2(new_n769), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n904), .A2(new_n650), .A3(new_n958), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(G211gat), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT63), .Z(new_n975));
  NAND4_X1  g774(.A1(new_n963), .A2(new_n333), .A3(new_n650), .A4(new_n965), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1354gat));
  NOR3_X1   g776(.A1(new_n960), .A2(new_n334), .A3(new_n696), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n667), .A3(new_n965), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n978), .B1(new_n979), .B2(new_n334), .ZN(G1355gat));
endmodule


