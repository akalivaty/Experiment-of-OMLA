//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n439, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(new_n439));
  INV_X1    g014(.A(new_n439), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(G234));
  NAND2_X1  g026(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(new_n439), .A2(G57), .A3(G69), .A4(G108), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT69), .Z(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT70), .Z(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT71), .B(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  INV_X1    g046(.A(new_n469), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n474), .A2(new_n482), .ZN(G160));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n470), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT72), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n470), .A2(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G112), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n476), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n488), .A2(G124), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n487), .A2(new_n492), .ZN(G162));
  AND2_X1   g068(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT3), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(G126), .A3(new_n467), .ZN(new_n497));
  NAND2_X1  g072(.A1(G114), .A2(G2104), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n484), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT4), .A2(G138), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n496), .A2(new_n484), .A3(new_n467), .A4(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n467), .A2(new_n477), .A3(G138), .A4(new_n484), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n484), .A2(G102), .A3(G2104), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n501), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n499), .A2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT73), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  INV_X1    g090(.A(new_n509), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G75), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n508), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n514), .A2(G88), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n516), .A2(G62), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n518), .A2(new_n525), .ZN(G166));
  NOR2_X1   g101(.A1(new_n513), .A2(new_n508), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT5), .B(G543), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n514), .A2(G89), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n522), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n528), .A2(new_n530), .A3(new_n535), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NOR2_X1   g114(.A1(new_n513), .A2(new_n522), .ZN(new_n540));
  AOI22_X1  g115(.A1(G52), .A2(new_n527), .B1(new_n540), .B2(G90), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n509), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n541), .B(KEYINPUT75), .C1(new_n509), .C2(new_n542), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n540), .A2(G81), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n514), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n534), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n509), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  OR2_X1    g135(.A1(KEYINPUT76), .A2(G65), .ZN(new_n561));
  NAND2_X1  g136(.A1(KEYINPUT76), .A2(G65), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n529), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n563), .A2(KEYINPUT77), .A3(new_n564), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n567), .A2(G651), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n540), .A2(G91), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n510), .A2(G53), .A3(G543), .A4(new_n512), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  OR2_X1    g150(.A1(new_n518), .A2(new_n525), .ZN(G303));
  NOR2_X1   g151(.A1(new_n522), .A2(new_n531), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(G74), .A2(G651), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n579), .A2(KEYINPUT78), .A3(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n582), .B(G651), .C1(new_n534), .C2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n510), .A2(G49), .A3(G543), .A4(new_n512), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n510), .A2(G87), .A3(new_n512), .A4(new_n529), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n516), .A2(G73), .ZN(new_n590));
  INV_X1    g165(.A(G48), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n513), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n516), .A2(G61), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n513), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(new_n529), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n534), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n509), .ZN(new_n600));
  AOI22_X1  g175(.A1(G47), .A2(new_n527), .B1(new_n540), .B2(G85), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n540), .A2(G92), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n529), .A2(G66), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT79), .ZN(new_n609));
  OAI21_X1  g184(.A(G651), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G54), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n550), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT80), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n606), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n603), .B1(G868), .B2(new_n617), .ZN(G284));
  OAI21_X1  g193(.A(new_n603), .B1(G868), .B2(new_n617), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  NOR2_X1   g200(.A1(new_n554), .A2(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n617), .A2(new_n624), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR3_X1   g205(.A1(new_n478), .A2(new_n469), .A3(G2105), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2100), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n486), .A2(G135), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(G111), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n476), .B1(new_n637), .B2(G2105), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n488), .A2(G123), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n634), .A2(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT82), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G1341), .B(G1348), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G14), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT83), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  XOR2_X1   g238(.A(new_n661), .B(KEYINPUT84), .Z(new_n664));
  OAI21_X1  g239(.A(KEYINPUT17), .B1(new_n664), .B2(new_n660), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(new_n659), .Z(new_n666));
  AND2_X1   g241(.A1(new_n664), .A2(new_n660), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n663), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2096), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n678));
  INV_X1    g253(.A(new_n673), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  AOI22_X1  g255(.A1(new_n677), .A2(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n680), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n682), .A2(new_n673), .A3(new_n676), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n681), .B(new_n683), .C1(new_n677), .C2(new_n678), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1986), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1991), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n686), .B(new_n689), .ZN(G229));
  NOR2_X1   g265(.A1(G5), .A2(G16), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G171), .B2(G16), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1961), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  OAI21_X1  g269(.A(KEYINPUT23), .B1(new_n621), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(G20), .ZN(new_n696));
  MUX2_X1   g271(.A(KEYINPUT23), .B(new_n695), .S(new_n696), .Z(new_n697));
  AOI21_X1  g272(.A(new_n693), .B1(G1956), .B2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G26), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  OR2_X1    g276(.A1(G104), .A2(G2105), .ZN(new_n702));
  INV_X1    g277(.A(G116), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n476), .B1(new_n703), .B2(G2105), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n488), .A2(G128), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT72), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n485), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G140), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n705), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n709), .A2(KEYINPUT88), .A3(G29), .ZN(new_n710));
  AOI21_X1  g285(.A(KEYINPUT88), .B1(new_n709), .B2(G29), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n701), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n699), .A2(G35), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G162), .B2(new_n699), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT29), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n698), .B1(G2067), .B2(new_n712), .C1(G2090), .C2(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n697), .A2(G1956), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(G2090), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n699), .A2(G33), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n484), .A2(G103), .A3(G2104), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT89), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT25), .ZN(new_n722));
  NAND2_X1  g297(.A1(G115), .A2(G2104), .ZN(new_n723));
  INV_X1    g298(.A(G127), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n478), .B2(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT90), .Z(new_n726));
  INV_X1    g301(.A(G139), .ZN(new_n727));
  OAI221_X1 g302(.A(new_n722), .B1(new_n726), .B2(new_n484), .C1(new_n707), .C2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT91), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n719), .B1(new_n729), .B2(G29), .ZN(new_n730));
  INV_X1    g305(.A(G2072), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n712), .A2(G2067), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n717), .A2(new_n718), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n730), .A2(new_n731), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n694), .A2(G4), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n617), .B2(new_n694), .ZN(new_n737));
  INV_X1    g312(.A(G1348), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n694), .A2(G19), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n554), .B2(new_n694), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G1341), .ZN(new_n742));
  INV_X1    g317(.A(G28), .ZN(new_n743));
  OR3_X1    g318(.A1(new_n743), .A2(KEYINPUT92), .A3(KEYINPUT30), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(KEYINPUT30), .ZN(new_n745));
  OAI21_X1  g320(.A(KEYINPUT92), .B1(new_n743), .B2(KEYINPUT30), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n744), .A2(new_n699), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n742), .B(new_n747), .C1(new_n699), .C2(new_n640), .ZN(new_n748));
  OR2_X1    g323(.A1(KEYINPUT24), .A2(G34), .ZN(new_n749));
  NAND2_X1  g324(.A1(KEYINPUT24), .A2(G34), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n749), .A2(new_n699), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G160), .B2(new_n699), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G2084), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n741), .B2(G1341), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT31), .B(G11), .Z(new_n755));
  NOR2_X1   g330(.A1(G27), .A2(G29), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G164), .B2(G29), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G2078), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(G2078), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n758), .B(new_n759), .C1(G2084), .C2(new_n752), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n748), .A2(new_n754), .A3(new_n755), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n694), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G168), .B2(new_n694), .ZN(new_n763));
  INV_X1    g338(.A(G1966), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n735), .A2(new_n739), .A3(new_n761), .A4(new_n765), .ZN(new_n766));
  OR3_X1    g341(.A1(new_n716), .A2(new_n734), .A3(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n699), .A2(G25), .ZN(new_n768));
  OR2_X1    g343(.A1(G95), .A2(G2105), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n769), .B(G2104), .C1(G107), .C2(new_n484), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT86), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n488), .A2(G119), .ZN(new_n772));
  INV_X1    g347(.A(G131), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n771), .B(new_n772), .C1(new_n707), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n768), .B1(new_n774), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT35), .B(G1991), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G290), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(new_n694), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n694), .B2(G24), .ZN(new_n781));
  INV_X1    g356(.A(G1986), .ZN(new_n782));
  OAI22_X1  g357(.A1(new_n781), .A2(new_n782), .B1(new_n777), .B2(new_n775), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n694), .A2(G22), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G166), .B2(new_n694), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1971), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT33), .B(G1976), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n694), .A2(G23), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT87), .B1(new_n584), .B2(new_n588), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT87), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n790), .B(new_n587), .C1(new_n581), .C2(new_n583), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n788), .B1(new_n793), .B2(new_n694), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n786), .B1(new_n787), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n694), .A2(G6), .ZN(new_n796));
  INV_X1    g371(.A(G305), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n694), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT32), .B(G1981), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n795), .B(new_n800), .C1(new_n787), .C2(new_n794), .ZN(new_n801));
  AOI211_X1 g376(.A(new_n778), .B(new_n783), .C1(new_n801), .C2(KEYINPUT34), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n781), .A2(new_n782), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT36), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(KEYINPUT36), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n767), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G29), .A2(G32), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n486), .A2(G141), .ZN(new_n810));
  NAND3_X1  g385(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT26), .Z(new_n812));
  NOR2_X1   g387(.A1(new_n469), .A2(G2105), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n488), .A2(G129), .B1(G105), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n810), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n809), .B1(new_n816), .B2(G29), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT27), .B(G1996), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n808), .A2(new_n820), .ZN(G311));
  NAND2_X1  g396(.A1(new_n808), .A2(new_n820), .ZN(G150));
  XNOR2_X1  g397(.A(KEYINPUT93), .B(G93), .ZN(new_n823));
  AOI22_X1  g398(.A1(G55), .A2(new_n527), .B1(new_n540), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n534), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n509), .B2(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT94), .B(G860), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n617), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  INV_X1    g406(.A(new_n826), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n551), .A2(new_n553), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n554), .A2(new_n826), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT39), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n831), .B(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n829), .B1(new_n838), .B2(new_n827), .ZN(G145));
  XOR2_X1   g414(.A(new_n709), .B(G164), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n815), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n729), .A2(KEYINPUT95), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n729), .A2(KEYINPUT95), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n840), .A2(new_n815), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n840), .A2(new_n815), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n845), .A2(KEYINPUT95), .A3(new_n729), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n488), .A2(G130), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n484), .A2(G118), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n476), .B1(new_n850), .B2(KEYINPUT96), .ZN(new_n851));
  OAI221_X1 g426(.A(new_n851), .B1(KEYINPUT96), .B2(new_n850), .C1(G106), .C2(G2105), .ZN(new_n852));
  INV_X1    g427(.A(G142), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n849), .B(new_n852), .C1(new_n707), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n774), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT97), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n632), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n855), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n632), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n848), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n844), .A2(new_n857), .A3(new_n861), .A4(new_n847), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n640), .B(G160), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G162), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT98), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n870));
  INV_X1    g445(.A(new_n867), .ZN(new_n871));
  AOI211_X1 g446(.A(new_n870), .B(new_n871), .C1(new_n863), .C2(new_n864), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n864), .A2(KEYINPUT99), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n857), .A2(new_n861), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n867), .B1(new_n879), .B2(new_n848), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n876), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n876), .A3(new_n880), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n874), .A2(new_n875), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n877), .A2(new_n876), .A3(new_n880), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(new_n881), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n868), .B2(new_n872), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT40), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n890), .ZN(G395));
  NAND2_X1  g466(.A1(new_n779), .A2(G303), .ZN(new_n892));
  NAND2_X1  g467(.A1(G166), .A2(G290), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(G305), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(G305), .B1(new_n892), .B2(new_n893), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n793), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n896), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(new_n792), .A3(new_n894), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n902));
  OR2_X1    g477(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(KEYINPUT101), .A3(KEYINPUT42), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n907));
  INV_X1    g482(.A(new_n836), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n627), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n616), .A2(G299), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n612), .B(new_n613), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n621), .A2(new_n911), .A3(new_n606), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n910), .A2(new_n912), .A3(KEYINPUT41), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT41), .B1(new_n910), .B2(new_n912), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n914), .B1(new_n917), .B2(new_n909), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n906), .B1(new_n907), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n918), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT102), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n906), .A3(KEYINPUT102), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(G868), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT103), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n922), .A2(new_n923), .A3(new_n926), .A4(G868), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n925), .B(new_n927), .C1(G868), .C2(new_n832), .ZN(G295));
  OAI211_X1 g503(.A(new_n925), .B(new_n927), .C1(G868), .C2(new_n832), .ZN(G331));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g505(.A1(G171), .A2(G286), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n545), .A2(G168), .A3(new_n546), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n836), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n908), .A2(new_n931), .A3(new_n932), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n915), .A2(new_n916), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n933), .A2(KEYINPUT104), .A3(new_n836), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n934), .A2(new_n935), .A3(new_n913), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n900), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(KEYINPUT105), .A3(new_n888), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n901), .B1(new_n940), .B2(new_n941), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(new_n946), .B2(G37), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n940), .A2(new_n901), .A3(new_n941), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n944), .A2(new_n947), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n930), .B1(new_n950), .B2(KEYINPUT106), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT105), .B1(new_n943), .B2(new_n888), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n946), .A2(new_n945), .A3(G37), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n954), .A2(new_n955), .A3(new_n948), .A4(new_n949), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n937), .A2(new_n939), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n934), .A2(new_n935), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n957), .A2(new_n913), .B1(new_n938), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n888), .B(new_n949), .C1(new_n959), .C2(new_n901), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n951), .A2(new_n956), .A3(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n944), .A2(new_n947), .A3(KEYINPUT43), .A4(new_n949), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n948), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n930), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(G397));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n499), .B2(new_n506), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n971));
  OAI211_X1 g546(.A(G40), .B(new_n481), .C1(new_n971), .C2(G2105), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(new_n815), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n709), .B(G2067), .Z(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n974), .B2(new_n816), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n973), .B(KEYINPUT108), .Z(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n976), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n774), .A2(new_n776), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n774), .A2(new_n776), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n779), .A2(new_n973), .A3(new_n782), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n973), .A2(G1986), .A3(G290), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n989), .B(KEYINPUT107), .Z(new_n990));
  NOR2_X1   g565(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  INV_X1    g567(.A(new_n972), .ZN(new_n993));
  INV_X1    g568(.A(new_n968), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(G305), .B(G1981), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n998), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n1000), .A3(new_n995), .ZN(new_n1001));
  INV_X1    g576(.A(G1976), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1001), .A2(new_n1002), .A3(new_n588), .A4(new_n584), .ZN(new_n1003));
  INV_X1    g578(.A(G1981), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n797), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n996), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n1007));
  NAND3_X1  g582(.A1(G303), .A2(new_n1007), .A3(G8), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1007), .B1(G303), .B2(G8), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT112), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1010), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n1013), .A3(new_n1008), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n968), .A2(new_n969), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n993), .B1(new_n1017), .B2(KEYINPUT109), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT45), .B(new_n967), .C1(new_n499), .C2(new_n506), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n970), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1016), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1020), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT109), .B1(new_n1017), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n972), .B1(new_n970), .B2(new_n1019), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(KEYINPUT110), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1971), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n968), .A2(KEYINPUT50), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n972), .B1(new_n1028), .B2(KEYINPUT111), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(new_n967), .C1(new_n499), .C2(new_n506), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n968), .A2(new_n1032), .A3(KEYINPUT50), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(G2090), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1015), .B(G8), .C1(new_n1027), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(KEYINPUT113), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G288), .A2(new_n790), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n584), .A2(KEYINPUT87), .A3(new_n588), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1002), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1039), .B1(new_n1042), .B2(new_n996), .ZN(new_n1043));
  NAND3_X1  g618(.A1(G288), .A2(new_n1037), .A3(new_n1002), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n995), .B(new_n1038), .C1(new_n792), .C2(new_n1002), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n1001), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1036), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1012), .A2(new_n1008), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1027), .A2(new_n1035), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(new_n1050), .B2(new_n992), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1033), .A2(new_n1031), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1032), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n1053));
  NOR4_X1   g628(.A1(new_n1052), .A2(new_n1053), .A3(G2084), .A4(new_n972), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n970), .A2(new_n993), .A3(new_n1020), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n764), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(G286), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1051), .A2(new_n1059), .A3(new_n1001), .A4(new_n1046), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n1006), .B(new_n1048), .C1(new_n1060), .C2(KEYINPUT63), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n1062));
  NAND3_X1  g637(.A1(G286), .A2(new_n1062), .A3(G8), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(G286), .B2(G8), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1065), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1063), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1069), .B2(KEYINPUT124), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1058), .A2(new_n1066), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT51), .B1(new_n1066), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G2084), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1029), .A2(new_n1074), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n992), .B1(new_n1075), .B2(new_n1056), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1073), .B1(new_n1076), .B2(new_n1069), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1069), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1071), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT125), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1071), .A2(new_n1077), .A3(KEYINPUT125), .A4(new_n1078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G2078), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1022), .A2(new_n1084), .A3(new_n1026), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1961), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1034), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1055), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1086), .A2(G2078), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1087), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  XOR2_X1   g668(.A(G171), .B(KEYINPUT54), .Z(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1083), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1047), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1046), .A2(KEYINPUT116), .A3(new_n1001), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1031), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n972), .B1(new_n1031), .B2(new_n1102), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(new_n1028), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(G2090), .B1(new_n1105), .B2(KEYINPUT115), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1103), .A2(new_n1104), .A3(new_n1107), .A4(new_n1028), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(G8), .B1(new_n1109), .B2(new_n1027), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1049), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1101), .A2(new_n1111), .A3(new_n1112), .A4(new_n1036), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT126), .B1(new_n1097), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1036), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1046), .A2(KEYINPUT116), .A3(new_n1001), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT116), .B1(new_n1046), .B2(new_n1001), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1095), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1112), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1114), .A2(new_n1122), .ZN(new_n1123));
  OR2_X1    g698(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n573), .A2(new_n570), .A3(new_n569), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT56), .B(G2072), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1024), .A2(new_n1025), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(G1956), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1105), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1034), .A2(new_n738), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n993), .A2(new_n994), .A3(KEYINPUT118), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT118), .B1(new_n993), .B2(new_n994), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1135), .A2(new_n1136), .A3(G2067), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n617), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1127), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1133), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1127), .B1(new_n1131), .B2(new_n1129), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT61), .B1(new_n1133), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1141), .A2(new_n1146), .A3(new_n1132), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT119), .B(G1996), .Z(new_n1149));
  NAND3_X1  g724(.A1(new_n1024), .A2(new_n1025), .A3(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT58), .B(G1341), .Z(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n833), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT121), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1157), .B1(new_n1153), .B2(KEYINPUT121), .ZN(new_n1158));
  NAND2_X1  g733(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1153), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1156), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1143), .B1(new_n1148), .B2(new_n1161), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1160), .A2(new_n1158), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1163), .A2(new_n1164), .A3(KEYINPUT122), .A4(new_n1156), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1167), .A2(KEYINPUT60), .A3(new_n616), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n616), .B1(new_n1167), .B2(KEYINPUT60), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n1168), .A2(new_n1169), .B1(KEYINPUT60), .B2(new_n1167), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1142), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1061), .B1(new_n1123), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1119), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1083), .A2(KEYINPUT62), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1081), .A2(new_n1175), .A3(new_n1082), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1174), .A2(G171), .A3(new_n1093), .A4(new_n1176), .ZN(new_n1177));
  OR3_X1    g752(.A1(new_n1058), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1173), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n991), .B1(new_n1172), .B2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n975), .B(KEYINPUT46), .Z(new_n1181));
  NAND2_X1  g756(.A1(new_n977), .A2(new_n816), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1181), .B1(new_n980), .B2(new_n1182), .ZN(new_n1183));
  XOR2_X1   g758(.A(new_n1183), .B(KEYINPUT47), .Z(new_n1184));
  NOR2_X1   g759(.A1(new_n709), .A2(G2067), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1185), .B1(new_n981), .B2(new_n982), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n987), .B(KEYINPUT48), .Z(new_n1187));
  OAI221_X1 g762(.A(new_n1184), .B1(new_n979), .B2(new_n1186), .C1(new_n986), .C2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n1188), .B(KEYINPUT127), .Z(new_n1189));
  NAND2_X1  g764(.A1(new_n1180), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g765(.A1(new_n656), .A2(new_n670), .ZN(new_n1192));
  INV_X1    g766(.A(new_n1192), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1193), .B1(new_n887), .B2(new_n889), .ZN(new_n1194));
  NOR2_X1   g768(.A1(G229), .A2(new_n464), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n963), .A2(new_n964), .A3(new_n1195), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n1194), .A2(new_n1196), .ZN(G308));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1198));
  OAI211_X1 g772(.A(new_n1198), .B(new_n1193), .C1(new_n889), .C2(new_n887), .ZN(G225));
endmodule


