//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957;
  INV_X1    g000(.A(G50gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G43gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(G43gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT15), .ZN(new_n206));
  NAND2_X1  g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NOR3_X1   g008(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n206), .B(new_n207), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(KEYINPUT86), .B(KEYINPUT15), .Z(new_n212));
  INV_X1    g011(.A(KEYINPUT87), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n203), .B1(new_n213), .B2(new_n205), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n202), .A2(KEYINPUT87), .A3(G43gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n210), .B1(KEYINPUT85), .B2(new_n208), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(KEYINPUT85), .B2(new_n208), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n206), .B1(new_n219), .B2(new_n207), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G1gat), .B2(new_n223), .ZN(new_n226));
  INV_X1    g025(.A(G8gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  OR3_X1    g028(.A1(new_n222), .A2(new_n229), .A3(KEYINPUT88), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n222), .A2(new_n229), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT88), .B1(new_n222), .B2(new_n229), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n234), .B(KEYINPUT13), .Z(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n228), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(new_n234), .A3(new_n231), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n239), .A2(KEYINPUT18), .A3(new_n234), .A4(new_n231), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n236), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(G169gat), .B(G197gat), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT12), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n236), .A2(new_n242), .A3(new_n243), .A4(new_n250), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(G211gat), .A2(G218gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT22), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n256), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n256), .B1(new_n260), .B2(new_n257), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G183gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT66), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G183gat), .ZN(new_n267));
  INV_X1    g066(.A(G190gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT24), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT24), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(G183gat), .A3(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G169gat), .ZN(new_n276));
  INV_X1    g075(.A(G176gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT23), .ZN(new_n278));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n278), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT23), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(G169gat), .B2(G176gat), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n285), .A2(KEYINPUT25), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n275), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n271), .A2(new_n273), .B1(new_n264), .B2(new_n268), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n278), .A2(new_n285), .A3(new_n279), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n294), .A2(new_n279), .ZN(new_n295));
  OR3_X1    g094(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n295), .A2(new_n296), .B1(G183gat), .B2(G190gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT27), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n268), .B1(new_n264), .B2(KEYINPUT27), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT28), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT27), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(G183gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n299), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n297), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n292), .A2(new_n293), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(new_n292), .B2(new_n306), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n263), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n292), .A2(new_n293), .A3(new_n306), .ZN(new_n313));
  INV_X1    g112(.A(new_n263), .ZN(new_n314));
  INV_X1    g113(.A(new_n305), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT66), .B(G183gat), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n299), .B1(new_n316), .B2(KEYINPUT27), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n317), .B2(KEYINPUT28), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n318), .A2(new_n297), .B1(new_n287), .B2(new_n291), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n313), .B(new_n314), .C1(new_n319), .C2(new_n310), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n312), .A2(KEYINPUT72), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT72), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n322), .B(new_n263), .C1(new_n307), .C2(new_n311), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT37), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT73), .ZN(new_n328));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(KEYINPUT38), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n312), .A2(new_n320), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n333), .B1(new_n334), .B2(KEYINPUT37), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n326), .A2(KEYINPUT83), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT83), .ZN(new_n337));
  INV_X1    g136(.A(new_n320), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n292), .A2(new_n306), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n309), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n314), .B1(new_n340), .B2(new_n313), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT37), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n332), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT37), .B1(new_n321), .B2(new_n323), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n337), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n336), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n324), .A2(new_n331), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n330), .B1(new_n324), .B2(new_n325), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT38), .B1(new_n348), .B2(new_n344), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT5), .ZN(new_n351));
  INV_X1    g150(.A(G127gat), .ZN(new_n352));
  INV_X1    g151(.A(G134gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G127gat), .A2(G134gat), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT1), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G120gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G113gat), .ZN(new_n358));
  INV_X1    g157(.A(G113gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G120gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n360), .A3(KEYINPUT68), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT69), .ZN(new_n362));
  OR3_X1    g161(.A1(new_n359), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n361), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n356), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G162gat), .ZN(new_n367));
  OR2_X1    g166(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT2), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT76), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n374));
  OAI21_X1  g173(.A(G162gat), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT2), .ZN(new_n377));
  INV_X1    g176(.A(G141gat), .ZN(new_n378));
  INV_X1    g177(.A(G148gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G141gat), .A2(G148gat), .ZN(new_n381));
  AND2_X1   g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n372), .A2(new_n377), .A3(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(KEYINPUT67), .B(G134gat), .Z(new_n387));
  AND2_X1   g186(.A1(new_n358), .A2(new_n360), .ZN(new_n388));
  OAI221_X1 g187(.A(new_n354), .B1(new_n387), .B2(new_n352), .C1(KEYINPUT1), .C2(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n371), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT74), .ZN(new_n391));
  OR2_X1    g190(.A1(new_n382), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n391), .B1(new_n382), .B2(new_n383), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n366), .A2(new_n386), .A3(new_n389), .A4(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G225gat), .A2(G233gat), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n375), .A2(KEYINPUT2), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n384), .B1(new_n400), .B2(KEYINPUT76), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n401), .B2(new_n377), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n402), .A2(KEYINPUT4), .A3(new_n366), .A4(new_n389), .ZN(new_n403));
  AND4_X1   g202(.A1(new_n351), .A2(new_n397), .A3(new_n398), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n394), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n405), .A2(KEYINPUT3), .B1(new_n366), .B2(new_n389), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT78), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT77), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n386), .A2(KEYINPUT77), .A3(new_n408), .A4(new_n394), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n406), .B(new_n407), .C1(new_n409), .C2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n386), .A2(new_n408), .A3(new_n394), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT77), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n410), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n407), .B1(new_n417), .B2(new_n406), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n404), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(G1gat), .B(G29gat), .Z(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G57gat), .B(G85gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n397), .A2(new_n398), .A3(new_n403), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n406), .B1(new_n409), .B2(new_n411), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT78), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n426), .B1(new_n428), .B2(new_n412), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n366), .A2(new_n389), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(new_n402), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT5), .B1(new_n431), .B2(new_n398), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n419), .B(new_n425), .C1(new_n429), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT80), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n419), .B1(new_n429), .B2(new_n432), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n424), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT6), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n426), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n413), .B2(new_n418), .ZN(new_n439));
  INV_X1    g238(.A(new_n432), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n428), .A2(new_n412), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n424), .B1(new_n442), .B2(new_n404), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n445), .A2(new_n446), .B1(new_n435), .B2(new_n424), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n350), .B1(new_n437), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT39), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n431), .B2(new_n398), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n397), .A2(new_n403), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n428), .B2(new_n412), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n452), .B2(new_n398), .ZN(new_n453));
  INV_X1    g252(.A(new_n451), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(new_n413), .B2(new_n418), .ZN(new_n455));
  INV_X1    g254(.A(new_n398), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n449), .A3(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n453), .A2(new_n457), .A3(KEYINPUT40), .A4(new_n425), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT30), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n347), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n321), .A2(new_n323), .A3(new_n330), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n324), .A2(KEYINPUT30), .A3(new_n331), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n436), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n398), .B1(new_n442), .B2(new_n454), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n424), .B1(new_n465), .B2(new_n449), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT40), .B1(new_n466), .B2(new_n453), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT82), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n405), .A2(new_n308), .A3(new_n314), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n405), .A2(KEYINPUT3), .ZN(new_n470));
  AND2_X1   g269(.A1(G228gat), .A2(G233gat), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT29), .B1(new_n416), .B2(new_n410), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(new_n314), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n308), .B1(new_n261), .B2(new_n262), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n475), .A2(KEYINPUT81), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT3), .B1(new_n475), .B2(KEYINPUT81), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n402), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n308), .B1(new_n409), .B2(new_n411), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n478), .B1(new_n479), .B2(new_n263), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n474), .B1(new_n480), .B2(new_n471), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G22gat), .ZN(new_n482));
  INV_X1    g281(.A(G22gat), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n474), .B(new_n483), .C1(new_n480), .C2(new_n471), .ZN(new_n484));
  XNOR2_X1  g283(.A(G78gat), .B(G106gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT31), .B(G50gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n482), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n482), .B2(new_n484), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n462), .A2(new_n461), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n492), .A2(new_n460), .B1(new_n435), .B2(new_n424), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n453), .A2(new_n457), .A3(new_n425), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT40), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT82), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n493), .A2(new_n496), .A3(new_n497), .A4(new_n458), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n448), .A2(new_n468), .A3(new_n491), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n444), .B1(new_n441), .B2(new_n443), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n425), .B1(new_n441), .B2(new_n419), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n446), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n446), .B1(new_n433), .B2(KEYINPUT80), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n436), .ZN(new_n504));
  INV_X1    g303(.A(new_n463), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT70), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n339), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n292), .A2(KEYINPUT70), .A3(new_n306), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(new_n430), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G227gat), .A2(G233gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT64), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n339), .A2(new_n507), .A3(new_n366), .A4(new_n389), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(KEYINPUT71), .B(KEYINPUT33), .Z(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(G15gat), .B(G43gat), .Z(new_n517));
  XNOR2_X1  g316(.A(G71gat), .B(G99gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n510), .A2(new_n513), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n512), .A2(KEYINPUT34), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n510), .A2(new_n513), .B1(G227gat), .B2(G233gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT34), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n514), .A2(KEYINPUT32), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n521), .A2(new_n511), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT34), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n527), .B1(new_n531), .B2(new_n523), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n520), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n526), .A2(new_n528), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n527), .A3(new_n523), .ZN(new_n535));
  INV_X1    g334(.A(new_n520), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(KEYINPUT36), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT36), .ZN(new_n539));
  INV_X1    g338(.A(new_n537), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n536), .B1(new_n534), .B2(new_n535), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n506), .A2(new_n490), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n499), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n533), .B(new_n537), .C1(new_n488), .C2(new_n489), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n437), .A2(new_n447), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .A4(new_n505), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT35), .B1(new_n506), .B2(new_n545), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n255), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G57gat), .B(G64gat), .Z(new_n553));
  NAND2_X1  g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n558), .A2(new_n554), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT89), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n553), .B(new_n556), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n553), .A2(new_n556), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n554), .A2(new_n558), .B1(new_n556), .B2(new_n560), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G127gat), .B(G155gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT90), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n568), .B(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G183gat), .B(G211gat), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n229), .B1(KEYINPUT21), .B2(new_n565), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n573), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n574), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n577), .B1(new_n574), .B2(new_n578), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT91), .B(G92gat), .Z(new_n582));
  INV_X1    g381(.A(G85gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT7), .ZN(new_n586));
  INV_X1    g385(.A(G99gat), .ZN(new_n587));
  INV_X1    g386(.A(G106gat), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT8), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n584), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G99gat), .B(G106gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n584), .A2(new_n591), .A3(new_n586), .A4(new_n589), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n237), .A2(new_n238), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT92), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n593), .A2(new_n594), .ZN(new_n600));
  AND2_X1   g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n222), .A2(new_n600), .B1(KEYINPUT41), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n596), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n601), .A2(KEYINPUT41), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n599), .B1(new_n596), .B2(new_n602), .ZN(new_n609));
  OR3_X1    g408(.A1(new_n604), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n608), .B1(new_n604), .B2(new_n609), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n581), .A2(KEYINPUT93), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT93), .B1(new_n581), .B2(new_n612), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n590), .A2(KEYINPUT95), .A3(new_n592), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n592), .A2(KEYINPUT95), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n616), .A2(new_n565), .A3(new_n594), .A4(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n600), .A2(KEYINPUT94), .A3(new_n565), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT94), .ZN(new_n621));
  INV_X1    g420(.A(new_n565), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(new_n595), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n600), .A2(KEYINPUT96), .A3(KEYINPUT10), .A4(new_n565), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n565), .A2(KEYINPUT10), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n595), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n618), .B1(new_n620), .B2(new_n623), .ZN(new_n633));
  INV_X1    g432(.A(new_n631), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT97), .ZN(new_n636));
  XOR2_X1   g435(.A(G120gat), .B(G148gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT98), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n633), .A2(new_n642), .A3(new_n634), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n632), .A2(new_n636), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n645));
  INV_X1    g444(.A(new_n635), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n634), .B1(new_n624), .B2(new_n629), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n640), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n644), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n645), .B1(new_n644), .B2(new_n648), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n552), .A2(new_n615), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n548), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(G1gat), .Z(G1324gat));
  INV_X1    g453(.A(new_n652), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n227), .B1(new_n655), .B2(new_n463), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT16), .B(G8gat), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n652), .A2(new_n505), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT42), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(KEYINPUT42), .B2(new_n658), .ZN(G1325gat));
  NAND2_X1  g459(.A1(new_n542), .A2(new_n538), .ZN(new_n661));
  OAI21_X1  g460(.A(G15gat), .B1(new_n652), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n533), .A2(new_n537), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n663), .A2(G15gat), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n662), .B1(new_n652), .B2(new_n664), .ZN(G1326gat));
  NOR2_X1   g464(.A1(new_n652), .A2(new_n491), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT43), .B(G22gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  INV_X1    g467(.A(new_n581), .ZN(new_n669));
  INV_X1    g468(.A(new_n612), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n670), .A3(new_n651), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT100), .Z(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n552), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(G29gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n548), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  INV_X1    g477(.A(new_n651), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n679), .A2(new_n255), .A3(new_n581), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n544), .A2(new_n551), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n670), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n610), .A2(KEYINPUT101), .A3(new_n611), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT101), .B1(new_n610), .B2(new_n611), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n681), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n544), .B2(new_n551), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n680), .B1(new_n683), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT102), .ZN(new_n690));
  INV_X1    g489(.A(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n682), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n612), .B1(new_n544), .B2(new_n551), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(new_n681), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n695), .A3(new_n680), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n690), .A2(new_n676), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n678), .B1(new_n697), .B2(new_n675), .ZN(G1328gat));
  NOR3_X1   g497(.A1(new_n673), .A2(G36gat), .A3(new_n505), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT46), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n690), .A2(new_n463), .A3(new_n696), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G36gat), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n701), .A2(new_n702), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n700), .B1(new_n704), .B2(new_n705), .ZN(G1329gat));
  OAI21_X1  g505(.A(G43gat), .B1(new_n689), .B2(new_n661), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n673), .A2(G43gat), .A3(new_n663), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n707), .A2(KEYINPUT47), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n661), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n690), .A2(new_n711), .A3(new_n696), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n708), .B1(new_n712), .B2(G43gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n710), .B1(new_n713), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g513(.A(G50gat), .B1(new_n689), .B2(new_n491), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n673), .A2(G50gat), .A3(new_n491), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n715), .A2(KEYINPUT48), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n690), .A2(new_n490), .A3(new_n696), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n719), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT105), .B1(new_n719), .B2(G50gat), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n720), .A2(new_n721), .A3(new_n716), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT104), .B(KEYINPUT48), .Z(new_n723));
  OAI21_X1  g522(.A(new_n718), .B1(new_n722), .B2(new_n723), .ZN(G1331gat));
  NOR4_X1   g523(.A1(new_n613), .A2(new_n614), .A3(new_n254), .A4(new_n651), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n682), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n676), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g528(.A(new_n505), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT106), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n732), .B(new_n733), .Z(G1333gat));
  OAI21_X1  g533(.A(G71gat), .B1(new_n726), .B2(new_n661), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n663), .A2(G71gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n726), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g537(.A1(new_n727), .A2(new_n490), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g539(.A1(new_n651), .A2(new_n581), .A3(new_n254), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n694), .A2(new_n676), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n583), .B1(new_n742), .B2(KEYINPUT107), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(KEYINPUT107), .B2(new_n742), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n581), .A2(new_n254), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n693), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT108), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n693), .A2(new_n749), .A3(KEYINPUT51), .A4(new_n745), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n748), .A2(new_n750), .B1(new_n747), .B2(new_n746), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n676), .A2(new_n679), .A3(new_n583), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n744), .B1(new_n751), .B2(new_n752), .ZN(G1336gat));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n651), .A2(G92gat), .A3(new_n505), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n582), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n694), .A2(new_n741), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(new_n505), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n754), .B1(new_n757), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n750), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n747), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n755), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n767), .A2(KEYINPUT111), .A3(new_n761), .A4(new_n760), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n746), .A2(KEYINPUT109), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT51), .B1(new_n746), .B2(KEYINPUT109), .ZN(new_n771));
  AOI22_X1  g570(.A1(new_n770), .A2(new_n771), .B1(new_n748), .B2(new_n750), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n760), .B1(new_n772), .B2(new_n756), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n773), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT110), .B1(new_n773), .B2(KEYINPUT52), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n769), .B1(new_n775), .B2(new_n776), .ZN(G1337gat));
  OAI21_X1  g576(.A(G99gat), .B1(new_n759), .B2(new_n661), .ZN(new_n778));
  INV_X1    g577(.A(new_n663), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n679), .A2(new_n587), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT112), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n751), .B2(new_n781), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n694), .A2(new_n490), .A3(new_n741), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT53), .B1(new_n783), .B2(G106gat), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n651), .A2(new_n491), .A3(G106gat), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n766), .A2(KEYINPUT115), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT115), .B1(new_n766), .B2(new_n785), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n785), .B(KEYINPUT114), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n772), .A2(new_n789), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n783), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT113), .B1(new_n783), .B2(G106gat), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n788), .B1(new_n793), .B2(new_n794), .ZN(G1339gat));
  NAND3_X1  g594(.A1(new_n624), .A2(new_n634), .A3(new_n629), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n632), .A2(KEYINPUT54), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n641), .B1(new_n647), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(KEYINPUT55), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT116), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n797), .A2(new_n799), .A3(new_n802), .A4(KEYINPUT55), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT55), .B1(new_n797), .B2(new_n799), .ZN(new_n805));
  INV_X1    g604(.A(new_n644), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n804), .A2(new_n254), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n233), .A2(new_n235), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n234), .B1(new_n239), .B2(new_n231), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n249), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(new_n253), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n649), .B2(new_n650), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n686), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  AND4_X1   g613(.A1(new_n686), .A2(new_n804), .A3(new_n812), .A4(new_n807), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n669), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n615), .A2(new_n255), .A3(new_n651), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n548), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n546), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n505), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n254), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n816), .A2(new_n817), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n491), .ZN(new_n825));
  AOI211_X1 g624(.A(KEYINPUT117), .B(new_n490), .C1(new_n816), .C2(new_n817), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR4_X1   g626(.A1(new_n827), .A2(new_n548), .A3(new_n463), .A4(new_n663), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n255), .A2(new_n359), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n822), .B1(new_n828), .B2(new_n829), .ZN(G1340gat));
  AOI21_X1  g629(.A(G120gat), .B1(new_n821), .B2(new_n679), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n651), .A2(new_n357), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n828), .B2(new_n832), .ZN(G1341gat));
  AOI21_X1  g632(.A(new_n352), .B1(new_n828), .B2(new_n581), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n820), .A2(G127gat), .A3(new_n669), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n834), .A2(new_n835), .ZN(G1342gat));
  INV_X1    g635(.A(new_n387), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n819), .A2(new_n505), .A3(new_n670), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n828), .A2(new_n670), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n841), .B1(new_n843), .B2(new_n353), .ZN(G1343gat));
  NOR2_X1   g643(.A1(new_n711), .A2(new_n491), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT120), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n818), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n463), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n378), .A3(new_n254), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n813), .A2(KEYINPUT119), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n813), .A2(KEYINPUT119), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n808), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n815), .B1(new_n853), .B2(new_n612), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n817), .B1(new_n854), .B2(new_n581), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n850), .B1(new_n855), .B2(new_n490), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n824), .A2(new_n490), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(KEYINPUT57), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n548), .A2(new_n463), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n661), .ZN(new_n860));
  NOR4_X1   g659(.A1(new_n856), .A2(new_n858), .A3(new_n255), .A4(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n849), .B1(new_n861), .B2(new_n378), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n379), .A3(new_n679), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n804), .A2(new_n670), .A3(new_n807), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(KEYINPUT121), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(KEYINPUT121), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n812), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n612), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n581), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n817), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n850), .B(new_n490), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n857), .A2(KEYINPUT57), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n875), .A2(new_n661), .A3(new_n679), .A4(new_n859), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n865), .B1(new_n876), .B2(G148gat), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n856), .A2(new_n858), .A3(new_n860), .ZN(new_n878));
  AOI211_X1 g677(.A(KEYINPUT59), .B(new_n379), .C1(new_n878), .C2(new_n679), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n864), .B1(new_n877), .B2(new_n879), .ZN(G1345gat));
  NOR2_X1   g679(.A1(new_n373), .A2(new_n374), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n848), .A2(new_n881), .A3(new_n581), .ZN(new_n882));
  INV_X1    g681(.A(new_n878), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n669), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n884), .B2(new_n881), .ZN(G1346gat));
  INV_X1    g684(.A(new_n686), .ZN(new_n886));
  OAI21_X1  g685(.A(G162gat), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n670), .A2(new_n505), .A3(new_n367), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n847), .B2(new_n888), .ZN(G1347gat));
  AOI21_X1  g688(.A(new_n676), .B1(new_n816), .B2(new_n817), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n890), .A2(new_n463), .A3(new_n546), .ZN(new_n891));
  AOI21_X1  g690(.A(G169gat), .B1(new_n891), .B2(new_n254), .ZN(new_n892));
  INV_X1    g691(.A(new_n827), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n676), .A2(new_n505), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n663), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n255), .A2(new_n276), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n892), .B1(new_n898), .B2(new_n899), .ZN(G1348gat));
  OAI21_X1  g699(.A(G176gat), .B1(new_n897), .B2(new_n651), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n891), .A2(new_n277), .A3(new_n679), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1349gat));
  OAI211_X1 g702(.A(new_n581), .B(new_n896), .C1(new_n825), .C2(new_n826), .ZN(new_n904));
  INV_X1    g703(.A(new_n316), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n264), .A2(KEYINPUT27), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n669), .A2(new_n906), .A3(new_n303), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n904), .A2(new_n905), .B1(new_n891), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(G1350gat));
  OAI211_X1 g711(.A(new_n670), .B(new_n896), .C1(new_n825), .C2(new_n826), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G190gat), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT61), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT123), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n914), .A2(new_n917), .A3(KEYINPUT61), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT124), .B1(new_n914), .B2(KEYINPUT61), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n913), .A2(new_n920), .A3(new_n921), .A4(G190gat), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n916), .A2(new_n918), .A3(new_n919), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n891), .A2(new_n268), .A3(new_n686), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1351gat));
  NOR3_X1   g724(.A1(new_n711), .A2(new_n491), .A3(new_n505), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n890), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n254), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n873), .A2(new_n874), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n895), .A2(new_n711), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n254), .A2(G197gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(G1352gat));
  NAND3_X1  g733(.A1(new_n875), .A2(new_n679), .A3(new_n930), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT125), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n932), .A2(new_n937), .A3(new_n679), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n936), .A2(G204gat), .A3(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n927), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n940), .A2(G204gat), .A3(new_n651), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT62), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n939), .A2(new_n942), .ZN(G1353gat));
  NAND4_X1  g742(.A1(new_n873), .A2(new_n581), .A3(new_n874), .A4(new_n930), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G211gat), .ZN(new_n945));
  NOR2_X1   g744(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n945), .A2(new_n946), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n669), .A2(G211gat), .ZN(new_n951));
  OAI22_X1  g750(.A1(new_n949), .A2(new_n950), .B1(new_n940), .B2(new_n951), .ZN(G1354gat));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n670), .B1(new_n932), .B2(new_n953), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n929), .A2(KEYINPUT127), .A3(new_n931), .ZN(new_n955));
  OAI21_X1  g754(.A(G218gat), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OR3_X1    g755(.A1(new_n940), .A2(G218gat), .A3(new_n886), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1355gat));
endmodule


