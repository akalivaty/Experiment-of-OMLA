//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT80), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT77), .ZN(new_n190));
  XNOR2_X1  g004(.A(G116), .B(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT5), .ZN(new_n192));
  INV_X1    g006(.A(G113), .ZN(new_n193));
  INV_X1    g007(.A(G116), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT5), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  XOR2_X1   g011(.A(KEYINPUT2), .B(G113), .Z(new_n198));
  AOI22_X1  g012(.A1(new_n192), .A2(new_n197), .B1(new_n198), .B2(new_n191), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(new_n200), .B2(G107), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G104), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n200), .A2(G107), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n201), .A2(new_n204), .A3(new_n205), .A4(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n200), .A2(G107), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n203), .A2(G104), .ZN(new_n209));
  OAI21_X1  g023(.A(G101), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n199), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n201), .A2(new_n204), .A3(new_n206), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n213), .A2(KEYINPUT73), .A3(G101), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT73), .B1(new_n213), .B2(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n207), .A2(KEYINPUT4), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n198), .A2(new_n191), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT2), .B(G113), .ZN(new_n219));
  INV_X1    g033(.A(G119), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(G116), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n219), .B1(new_n195), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n213), .A2(new_n224), .A3(G101), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n190), .B(new_n212), .C1(new_n217), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n213), .A2(G101), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT73), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n213), .A2(KEYINPUT73), .A3(G101), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n230), .A2(KEYINPUT4), .A3(new_n207), .A4(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n223), .A2(new_n225), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n232), .A2(new_n233), .B1(new_n211), .B2(new_n199), .ZN(new_n234));
  INV_X1    g048(.A(new_n190), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT78), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n227), .B(KEYINPUT6), .C1(new_n234), .C2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n212), .B1(new_n217), .B2(new_n226), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT6), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n239), .A2(new_n236), .A3(new_n240), .A4(new_n235), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G224), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(G953), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT79), .ZN(new_n245));
  XNOR2_X1  g059(.A(G143), .B(G146), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT0), .A3(G128), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT0), .B(G128), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G125), .ZN(new_n250));
  INV_X1    g064(.A(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G143), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT1), .B1(new_n253), .B2(G146), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(G128), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n252), .B(new_n254), .C1(KEYINPUT1), .C2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(G125), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n245), .B1(new_n250), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G125), .ZN(new_n263));
  OR2_X1    g077(.A1(new_n246), .A2(new_n248), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(new_n247), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(KEYINPUT79), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n244), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT79), .B1(new_n265), .B2(new_n260), .ZN(new_n268));
  INV_X1    g082(.A(new_n244), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n250), .A2(new_n245), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n188), .B1(new_n242), .B2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n272), .A2(new_n238), .A3(KEYINPUT80), .A4(new_n241), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G902), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT81), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n212), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n199), .A2(new_n211), .A3(KEYINPUT81), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n199), .A2(new_n211), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n190), .B(KEYINPUT8), .Z(new_n283));
  OAI21_X1  g097(.A(new_n227), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n269), .A2(KEYINPUT7), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n265), .B2(new_n260), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT7), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n271), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n277), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n187), .B1(new_n276), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n187), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n292), .B(new_n289), .C1(new_n274), .C2(new_n275), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G214), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OR3_X1    g110(.A1(new_n294), .A2(KEYINPUT82), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(G234), .A2(G237), .ZN(new_n298));
  INV_X1    g112(.A(G953), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n298), .A2(G952), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT21), .B(G898), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT93), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n298), .A2(G902), .A3(G953), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT82), .B1(new_n294), .B2(new_n296), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n297), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n299), .A2(G227), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(KEYINPUT72), .ZN(new_n310));
  XNOR2_X1  g124(.A(G110), .B(G140), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT65), .ZN(new_n314));
  INV_X1    g128(.A(G137), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(G134), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT64), .B1(new_n317), .B2(G137), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n318), .B2(KEYINPUT11), .ZN(new_n319));
  INV_X1    g133(.A(G131), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT11), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT64), .B(new_n321), .C1(new_n317), .C2(G137), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n320), .B1(new_n319), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n314), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n318), .A2(KEYINPUT11), .ZN(new_n326));
  INV_X1    g140(.A(new_n316), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G131), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(KEYINPUT65), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n257), .A2(new_n259), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n207), .A2(new_n210), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n257), .A2(new_n207), .A3(new_n210), .A4(new_n259), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT12), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT75), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n325), .A2(new_n331), .B1(new_n336), .B2(new_n335), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(KEYINPUT12), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n323), .A2(new_n324), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT12), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n339), .A2(new_n342), .B1(new_n337), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n336), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n257), .A2(new_n259), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n211), .A3(KEYINPUT10), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n225), .A2(new_n264), .A3(new_n247), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n348), .B(new_n350), .C1(new_n217), .C2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT74), .B1(new_n352), .B2(new_n332), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n350), .A2(new_n348), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n323), .A2(new_n324), .A3(new_n314), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT65), .B1(new_n329), .B2(new_n330), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT74), .ZN(new_n358));
  INV_X1    g172(.A(new_n249), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n232), .A2(new_n359), .A3(new_n225), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n354), .A2(new_n357), .A3(new_n358), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n353), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n313), .B1(new_n346), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n352), .A2(new_n332), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n312), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT76), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n313), .B1(new_n353), .B2(new_n361), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(KEYINPUT76), .ZN(new_n370));
  OAI211_X1 g184(.A(G469), .B(new_n364), .C1(new_n368), .C2(new_n370), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n353), .A2(new_n361), .B1(new_n332), .B2(new_n352), .ZN(new_n372));
  OAI22_X1  g186(.A1(new_n366), .A2(new_n346), .B1(new_n372), .B2(new_n312), .ZN(new_n373));
  INV_X1    g187(.A(G469), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n277), .ZN(new_n375));
  NAND2_X1  g189(.A1(G469), .A2(G902), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n371), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT9), .B(G234), .ZN(new_n378));
  OAI21_X1  g192(.A(G221), .B1(new_n378), .B2(G902), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n194), .A2(G122), .ZN(new_n382));
  INV_X1    g196(.A(G122), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(G116), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(new_n203), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT88), .B1(new_n258), .B2(G143), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT88), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n253), .A3(G128), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n258), .A2(G143), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n317), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT13), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n391), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT89), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n390), .A2(new_n397), .A3(new_n394), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n397), .B1(new_n390), .B2(new_n394), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n393), .B1(G134), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n385), .A2(new_n203), .ZN(new_n403));
  INV_X1    g217(.A(new_n392), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n317), .B1(new_n390), .B2(new_n391), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT14), .B1(new_n383), .B2(G116), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT90), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n382), .B1(new_n409), .B2(new_n384), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n203), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G217), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n378), .A2(new_n413), .A3(G953), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n402), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n401), .A2(G134), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n386), .A2(new_n392), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n406), .A2(new_n411), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n414), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(KEYINPUT92), .B(new_n277), .C1(new_n416), .C2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G478), .ZN(new_n423));
  NOR2_X1   g237(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n415), .B1(new_n402), .B2(new_n412), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n419), .A2(new_n420), .A3(new_n414), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n427), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n431), .A2(KEYINPUT92), .A3(new_n277), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT17), .ZN(new_n436));
  INV_X1    g250(.A(G237), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n299), .A3(G214), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(new_n253), .ZN(new_n440));
  NOR2_X1   g254(.A1(G237), .A2(G953), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n441), .B(G214), .C1(KEYINPUT83), .C2(G143), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G131), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n320), .B1(new_n440), .B2(new_n442), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n436), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n445), .A2(new_n436), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n449));
  INV_X1    g263(.A(G140), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G125), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n263), .A2(G140), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT16), .ZN(new_n453));
  OR3_X1    g267(.A1(new_n263), .A2(KEYINPUT16), .A3(G140), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n453), .A2(G146), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(G146), .B1(new_n453), .B2(new_n454), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT69), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AND4_X1   g272(.A1(new_n457), .A2(new_n453), .A3(G146), .A4(new_n454), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n449), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n456), .A2(new_n457), .ZN(new_n461));
  INV_X1    g275(.A(new_n455), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n459), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(KEYINPUT85), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n448), .A2(new_n460), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G113), .B(G122), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(new_n200), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n451), .A2(new_n452), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(new_n251), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n443), .A2(KEYINPUT18), .A3(G131), .ZN(new_n471));
  NAND2_X1  g285(.A1(KEYINPUT18), .A2(G131), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n440), .A2(new_n472), .A3(new_n442), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n466), .A2(new_n468), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT19), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT84), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n478));
  MUX2_X1   g292(.A(new_n477), .B(new_n478), .S(new_n469), .Z(new_n479));
  OAI21_X1  g293(.A(new_n462), .B1(new_n479), .B2(G146), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n444), .A2(new_n445), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n474), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n468), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n475), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n486));
  NOR2_X1   g300(.A1(G475), .A2(G902), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT20), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n466), .A2(new_n474), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n483), .ZN(new_n490));
  AOI21_X1  g304(.A(G902), .B1(new_n490), .B2(new_n475), .ZN(new_n491));
  INV_X1    g305(.A(G475), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n486), .A2(KEYINPUT20), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n486), .A2(KEYINPUT20), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI211_X1 g310(.A(new_n494), .B(new_n496), .C1(new_n485), .C2(new_n487), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT87), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n494), .B1(new_n485), .B2(new_n487), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n495), .ZN(new_n500));
  INV_X1    g314(.A(new_n475), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n468), .B1(new_n466), .B2(new_n474), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n277), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G475), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n500), .A2(new_n504), .A3(new_n505), .A4(new_n488), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n381), .A2(new_n435), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n308), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n359), .B1(new_n355), .B2(new_n356), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n317), .A2(G137), .ZN(new_n511));
  OAI21_X1  g325(.A(G131), .B1(new_n511), .B2(new_n316), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n349), .A2(new_n330), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(KEYINPUT30), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n513), .B1(new_n343), .B2(new_n249), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT30), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n223), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n513), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n332), .B2(new_n359), .ZN(new_n520));
  INV_X1    g334(.A(new_n223), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT66), .B(KEYINPUT27), .Z(new_n524));
  NAND2_X1  g338(.A1(new_n441), .A2(G210), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT26), .B(G101), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n515), .A2(new_n223), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT28), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n520), .B2(new_n521), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n249), .B1(new_n325), .B2(new_n331), .ZN(new_n533));
  NOR4_X1   g347(.A1(new_n533), .A2(new_n519), .A3(KEYINPUT28), .A4(new_n223), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n530), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n528), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT29), .B1(new_n529), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n223), .B1(new_n533), .B2(new_n519), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n532), .B2(new_n534), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n536), .A2(KEYINPUT29), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n277), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G472), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n528), .B1(new_n520), .B2(new_n521), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n518), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT67), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT67), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n518), .A2(new_n546), .A3(new_n549), .A4(new_n545), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n518), .A2(new_n546), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n535), .A2(new_n528), .B1(new_n552), .B2(KEYINPUT31), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(G472), .A2(G902), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n544), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n555), .ZN(new_n557));
  AOI211_X1 g371(.A(KEYINPUT32), .B(new_n557), .C1(new_n551), .C2(new_n553), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n543), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n413), .B1(G234), .B2(new_n277), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n258), .B(G119), .C1(KEYINPUT68), .C2(KEYINPUT23), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT23), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n220), .B2(G128), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT68), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n220), .B2(G128), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n561), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(G119), .B(G128), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT24), .B(G110), .Z(new_n568));
  AOI22_X1  g382(.A1(new_n566), .A2(G110), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n463), .A2(new_n464), .A3(new_n569), .ZN(new_n570));
  OAI22_X1  g384(.A1(new_n566), .A2(G110), .B1(new_n567), .B2(new_n568), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n469), .A2(new_n251), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n462), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n299), .A2(G221), .A3(G234), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT70), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT22), .B(G137), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n574), .B(new_n578), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n579), .A2(KEYINPUT25), .A3(new_n277), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT25), .B1(new_n579), .B2(new_n277), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n560), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n560), .A2(G902), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT71), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n559), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n509), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n276), .A2(new_n290), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n292), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n276), .A2(new_n187), .A3(new_n290), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(KEYINPUT94), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n296), .B1(new_n293), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n306), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n423), .A2(new_n277), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n416), .A2(new_n421), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(G902), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n599), .B1(new_n601), .B2(new_n423), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n431), .A2(KEYINPUT33), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n431), .A2(KEYINPUT33), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(G478), .A3(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n498), .A2(new_n606), .A3(new_n506), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n591), .B1(new_n598), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n276), .A2(new_n596), .A3(new_n187), .A4(new_n290), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n295), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n294), .B2(KEYINPUT94), .ZN(new_n611));
  INV_X1    g425(.A(new_n607), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n611), .A2(new_n612), .A3(KEYINPUT95), .A4(new_n306), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n380), .A2(new_n586), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n551), .B2(new_n553), .ZN(new_n616));
  INV_X1    g430(.A(G472), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n557), .B1(new_n551), .B2(new_n553), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(new_n200), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT96), .B(KEYINPUT34), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  NOR2_X1   g439(.A1(new_n493), .A2(new_n497), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n611), .A2(new_n306), .A3(new_n434), .A4(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  INV_X1    g445(.A(KEYINPUT36), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n578), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n574), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n584), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n582), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n618), .A2(new_n619), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n509), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  AND3_X1   g455(.A1(new_n559), .A2(new_n381), .A3(new_n636), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n434), .A2(new_n500), .A3(new_n504), .A4(new_n488), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT97), .B(G900), .Z(new_n644));
  AOI21_X1  g458(.A(new_n300), .B1(new_n644), .B2(new_n304), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT98), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n647));
  INV_X1    g461(.A(new_n645), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n626), .A2(new_n647), .A3(new_n434), .A4(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(KEYINPUT99), .A3(new_n611), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n646), .A2(new_n649), .A3(new_n595), .A4(new_n597), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n642), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT100), .B(G128), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G30));
  NOR2_X1   g471(.A1(new_n523), .A2(new_n528), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n522), .A2(new_n528), .A3(new_n539), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n277), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n661), .B1(new_n556), .B2(new_n558), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(KEYINPUT102), .Z(new_n663));
  XOR2_X1   g477(.A(new_n645), .B(KEYINPUT39), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n381), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT40), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n294), .B(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n507), .A2(new_n435), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n295), .A3(new_n637), .ZN(new_n670));
  OR4_X1    g484(.A1(new_n663), .A2(new_n666), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G143), .ZN(G45));
  NAND4_X1  g486(.A1(new_n498), .A2(new_n606), .A3(new_n506), .A4(new_n648), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n611), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n642), .A2(KEYINPUT103), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n559), .A2(new_n381), .A3(new_n636), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n678), .B1(new_n679), .B2(new_n675), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  NAND2_X1  g496(.A1(new_n373), .A2(new_n277), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n374), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n373), .B(new_n277), .C1(new_n684), .C2(new_n374), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n379), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n559), .A2(new_n587), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n614), .A2(new_n691), .A3(KEYINPUT105), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT105), .B1(new_n614), .B2(new_n691), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT41), .B(G113), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT106), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n694), .B(new_n696), .ZN(G15));
  NAND3_X1  g511(.A1(new_n691), .A2(new_n628), .A3(KEYINPUT107), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(new_n690), .B2(new_n627), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT108), .B(G116), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G18));
  NAND2_X1  g517(.A1(new_n595), .A2(new_n597), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n688), .ZN(new_n705));
  AOI211_X1 g519(.A(new_n305), .B(new_n434), .C1(new_n498), .C2(new_n506), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n559), .A3(new_n636), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  NAND2_X1  g522(.A1(new_n554), .A2(new_n277), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G472), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n540), .A2(new_n528), .B1(new_n552), .B2(KEYINPUT31), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n551), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n555), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n710), .A2(new_n587), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n688), .A2(new_n305), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n611), .A3(new_n669), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G122), .ZN(G24));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n713), .B(new_n636), .C1(new_n617), .C2(new_n616), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT109), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n710), .A2(new_n721), .A3(new_n636), .A4(new_n713), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n718), .A2(new_n723), .A3(new_n674), .A4(new_n705), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n673), .B1(new_n720), .B2(new_n722), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n718), .B1(new_n725), .B2(new_n705), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n263), .ZN(G27));
  AND4_X1   g542(.A1(new_n295), .A2(new_n377), .A3(new_n294), .A4(new_n379), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(KEYINPUT42), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n588), .A2(new_n674), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n729), .A2(new_n587), .A3(new_n559), .A4(new_n674), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n731), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  AND3_X1   g551(.A1(new_n729), .A2(new_n587), .A3(new_n559), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n650), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT112), .B(G134), .Z(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G36));
  OR2_X1    g555(.A1(new_n368), .A2(new_n370), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n364), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n374), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(KEYINPUT113), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n742), .A2(KEYINPUT45), .A3(new_n364), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT114), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(KEYINPUT113), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n376), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(KEYINPUT46), .A3(new_n376), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n375), .A3(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n755), .A2(new_n379), .A3(new_n664), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n291), .A2(new_n293), .A3(new_n296), .ZN(new_n757));
  XOR2_X1   g571(.A(new_n757), .B(KEYINPUT115), .Z(new_n758));
  AND2_X1   g572(.A1(new_n498), .A2(new_n506), .ZN(new_n759));
  INV_X1    g573(.A(new_n606), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT43), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n620), .A2(new_n637), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n758), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n756), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  INV_X1    g584(.A(new_n559), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n586), .A3(new_n674), .A4(new_n757), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n755), .A2(KEYINPUT47), .A3(new_n379), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT47), .B1(new_n755), .B2(new_n379), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n379), .A2(new_n377), .A3(new_n637), .A4(new_n648), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(new_n662), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n704), .A2(new_n435), .A3(new_n507), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT103), .B1(new_n642), .B2(new_n676), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n679), .A2(new_n675), .A3(new_n678), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n655), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n779), .B1(new_n786), .B2(new_n727), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n725), .A2(new_n705), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT110), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n725), .A2(new_n718), .A3(new_n705), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n652), .A2(new_n653), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n679), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n793), .A2(new_n654), .B1(new_n782), .B2(new_n781), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n791), .A2(KEYINPUT52), .A3(new_n681), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n509), .B1(new_n588), .B2(new_n638), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n507), .A2(new_n435), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n760), .A2(new_n498), .A3(new_n506), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n615), .A2(new_n798), .A3(new_n620), .A4(new_n799), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(new_n308), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n707), .A2(new_n716), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n701), .A2(new_n797), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n434), .A2(new_n645), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n559), .A2(new_n626), .A3(new_n636), .A4(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n729), .B1(new_n725), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n736), .A2(new_n739), .A3(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n803), .A2(new_n694), .A3(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n796), .A2(KEYINPUT53), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n811), .B(new_n779), .C1(new_n786), .C2(new_n727), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n795), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n794), .B(new_n681), .C1(new_n724), .C2(new_n726), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n811), .B1(new_n814), .B2(new_n779), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n808), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n809), .B1(new_n810), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n778), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n787), .A2(KEYINPUT117), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n812), .A3(new_n795), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT53), .B1(new_n821), .B2(new_n808), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT118), .B(KEYINPUT54), .C1(new_n822), .C2(new_n809), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n796), .A2(new_n810), .A3(new_n808), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(KEYINPUT53), .B2(new_n816), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n825), .B1(new_n827), .B2(KEYINPUT54), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n816), .A2(KEYINPUT53), .ZN(new_n829));
  INV_X1    g643(.A(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(KEYINPUT119), .A3(new_n818), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n755), .A2(new_n379), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT47), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n755), .A2(KEYINPUT47), .A3(new_n379), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n686), .A2(new_n687), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n379), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n835), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n762), .A2(new_n300), .A3(new_n714), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n842), .A2(new_n758), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n689), .A2(new_n757), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n845), .A2(new_n587), .A3(new_n300), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n663), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT122), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n759), .A2(new_n606), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n762), .A2(new_n300), .A3(new_n845), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n723), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n855));
  OR2_X1    g669(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n668), .A2(new_n296), .A3(new_n689), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n842), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(KEYINPUT120), .B(KEYINPUT50), .C1(new_n841), .C2(new_n857), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n859), .A2(new_n860), .A3(KEYINPUT51), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n844), .A2(new_n854), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n851), .A2(new_n588), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT48), .ZN(new_n864));
  INV_X1    g678(.A(G952), .ZN(new_n865));
  AOI211_X1 g679(.A(new_n865), .B(G953), .C1(new_n842), .C2(new_n705), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n612), .B2(new_n848), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n853), .B1(new_n840), .B2(new_n843), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n859), .A2(new_n860), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n871), .B(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT51), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n824), .A2(new_n828), .A3(new_n832), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n865), .A2(new_n299), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n587), .A2(new_n295), .A3(new_n379), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n837), .B2(KEYINPUT49), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(new_n668), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n837), .A2(KEYINPUT49), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT116), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n663), .A2(new_n761), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n878), .A2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n831), .A2(new_n277), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(G210), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n242), .B(KEYINPUT123), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n272), .B(KEYINPUT55), .Z(new_n890));
  XNOR2_X1  g704(.A(new_n889), .B(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n887), .B2(new_n888), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n299), .A2(G952), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(G51));
  XNOR2_X1  g709(.A(new_n827), .B(new_n818), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n376), .B(KEYINPUT57), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n373), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OR3_X1    g712(.A1(new_n831), .A2(new_n277), .A3(new_n750), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(G54));
  NAND3_X1  g714(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n475), .A3(new_n484), .ZN(new_n902));
  INV_X1    g716(.A(new_n894), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .A4(new_n485), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G60));
  NAND2_X1  g719(.A1(new_n603), .A2(new_n604), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n599), .B(KEYINPUT59), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n903), .B1(new_n896), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n816), .A2(new_n810), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n796), .A2(new_n808), .A3(KEYINPUT53), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT118), .B1(new_n913), .B2(KEYINPUT54), .ZN(new_n914));
  AOI211_X1 g728(.A(new_n778), .B(new_n818), .C1(new_n911), .C2(new_n912), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n828), .A2(new_n832), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n908), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n906), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n910), .B1(new_n918), .B2(new_n919), .ZN(G63));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT60), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n827), .A2(new_n634), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n831), .A2(new_n922), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n903), .B(new_n924), .C1(new_n925), .C2(new_n579), .ZN(new_n926));
  XOR2_X1   g740(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(G66));
  OAI21_X1  g742(.A(G953), .B1(new_n303), .B2(new_n243), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n803), .A2(new_n694), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT125), .Z(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n931), .B2(G953), .ZN(new_n932));
  INV_X1    g746(.A(new_n889), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(G898), .B2(new_n299), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n932), .B(new_n934), .ZN(G69));
  AND2_X1   g749(.A1(new_n514), .A2(new_n517), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(new_n479), .Z(new_n937));
  AOI21_X1  g751(.A(new_n772), .B1(new_n835), .B2(new_n836), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n755), .A2(new_n379), .A3(new_n664), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n736), .B(new_n739), .C1(new_n939), .C2(new_n767), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n791), .A2(new_n655), .A3(new_n681), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n588), .A2(new_n782), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n941), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n938), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n944), .A2(G953), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n299), .A2(G900), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n937), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n738), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n798), .A2(new_n664), .A3(new_n799), .ZN(new_n949));
  OAI22_X1  g763(.A1(new_n939), .A2(new_n767), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n938), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n941), .A2(new_n671), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n941), .A2(new_n671), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n951), .A2(KEYINPUT126), .A3(new_n953), .A4(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n948), .A2(new_n949), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n756), .B2(new_n768), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n776), .A2(new_n958), .A3(new_n955), .A4(new_n953), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(G953), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n947), .B1(new_n962), .B2(new_n937), .ZN(new_n963));
  INV_X1    g777(.A(G227), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n946), .B1(new_n964), .B2(G953), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n966), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n947), .B(new_n968), .C1(new_n962), .C2(new_n937), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(G72));
  INV_X1    g784(.A(new_n658), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n956), .A2(new_n961), .A3(new_n931), .ZN(new_n972));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT63), .Z(new_n974));
  AOI21_X1  g788(.A(new_n971), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n974), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n944), .B2(new_n931), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n903), .B1(new_n977), .B2(new_n529), .ZN(new_n978));
  AND4_X1   g792(.A1(new_n529), .A2(new_n913), .A3(new_n971), .A4(new_n974), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(G57));
endmodule


