//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT64), .B(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G58), .A2(G232), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n205), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n208), .B(new_n214), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(KEYINPUT13), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT3), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n248));
  OAI21_X1  g0048(.A(KEYINPUT68), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n245), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT68), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n249), .A2(G226), .A3(new_n250), .A4(new_n254), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n249), .A2(G232), .A3(G1698), .A4(new_n254), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G97), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT66), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n261), .A2(new_n265), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(G1), .A2(G13), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n269), .B1(new_n276), .B2(new_n217), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n244), .B1(new_n260), .B2(new_n278), .ZN(new_n279));
  AOI211_X1 g0079(.A(KEYINPUT13), .B(new_n277), .C1(new_n258), .C2(new_n259), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT75), .A2(G169), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT14), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT14), .ZN(new_n284));
  INV_X1    g0084(.A(new_n282), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n284), .B(new_n285), .C1(new_n279), .C2(new_n280), .ZN(new_n286));
  AOI21_X1  g0086(.A(KEYINPUT76), .B1(new_n281), .B2(G179), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT76), .ZN(new_n288));
  INV_X1    g0088(.A(G179), .ZN(new_n289));
  NOR4_X1   g0089(.A1(new_n279), .A2(new_n280), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n283), .B(new_n286), .C1(new_n287), .C2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n211), .ZN(new_n293));
  INV_X1    g0093(.A(G77), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n212), .A2(G33), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n215), .A2(new_n212), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G50), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n296), .A2(KEYINPUT74), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n296), .A2(KEYINPUT74), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n293), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT11), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G13), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n305), .A2(new_n212), .A3(G1), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(new_n293), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n271), .A2(G20), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(G68), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT12), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n305), .A2(G1), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G20), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n310), .B1(new_n312), .B2(G68), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n216), .A2(KEYINPUT12), .A3(G20), .A4(new_n311), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n309), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n302), .B2(new_n303), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n304), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n291), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n281), .A2(G190), .ZN(new_n320));
  OAI21_X1  g0120(.A(G200), .B1(new_n279), .B2(new_n280), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n249), .A2(G222), .A3(new_n250), .A4(new_n254), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n249), .A2(G223), .A3(G1698), .A4(new_n254), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n249), .A2(new_n254), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n325), .B(new_n326), .C1(new_n328), .C2(new_n294), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n259), .ZN(new_n330));
  INV_X1    g0130(.A(G226), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n269), .B1(new_n276), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT67), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n324), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n334), .A2(KEYINPUT73), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n330), .A2(new_n333), .A3(G190), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT8), .B(G58), .ZN(new_n337));
  INV_X1    g0137(.A(G150), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n337), .A2(new_n295), .B1(new_n338), .B2(new_n299), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n212), .B1(new_n201), .B2(new_n297), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n293), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n297), .B1(new_n271), .B2(G20), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n307), .A2(new_n342), .B1(new_n297), .B2(new_n306), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n341), .A2(KEYINPUT9), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT9), .B1(new_n341), .B2(new_n343), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n336), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n334), .A2(KEYINPUT73), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n335), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT10), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT10), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n335), .A2(new_n347), .A3(new_n351), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n341), .A2(new_n343), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n330), .A2(new_n333), .ZN(new_n355));
  AND2_X1   g0155(.A1(KEYINPUT69), .A2(G179), .ZN(new_n356));
  NOR2_X1   g0156(.A1(KEYINPUT69), .A2(G179), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G169), .ZN(new_n360));
  AOI211_X1 g0160(.A(new_n354), .B(new_n359), .C1(new_n360), .C2(new_n355), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n353), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n328), .A2(G238), .A3(G1698), .ZN(new_n364));
  INV_X1    g0164(.A(G107), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n328), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n327), .A2(new_n228), .A3(G1698), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n259), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G244), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n269), .B1(new_n276), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT70), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n360), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT15), .B(G87), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n374), .A2(new_n295), .B1(new_n212), .B2(new_n294), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n337), .B(KEYINPUT71), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n298), .ZN(new_n377));
  INV_X1    g0177(.A(new_n293), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT72), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n307), .A2(G77), .A3(new_n308), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G77), .B2(new_n312), .ZN(new_n382));
  OR3_X1    g0182(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n380), .B1(new_n379), .B2(new_n382), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n373), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n368), .A2(new_n371), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n356), .A2(new_n357), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n387), .A2(new_n324), .ZN(new_n391));
  INV_X1    g0191(.A(G190), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n384), .B(new_n383), .C1(new_n372), .C2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n390), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n251), .A2(new_n252), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n395), .B2(new_n212), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  AOI211_X1 g0197(.A(new_n397), .B(G20), .C1(new_n251), .C2(new_n252), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(KEYINPUT64), .A2(G68), .ZN(new_n400));
  NOR2_X1   g0200(.A1(KEYINPUT64), .A2(G68), .ZN(new_n401));
  OAI21_X1  g0201(.A(G58), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n202), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n403), .A2(G20), .B1(G159), .B2(new_n298), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n399), .A2(KEYINPUT16), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n201), .B1(new_n215), .B2(G58), .ZN(new_n406));
  INV_X1    g0206(.A(G159), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n406), .A2(new_n212), .B1(new_n407), .B2(new_n299), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n395), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n409));
  AOI21_X1  g0209(.A(G20), .B1(new_n249), .B2(new_n254), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(KEYINPUT7), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n408), .B1(new_n411), .B2(new_n215), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n293), .B(new_n405), .C1(new_n412), .C2(KEYINPUT16), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT78), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n269), .B1(new_n276), .B2(new_n228), .ZN(new_n415));
  OR2_X1    g0215(.A1(G223), .A2(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n331), .A2(G1698), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n251), .A2(new_n416), .A3(new_n252), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n275), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n415), .A2(new_n420), .A3(G190), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n419), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n259), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n271), .A2(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(G232), .B1(new_n266), .B2(new_n268), .ZN(new_n425));
  AOI21_X1  g0225(.A(G200), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n414), .B1(new_n421), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n392), .A3(new_n425), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n415), .A2(new_n420), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n428), .B(KEYINPUT78), .C1(new_n429), .C2(G200), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n307), .ZN(new_n432));
  INV_X1    g0232(.A(new_n337), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n308), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n432), .A2(new_n434), .B1(new_n312), .B2(new_n433), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n413), .A2(new_n431), .A3(KEYINPUT79), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n253), .B1(new_n251), .B2(new_n252), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n212), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n398), .B1(new_n442), .B2(new_n397), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n404), .B1(new_n443), .B2(new_n216), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT16), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n405), .A2(new_n293), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n435), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n448), .A2(KEYINPUT79), .A3(KEYINPUT17), .A4(new_n431), .ZN(new_n449));
  OAI21_X1  g0249(.A(G169), .B1(new_n415), .B2(new_n420), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n423), .A2(new_n358), .A3(new_n425), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT77), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT77), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT18), .B1(new_n448), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n454), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n452), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT18), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n405), .A2(new_n293), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n445), .B2(new_n444), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n458), .B(new_n459), .C1(new_n461), .C2(new_n435), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n439), .A2(new_n449), .A3(new_n456), .A4(new_n462), .ZN(new_n463));
  NOR4_X1   g0263(.A1(new_n323), .A2(new_n363), .A3(new_n394), .A4(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n311), .ZN(new_n465));
  INV_X1    g0265(.A(G116), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G20), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  INV_X1    g0269(.A(G97), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n469), .B(new_n212), .C1(G33), .C2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(new_n293), .A3(new_n467), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT20), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n473), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT86), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n271), .A2(G33), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n378), .A2(new_n312), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n479), .B2(new_n466), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n307), .A2(KEYINPUT86), .A3(G116), .A4(new_n478), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n262), .A2(new_n264), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT5), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n271), .B(G45), .C1(new_n485), .C2(G41), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n486), .A2(new_n488), .A3(G274), .A4(new_n275), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT5), .B1(new_n262), .B2(new_n264), .ZN(new_n490));
  OAI211_X1 g0290(.A(G270), .B(new_n275), .C1(new_n490), .C2(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G303), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n249), .B2(new_n254), .ZN(new_n495));
  XNOR2_X1  g0295(.A(KEYINPUT3), .B(G33), .ZN(new_n496));
  INV_X1    g0296(.A(G257), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n250), .ZN(new_n498));
  OR2_X1    g0298(.A1(new_n250), .A2(G264), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n259), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n483), .A2(new_n503), .A3(G169), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n327), .A2(G303), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n275), .B1(new_n507), .B2(new_n500), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n508), .A2(new_n289), .A3(new_n492), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n483), .ZN(new_n510));
  OAI21_X1  g0310(.A(G200), .B1(new_n508), .B2(new_n492), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n493), .A2(G190), .A3(new_n502), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n511), .A2(new_n482), .A3(new_n476), .A4(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n483), .A2(new_n503), .A3(KEYINPUT21), .A4(G169), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n506), .A2(new_n510), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT87), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n510), .A2(new_n514), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT87), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(new_n506), .A4(new_n513), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n217), .A2(new_n250), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n369), .A2(G1698), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n251), .A2(new_n521), .A3(new_n252), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n275), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(G250), .B1(new_n265), .B2(G1), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n268), .A2(G45), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n259), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT83), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT83), .ZN(new_n530));
  INV_X1    g0330(.A(new_n526), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n265), .A2(new_n267), .A3(G1), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n275), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G238), .A2(G1698), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n369), .B2(G1698), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(new_n496), .B1(G33), .B2(G116), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n530), .B(new_n533), .C1(new_n536), .C2(new_n275), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n529), .A2(new_n537), .A3(new_n360), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n358), .B1(new_n529), .B2(new_n537), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT84), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n529), .A2(new_n537), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n388), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT84), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n529), .A2(new_n537), .A3(new_n360), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n496), .A2(new_n212), .A3(G68), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n212), .B1(new_n257), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G87), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(new_n470), .A3(new_n365), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n547), .B1(new_n295), .B2(new_n470), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n546), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n553), .A2(new_n293), .B1(new_n306), .B2(new_n374), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n479), .A2(new_n374), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n540), .A2(new_n545), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n553), .A2(new_n293), .ZN(new_n558));
  INV_X1    g0358(.A(new_n479), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n374), .A2(new_n306), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(G190), .B2(new_n541), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n324), .B2(new_n541), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n557), .A2(KEYINPUT85), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT85), .B1(new_n557), .B2(new_n564), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n306), .A2(new_n470), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n479), .B2(new_n470), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT6), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G97), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n570), .A2(G97), .A3(G107), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT80), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(G107), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n365), .A2(KEYINPUT80), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n572), .A2(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n470), .A2(new_n365), .A3(KEYINPUT6), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n365), .A2(KEYINPUT80), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(G107), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n578), .A2(new_n571), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n212), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n298), .A2(G77), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT81), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT81), .ZN(new_n586));
  AND4_X1   g0386(.A1(new_n578), .A2(new_n571), .A3(new_n579), .A4(new_n580), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n578), .A2(new_n571), .B1(new_n579), .B2(new_n580), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n586), .B(new_n583), .C1(new_n589), .C2(new_n212), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n585), .B(new_n590), .C1(new_n365), .C2(new_n443), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n569), .B1(new_n591), .B2(new_n293), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n249), .A2(G250), .A3(G1698), .A4(new_n254), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n369), .A2(G1698), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(new_n251), .A3(new_n252), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT4), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n595), .A2(KEYINPUT82), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT82), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n596), .A2(new_n369), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n249), .A2(new_n250), .A3(new_n254), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n469), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n259), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(G257), .B(new_n275), .C1(new_n490), .C2(new_n487), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n489), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G200), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(new_n605), .A3(G190), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n592), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n360), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n603), .A2(new_n605), .A3(new_n388), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n609), .B1(new_n592), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(G250), .A2(G1698), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n497), .B2(G1698), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(new_n496), .B1(G33), .B2(G294), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n616), .A2(new_n275), .ZN(new_n617));
  OAI211_X1 g0417(.A(G264), .B(new_n275), .C1(new_n490), .C2(new_n487), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n617), .A2(G179), .A3(new_n489), .A4(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n489), .B(new_n618), .C1(new_n275), .C2(new_n616), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G169), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT90), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT90), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n619), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT22), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n212), .A3(G87), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n395), .A2(G20), .A3(new_n549), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n327), .A2(new_n627), .B1(new_n628), .B2(new_n626), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT23), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(new_n365), .A3(G20), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT88), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n630), .B2(new_n365), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n635));
  OAI22_X1  g0435(.A1(new_n631), .A2(new_n632), .B1(new_n635), .B2(G20), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n629), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT24), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT24), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n629), .A2(new_n640), .A3(new_n637), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n378), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n306), .A2(KEYINPUT25), .A3(new_n365), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT89), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT25), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n312), .B2(G107), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n646), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n647), .A2(new_n648), .B1(G107), .B2(new_n559), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n623), .B(new_n625), .C1(new_n642), .C2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n620), .A2(G200), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n620), .A2(new_n392), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n629), .A2(new_n640), .A3(new_n637), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n640), .B1(new_n629), .B2(new_n637), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n293), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(new_n657), .A3(new_n649), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n613), .A2(new_n659), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n464), .A2(new_n520), .A3(new_n567), .A4(new_n660), .ZN(G372));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n591), .A2(new_n293), .ZN(new_n663));
  INV_X1    g0463(.A(new_n569), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n610), .A3(new_n611), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n662), .B1(new_n567), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n610), .A2(new_n611), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n533), .B1(new_n536), .B2(new_n275), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G200), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n554), .A2(new_n555), .B1(new_n671), .B2(new_n360), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n563), .A2(new_n672), .B1(new_n542), .B2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n670), .A2(new_n662), .A3(new_n665), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n542), .A2(new_n673), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n657), .A2(new_n649), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n622), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n679), .A2(new_n517), .A3(new_n506), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n658), .A2(new_n674), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n666), .A4(new_n609), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n669), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n464), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n439), .A2(new_n449), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n386), .A2(new_n322), .A3(new_n389), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n687), .B1(new_n319), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n413), .A2(new_n436), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n450), .A2(new_n451), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n459), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n691), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT18), .B1(new_n448), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n353), .B1(new_n689), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n686), .A2(new_n362), .A3(new_n696), .ZN(G369));
  AND2_X1   g0497(.A1(new_n517), .A2(new_n506), .ZN(new_n698));
  OR3_X1    g0498(.A1(new_n465), .A2(KEYINPUT27), .A3(G20), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT27), .B1(new_n465), .B2(G20), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n483), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n698), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n520), .B2(new_n704), .ZN(new_n706));
  INV_X1    g0506(.A(G330), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n659), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n678), .A2(new_n703), .ZN(new_n710));
  INV_X1    g0510(.A(new_n651), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n709), .A2(new_n710), .B1(new_n711), .B2(new_n703), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n679), .A2(new_n703), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n698), .A2(new_n703), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(new_n709), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n206), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n484), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n550), .A2(G116), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G1), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n209), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT91), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n703), .B1(new_n669), .B2(new_n684), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT29), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n557), .A2(new_n564), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT85), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n557), .A2(KEYINPUT85), .A3(new_n564), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n732), .A2(new_n662), .A3(new_n733), .A4(new_n667), .ZN(new_n734));
  INV_X1    g0534(.A(new_n676), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n670), .A2(new_n665), .A3(new_n674), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(KEYINPUT26), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT92), .ZN(new_n739));
  INV_X1    g0539(.A(new_n613), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n740), .A2(new_n681), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n698), .A2(new_n651), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n738), .A2(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n734), .A2(KEYINPUT92), .A3(new_n737), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n703), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n729), .B1(new_n745), .B2(new_n728), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n703), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n567), .A2(new_n660), .A3(new_n520), .A4(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n618), .B1(new_n616), .B2(new_n275), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n529), .B2(new_n537), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n509), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n750), .B1(new_n753), .B2(new_n606), .ZN(new_n754));
  INV_X1    g0554(.A(new_n606), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n755), .A2(KEYINPUT30), .A3(new_n509), .A4(new_n752), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n671), .A2(new_n388), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n606), .A2(new_n503), .A3(new_n620), .A4(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n754), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n760));
  AOI21_X1  g0560(.A(KEYINPUT31), .B1(new_n759), .B2(new_n703), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n749), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G330), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n747), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n726), .B1(new_n766), .B2(G1), .ZN(G364));
  AOI21_X1  g0567(.A(new_n211), .B1(G20), .B2(new_n360), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n212), .A2(new_n324), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n358), .A2(G190), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n212), .A2(new_n392), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n358), .A2(new_n324), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G58), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n297), .A2(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR4_X1   g0574(.A1(new_n388), .A2(new_n212), .A3(G190), .A4(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(KEYINPUT93), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n212), .A2(G190), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n358), .A2(new_n324), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT93), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n774), .B1(new_n782), .B2(G77), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G179), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n777), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n407), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT95), .B(KEYINPUT32), .Z(new_n788));
  XNOR2_X1  g0588(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n785), .A2(G190), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n789), .B1(new_n470), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n358), .A2(new_n392), .A3(new_n769), .ZN(new_n794));
  INV_X1    g0594(.A(G68), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n324), .A2(G179), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n777), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G107), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n771), .A2(new_n797), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n328), .B(new_n800), .C1(new_n549), .C2(new_n801), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n784), .A2(new_n793), .A3(new_n796), .A4(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n786), .B(KEYINPUT96), .Z(new_n804));
  INV_X1    g0604(.A(new_n772), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n804), .A2(G329), .B1(G322), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(KEYINPUT33), .B(G317), .Z(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n794), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n801), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G303), .A2(new_n809), .B1(new_n799), .B2(G283), .ZN(new_n810));
  INV_X1    g0610(.A(G294), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n810), .B(new_n327), .C1(new_n811), .C2(new_n792), .ZN(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  INV_X1    g0613(.A(G326), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n813), .A2(new_n778), .B1(new_n770), .B2(new_n814), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n808), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n768), .B1(new_n803), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n305), .A2(G20), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n271), .B1(new_n818), .B2(G45), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n720), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(G13), .A2(G33), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(G20), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n768), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n328), .A2(G355), .A3(new_n206), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(G116), .B2(new_n206), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n719), .A2(new_n496), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(G45), .B2(new_n209), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(new_n242), .B2(G45), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n825), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n817), .A2(new_n821), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n706), .B2(new_n824), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n708), .A2(new_n821), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n706), .A2(new_n707), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  AND4_X1   g0637(.A1(new_n389), .A2(new_n385), .A3(new_n373), .A4(new_n748), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n385), .A2(new_n703), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n391), .B2(new_n393), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n838), .B1(new_n390), .B2(new_n840), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n727), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n748), .C1(new_n668), .C2(new_n683), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n821), .B1(new_n844), .B2(new_n764), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n707), .B1(new_n749), .B2(new_n762), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n842), .A2(new_n846), .A3(new_n843), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n768), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n823), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G107), .A2(new_n809), .B1(new_n799), .B2(G87), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n851), .B(new_n327), .C1(new_n470), .C2(new_n792), .ZN(new_n852));
  INV_X1    g0652(.A(new_n794), .ZN(new_n853));
  INV_X1    g0653(.A(new_n770), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G283), .A2(new_n853), .B1(new_n854), .B2(G303), .ZN(new_n855));
  INV_X1    g0655(.A(new_n804), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n855), .B1(new_n811), .B2(new_n772), .C1(new_n813), .C2(new_n856), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n852), .B(new_n857), .C1(G116), .C2(new_n782), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n801), .A2(new_n297), .B1(new_n798), .B2(new_n795), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n395), .B1(new_n804), .B2(G132), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT97), .Z(new_n861));
  AOI211_X1 g0661(.A(new_n859), .B(new_n861), .C1(G58), .C2(new_n791), .ZN(new_n862));
  AOI22_X1  g0662(.A1(G137), .A2(new_n854), .B1(new_n805), .B2(G143), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n863), .B1(new_n338), .B2(new_n794), .C1(new_n781), .C2(new_n407), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT34), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n858), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n866), .A2(KEYINPUT98), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n768), .B1(new_n866), .B2(KEYINPUT98), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n821), .B1(G77), .B2(new_n850), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n869), .A2(KEYINPUT99), .ZN(new_n870));
  INV_X1    g0670(.A(new_n841), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n822), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(KEYINPUT99), .B2(new_n869), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n848), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  NAND2_X1  g0676(.A1(new_n318), .A2(new_n703), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n319), .A2(new_n322), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n322), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n318), .B(new_n703), .C1(new_n291), .C2(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n838), .B(KEYINPUT100), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n881), .B1(new_n843), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n413), .A2(new_n431), .A3(new_n436), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n448), .B2(new_n701), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n448), .B2(new_n455), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n405), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n397), .B1(new_n496), .B2(G20), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n795), .B1(new_n891), .B2(new_n409), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n445), .B1(new_n408), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n293), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT101), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n890), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n893), .A2(KEYINPUT101), .A3(new_n293), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n435), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT102), .B1(new_n898), .B2(new_n701), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT16), .B1(new_n399), .B2(new_n404), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n895), .B1(new_n900), .B2(new_n378), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n405), .A3(new_n897), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n436), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n903), .A2(new_n691), .B1(new_n448), .B2(new_n431), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT102), .ZN(new_n905));
  INV_X1    g0705(.A(new_n701), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n899), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n889), .B1(new_n908), .B2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n899), .A2(new_n907), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(new_n463), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n884), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n463), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n905), .B1(new_n903), .B2(new_n906), .ZN(new_n914));
  AOI211_X1 g0714(.A(KEYINPUT102), .B(new_n701), .C1(new_n902), .C2(new_n436), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n887), .B1(new_n916), .B2(new_n904), .ZN(new_n917));
  OAI211_X1 g0717(.A(KEYINPUT38), .B(new_n913), .C1(new_n917), .C2(new_n889), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n883), .A2(new_n919), .B1(new_n695), .B2(new_n701), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n319), .A2(new_n703), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n687), .A2(new_n695), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n690), .A2(new_n906), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n923), .B(new_n885), .C1(new_n448), .C2(new_n693), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n889), .B1(KEYINPUT37), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n884), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n927), .A2(new_n918), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT39), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n912), .B2(new_n918), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n921), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n920), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT104), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n920), .A2(new_n932), .A3(KEYINPUT104), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n696), .A2(new_n362), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n746), .B2(new_n464), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n878), .A2(new_n880), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n763), .A2(new_n941), .A3(new_n841), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n919), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT40), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n927), .B2(new_n918), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n943), .A2(new_n944), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n464), .A2(new_n763), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n707), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n947), .B2(new_n946), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n940), .A2(new_n949), .B1(new_n271), .B2(new_n818), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT105), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n940), .A2(new_n949), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n589), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT35), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(KEYINPUT35), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n957), .A2(G116), .A3(new_n213), .A4(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT36), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n210), .A2(G77), .A3(new_n402), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(G50), .B2(new_n795), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(G1), .A3(new_n305), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n955), .A2(new_n960), .A3(new_n963), .ZN(G367));
  INV_X1    g0764(.A(new_n828), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n825), .B1(new_n206), .B2(new_n374), .C1(new_n234), .C2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(G137), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n801), .A2(new_n773), .B1(new_n786), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n791), .A2(G68), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n328), .A2(new_n969), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n968), .B(new_n970), .C1(G77), .C2(new_n799), .ZN(new_n971));
  INV_X1    g0771(.A(G143), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n972), .A2(new_n770), .B1(new_n772), .B2(new_n338), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G159), .B2(new_n853), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n971), .B(new_n974), .C1(new_n297), .C2(new_n781), .ZN(new_n975));
  INV_X1    g0775(.A(G317), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n395), .B1(new_n786), .B2(new_n976), .C1(new_n470), .C2(new_n798), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G107), .B2(new_n791), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G303), .A2(new_n805), .B1(new_n854), .B2(G311), .ZN(new_n979));
  INV_X1    g0779(.A(G283), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n978), .B(new_n979), .C1(new_n980), .C2(new_n781), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n809), .A2(KEYINPUT46), .A3(G116), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT46), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n801), .B2(new_n466), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(new_n811), .C2(new_n794), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT110), .Z(new_n986));
  OAI21_X1  g0786(.A(new_n975), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT47), .Z(new_n988));
  OAI211_X1 g0788(.A(new_n821), .B(new_n966), .C1(new_n988), .C2(new_n849), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT111), .Z(new_n990));
  NAND2_X1  g0790(.A1(new_n562), .A2(new_n703), .ZN(new_n991));
  MUX2_X1   g0791(.A(new_n735), .B(new_n674), .S(new_n991), .Z(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT106), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n824), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT112), .Z(new_n996));
  INV_X1    g0796(.A(KEYINPUT43), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n993), .A2(new_n997), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n740), .B1(new_n592), .B2(new_n748), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n667), .A2(new_n703), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT107), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT107), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1000), .A2(new_n1004), .A3(new_n1001), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT42), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n716), .A2(new_n709), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1007), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1006), .A2(new_n711), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n703), .B1(new_n1014), .B2(new_n666), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n998), .B(new_n999), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n714), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n1006), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1015), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1020), .A2(new_n1021), .A3(new_n997), .A4(new_n993), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1016), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT108), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1016), .A2(KEYINPUT108), .A3(new_n1019), .A4(new_n1022), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n1018), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n720), .B(KEYINPUT41), .Z(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n1000), .A2(new_n1004), .A3(new_n1001), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1004), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n717), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT45), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1006), .A2(KEYINPUT45), .A3(new_n717), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n717), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1003), .A2(new_n1039), .A3(new_n1005), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT44), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1003), .A2(new_n1039), .A3(KEYINPUT44), .A4(new_n1005), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1038), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n1017), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1038), .A2(new_n1044), .A3(new_n714), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n708), .A2(KEYINPUT109), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n716), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1009), .B1(new_n712), .B2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1049), .B(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n747), .A2(new_n1052), .A3(new_n764), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1031), .B1(new_n1054), .B2(new_n765), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n819), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n996), .B1(new_n1029), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(G387));
  OAI22_X1  g0858(.A1(new_n781), .A2(new_n494), .B1(new_n976), .B2(new_n772), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT114), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G311), .A2(new_n853), .B1(new_n854), .B2(G322), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT115), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1064), .B(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT48), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1064), .B(KEYINPUT115), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT48), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n809), .A2(G294), .B1(new_n791), .B2(G283), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1067), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT49), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1067), .A2(new_n1070), .A3(KEYINPUT49), .A4(new_n1071), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n395), .B1(new_n786), .B2(new_n814), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G116), .B2(new_n799), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n395), .B1(new_n799), .B2(G97), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n294), .B2(new_n801), .C1(new_n338), .C2(new_n786), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n792), .A2(new_n374), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n795), .A2(new_n778), .B1(new_n794), .B2(new_n337), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n297), .A2(new_n772), .B1(new_n770), .B2(new_n407), .ZN(new_n1083));
  NOR4_X1   g0883(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n849), .B1(new_n1078), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT116), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n825), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n722), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n328), .A2(new_n206), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(G107), .B2(new_n206), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n231), .A2(G45), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT113), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n376), .A2(new_n297), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT50), .Z(new_n1095));
  AOI211_X1 g0895(.A(G45), .B(new_n1089), .C1(G68), .C2(G77), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n965), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1091), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n824), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n821), .B1(new_n1088), .B2(new_n1098), .C1(new_n713), .C2(new_n1099), .ZN(new_n1100));
  OR3_X1    g0900(.A1(new_n1086), .A2(new_n1087), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1087), .B1(new_n1086), .B2(new_n1100), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1101), .A2(new_n1102), .B1(new_n820), .B2(new_n1052), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1053), .A2(KEYINPUT117), .A3(new_n720), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1052), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n765), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT117), .B1(new_n1053), .B2(new_n720), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1103), .B1(new_n1107), .B2(new_n1108), .ZN(G393));
  AOI22_X1  g0909(.A1(new_n1037), .A2(new_n1036), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1110));
  OAI21_X1  g0910(.A(KEYINPUT119), .B1(new_n1110), .B2(new_n714), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT119), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1045), .A2(new_n1112), .A3(new_n1017), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT118), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1047), .B(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1114), .A2(new_n1116), .A3(new_n820), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n239), .A2(new_n828), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n825), .B1(new_n470), .B2(new_n206), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n821), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n792), .A2(new_n294), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n395), .B1(new_n799), .B2(G87), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n972), .B2(new_n786), .C1(new_n216), .C2(new_n801), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1121), .B(new_n1123), .C1(G50), .C2(new_n853), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n338), .A2(new_n770), .B1(new_n772), .B2(new_n407), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT51), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n782), .A2(new_n376), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT120), .ZN(new_n1129));
  INV_X1    g0929(.A(G322), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n800), .B1(new_n980), .B2(new_n801), .C1(new_n1130), .C2(new_n786), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n328), .B(new_n1131), .C1(G116), .C2(new_n791), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n813), .A2(new_n772), .B1(new_n770), .B2(new_n976), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT52), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n853), .A2(G303), .B1(new_n775), .B2(G294), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1129), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT121), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1120), .B1(new_n1138), .B2(new_n768), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1099), .B2(new_n1006), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1114), .A2(new_n1116), .B1(new_n766), .B2(new_n1052), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n720), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1117), .B(new_n1140), .C1(new_n1141), .C2(new_n1142), .ZN(G390));
  NOR3_X1   g0943(.A1(new_n764), .A2(new_n881), .A3(new_n871), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n927), .A2(new_n918), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n319), .B2(new_n703), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n738), .A2(new_n739), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n741), .A2(new_n742), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(new_n744), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n748), .A3(new_n841), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n882), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1146), .B1(new_n1151), .B2(new_n941), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n889), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT38), .B1(new_n1155), .B2(new_n913), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n909), .A2(new_n911), .A3(new_n884), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT39), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n927), .A2(new_n918), .A3(new_n928), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n843), .A2(new_n882), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n921), .B1(new_n1161), .B2(new_n941), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1144), .B1(new_n1152), .B2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1158), .B(new_n1159), .C1(new_n883), .C2(new_n921), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1144), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n881), .B1(new_n1150), .B2(new_n882), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1165), .B(new_n1166), .C1(new_n1167), .C2(new_n1146), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n464), .A2(new_n846), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n938), .B(new_n1170), .C1(new_n746), .C2(new_n464), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n941), .B1(new_n846), .B2(new_n841), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1144), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n882), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n745), .B2(new_n841), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1161), .B1(new_n1144), .B2(new_n1172), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1171), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1169), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1164), .A2(new_n1168), .A3(new_n1171), .A4(new_n1178), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n720), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1164), .A2(new_n820), .A3(new_n1168), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n821), .B1(new_n433), .B2(new_n850), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n770), .A2(new_n980), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n365), .A2(new_n794), .B1(new_n772), .B2(new_n466), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(G294), .C2(new_n804), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n801), .A2(new_n549), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n798), .A2(new_n795), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n328), .A2(new_n1121), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1187), .B(new_n1190), .C1(new_n470), .C2(new_n781), .ZN(new_n1191));
  INV_X1    g0991(.A(G125), .ZN(new_n1192));
  INV_X1    g0992(.A(G132), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n856), .A2(new_n1192), .B1(new_n1193), .B2(new_n772), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G137), .B2(new_n853), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n809), .A2(G150), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT53), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G159), .B2(new_n791), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n328), .B1(new_n297), .B2(new_n798), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G128), .B2(new_n854), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1195), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT54), .B(G143), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n781), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1191), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1184), .B1(new_n1204), .B2(new_n768), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1160), .B2(new_n823), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1182), .A2(new_n1183), .A3(new_n1206), .ZN(G378));
  NAND2_X1  g1007(.A1(new_n1181), .A2(new_n1171), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT125), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n354), .A2(new_n701), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n363), .A2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n353), .B(new_n362), .C1(new_n354), .C2(new_n701), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1213), .B(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n946), .B2(G330), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n912), .A2(new_n918), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n763), .A2(new_n941), .A3(new_n841), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n944), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n945), .A2(new_n942), .ZN(new_n1221));
  AND4_X1   g1021(.A1(G330), .A2(new_n1220), .A3(new_n1221), .A4(new_n1216), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n935), .B(new_n936), .C1(new_n1217), .C2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1220), .A2(G330), .A3(new_n1221), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1216), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n946), .A2(G330), .A3(new_n1216), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n920), .A2(new_n932), .A3(KEYINPUT104), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT104), .B1(new_n920), .B2(new_n932), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1226), .B(new_n1227), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1209), .B1(new_n1223), .B2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1217), .A2(new_n1222), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT125), .B1(new_n1232), .B2(new_n937), .ZN(new_n1233));
  OAI211_X1 g1033(.A(KEYINPUT57), .B(new_n1208), .C1(new_n1231), .C2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1223), .A2(new_n1230), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1208), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT57), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1234), .A2(new_n1238), .A3(new_n720), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1225), .A2(new_n822), .ZN(new_n1240));
  AOI211_X1 g1040(.A(G33), .B(G41), .C1(new_n799), .C2(G159), .ZN(new_n1241));
  INV_X1    g1041(.A(G124), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n770), .A2(new_n1192), .B1(new_n792), .B2(new_n338), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n1193), .A2(new_n794), .B1(new_n778), .B2(new_n967), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1202), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n805), .A2(G128), .B1(new_n809), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1247), .A2(KEYINPUT122), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(KEYINPUT122), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1243), .B(new_n1244), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT59), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1241), .B1(new_n1242), .B2(new_n786), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1251), .B2(new_n1250), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(G97), .A2(new_n853), .B1(new_n805), .B2(G107), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n374), .B2(new_n778), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n856), .A2(new_n980), .B1(new_n466), .B2(new_n770), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n496), .B(new_n484), .C1(new_n809), .C2(G77), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n799), .A2(G58), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n969), .A3(new_n1258), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1255), .A2(new_n1256), .A3(new_n1259), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1260), .A2(KEYINPUT58), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(KEYINPUT58), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n297), .B1(G33), .B2(G41), .C1(new_n484), .C2(new_n496), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n768), .B1(new_n1253), .B2(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT123), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n821), .B1(G50), .B2(new_n850), .ZN(new_n1267));
  XOR2_X1   g1067(.A(new_n1267), .B(KEYINPUT124), .Z(new_n1268));
  NOR2_X1   g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1235), .A2(new_n820), .B1(new_n1240), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1239), .A2(new_n1270), .ZN(G375));
  NAND2_X1  g1071(.A1(new_n881), .A2(new_n822), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n821), .B1(G68), .B2(new_n850), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n770), .A2(new_n811), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n466), .A2(new_n794), .B1(new_n772), .B2(new_n980), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n1274), .B(new_n1275), .C1(G303), .C2(new_n804), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n801), .A2(new_n470), .B1(new_n798), .B2(new_n294), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n328), .A2(new_n1081), .A3(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1276), .B(new_n1278), .C1(new_n365), .C2(new_n781), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n801), .A2(new_n407), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1258), .A2(new_n496), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1280), .B(new_n1281), .C1(G50), .C2(new_n791), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n854), .A2(G132), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n853), .A2(new_n1245), .B1(new_n775), .B2(G150), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n804), .A2(G128), .B1(G137), .B2(new_n805), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1279), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1273), .B1(new_n1287), .B2(new_n768), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n1178), .A2(new_n820), .B1(new_n1272), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1179), .A2(new_n1031), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1178), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1170), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n939), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1290), .B1(new_n1292), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(G381));
  NOR3_X1   g1098(.A1(G381), .A2(G390), .A3(G384), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n836), .B(new_n1103), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1057), .A3(new_n1301), .ZN(new_n1302));
  OR3_X1    g1102(.A1(new_n1302), .A2(G378), .A3(G375), .ZN(G407));
  INV_X1    g1103(.A(G378), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n702), .A2(G213), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G407), .B(G213), .C1(G375), .C2(new_n1307), .ZN(G409));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1239), .A2(G378), .A3(new_n1270), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n820), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1240), .A2(new_n1269), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1236), .A2(new_n1030), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1304), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1310), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1305), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1293), .A2(KEYINPUT60), .A3(new_n1295), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1318), .A2(new_n720), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1179), .A2(KEYINPUT60), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1296), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G384), .B1(new_n1322), .B2(new_n1289), .ZN(new_n1323));
  AOI211_X1 g1123(.A(new_n1290), .B(new_n875), .C1(new_n1319), .C2(new_n1321), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1309), .B1(new_n1317), .B2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(G2897), .B(new_n1306), .C1(new_n1323), .C2(new_n1324), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1322), .A2(new_n1289), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n875), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1322), .A2(G384), .A3(new_n1289), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1306), .A2(G2897), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1330), .A2(new_n1331), .A3(new_n1332), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1328), .A2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT61), .B1(new_n1317), .B2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(G393), .A2(G396), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1300), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT118), .B1(new_n1110), .B2(new_n714), .ZN(new_n1338));
  AND4_X1   g1138(.A1(KEYINPUT118), .A2(new_n1038), .A3(new_n1044), .A4(new_n714), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1111), .B(new_n1113), .C1(new_n1338), .C2(new_n1339), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1140), .B1(new_n1340), .B2(new_n819), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1053), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1142), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1341), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1337), .A2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(G390), .A2(new_n1336), .A3(new_n1300), .ZN(new_n1346));
  AND3_X1   g1146(.A1(new_n1345), .A2(new_n1057), .A3(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1057), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1306), .B1(new_n1310), .B2(new_n1315), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1350), .A2(KEYINPUT63), .A3(new_n1325), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1327), .A2(new_n1335), .A3(new_n1349), .A4(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT62), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1350), .A2(new_n1353), .A3(new_n1325), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT61), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1328), .A2(new_n1333), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1355), .B1(new_n1350), .B2(new_n1356), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1353), .B1(new_n1350), .B2(new_n1325), .ZN(new_n1358));
  NOR3_X1   g1158(.A1(new_n1354), .A2(new_n1357), .A3(new_n1358), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1352), .B1(new_n1359), .B2(new_n1349), .ZN(G405));
  NAND2_X1  g1160(.A1(G375), .A2(new_n1304), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1310), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1326), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1364), .A2(G387), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1345), .A2(new_n1057), .A3(new_n1346), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1365), .A2(new_n1325), .A3(new_n1366), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT126), .ZN(new_n1368));
  AND3_X1   g1168(.A1(new_n1363), .A2(new_n1367), .A3(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1368), .B1(new_n1363), .B2(new_n1367), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n1362), .B1(new_n1369), .B2(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1363), .A2(new_n1367), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1372), .A2(KEYINPUT126), .ZN(new_n1373));
  INV_X1    g1173(.A(new_n1362), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1363), .A2(new_n1367), .A3(new_n1368), .ZN(new_n1375));
  NAND3_X1  g1175(.A1(new_n1373), .A2(new_n1374), .A3(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1371), .A2(new_n1376), .ZN(G402));
endmodule


