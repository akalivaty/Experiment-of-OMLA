//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979;
  OR2_X1    g000(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n203));
  AOI21_X1  g002(.A(G36gat), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  AND3_X1   g004(.A1(new_n205), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n204), .A2(KEYINPUT15), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G43gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G50gat), .ZN(new_n209));
  INV_X1    g008(.A(G50gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G43gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT87), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(new_n204), .B2(new_n206), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n207), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n217), .A2(new_n212), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT17), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT88), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(G1gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n225), .B2(G1gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n226), .A3(KEYINPUT89), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n227), .B(G8gat), .C1(KEYINPUT89), .C2(new_n226), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n226), .A2(KEYINPUT90), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(KEYINPUT90), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n224), .A4(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n219), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT17), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n222), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT91), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n233), .A2(new_n234), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n233), .B(new_n234), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n238), .B(KEYINPUT13), .Z(new_n244));
  AOI22_X1  g043(.A1(new_n240), .A2(new_n241), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G141gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(G169gat), .B(G197gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT12), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n246), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n242), .A2(new_n245), .A3(new_n252), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G8gat), .B(G36gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(G64gat), .B(G92gat), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n258), .B(new_n259), .Z(new_n260));
  XNOR2_X1  g059(.A(G197gat), .B(G204gat), .ZN(new_n261));
  INV_X1    g060(.A(G211gat), .ZN(new_n262));
  INV_X1    g061(.A(G218gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n261), .B1(KEYINPUT22), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G226gat), .ZN(new_n269));
  INV_X1    g068(.A(G233gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT27), .B(G183gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(KEYINPUT67), .ZN(new_n276));
  AOI21_X1  g075(.A(G190gat), .B1(new_n275), .B2(KEYINPUT67), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n276), .B1(new_n274), .B2(new_n277), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n273), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT26), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G169gat), .ZN(new_n284));
  INV_X1    g083(.A(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n284), .A3(new_n285), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n282), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT68), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n289), .A2(new_n293), .A3(new_n282), .A4(new_n290), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n287), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n297), .A2(G169gat), .A3(G176gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n281), .A2(KEYINPUT23), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n286), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n273), .ZN(new_n302));
  NAND4_X1  g101(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT65), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n296), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n302), .A2(new_n304), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(new_n299), .B2(new_n286), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n289), .A2(KEYINPUT23), .A3(new_n290), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  OAI22_X1  g112(.A1(new_n280), .A2(new_n295), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n292), .A2(new_n294), .ZN(new_n317));
  INV_X1    g116(.A(new_n287), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n273), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n274), .A2(new_n277), .ZN(new_n321));
  INV_X1    g120(.A(new_n276), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n320), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n300), .A2(new_n307), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(new_n296), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(KEYINPUT73), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n272), .B1(new_n316), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n271), .A2(KEYINPUT29), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n268), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n316), .A2(new_n330), .A3(new_n332), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n326), .A2(new_n329), .A3(new_n271), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(new_n267), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n260), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n338), .A3(new_n260), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT30), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n335), .A2(new_n338), .ZN(new_n343));
  INV_X1    g142(.A(new_n260), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n343), .A2(KEYINPUT30), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT5), .ZN(new_n348));
  XOR2_X1   g147(.A(G127gat), .B(G134gat), .Z(new_n349));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n350));
  INV_X1    g149(.A(G120gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G113gat), .ZN(new_n352));
  INV_X1    g151(.A(G113gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G120gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n350), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI211_X1 g156(.A(KEYINPUT70), .B(KEYINPUT1), .C1(new_n352), .C2(new_n354), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n349), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OR2_X1    g158(.A1(G141gat), .A2(G148gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(KEYINPUT75), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n363));
  AND2_X1   g162(.A1(G141gat), .A2(G148gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT2), .ZN(new_n368));
  INV_X1    g167(.A(G155gat), .ZN(new_n369));
  INV_X1    g168(.A(G162gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(new_n369), .B2(new_n370), .ZN(new_n372));
  AND2_X1   g171(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n373));
  NOR2_X1   g172(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n360), .B(new_n361), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G155gat), .B(G162gat), .Z(new_n376));
  AOI22_X1  g175(.A1(new_n367), .A2(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT69), .B1(new_n378), .B2(KEYINPUT1), .ZN(new_n379));
  INV_X1    g178(.A(new_n349), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT70), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n353), .A2(G120gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n351), .A2(G113gat), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n381), .B(new_n356), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n359), .A2(new_n377), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT77), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n359), .A2(new_n377), .A3(new_n388), .A4(new_n385), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n359), .A2(new_n385), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n364), .A2(new_n365), .A3(new_n363), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT75), .B1(new_n360), .B2(new_n361), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n372), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n376), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n387), .A2(new_n389), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G225gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n348), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n387), .A2(new_n401), .A3(new_n389), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n393), .A2(new_n403), .A3(new_n394), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT76), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n377), .A2(KEYINPUT76), .A3(new_n403), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(KEYINPUT3), .A2(new_n395), .B1(new_n359), .B2(new_n385), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n380), .B1(new_n379), .B2(new_n384), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(KEYINPUT4), .A3(new_n377), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n402), .A2(new_n410), .A3(new_n398), .A4(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n400), .A2(new_n415), .ZN(new_n416));
  AOI211_X1 g215(.A(KEYINPUT5), .B(new_n399), .C1(new_n408), .C2(new_n409), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n387), .A2(KEYINPUT4), .A3(new_n389), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n359), .A2(new_n377), .A3(new_n401), .A4(new_n385), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n419), .A2(KEYINPUT79), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT79), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n387), .A2(new_n422), .A3(KEYINPUT4), .A4(new_n389), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n417), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT80), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n417), .A2(new_n421), .A3(KEYINPUT80), .A4(new_n423), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n416), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  XOR2_X1   g228(.A(G1gat), .B(G29gat), .Z(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G57gat), .B(G85gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n428), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n435), .A2(new_n429), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n434), .A2(KEYINPUT6), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n428), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n347), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT81), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n427), .ZN(new_n444));
  INV_X1    g243(.A(new_n416), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n438), .ZN(new_n447));
  INV_X1    g246(.A(new_n439), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n436), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(KEYINPUT81), .A3(new_n347), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n403), .B1(new_n267), .B2(KEYINPUT29), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n395), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT29), .B1(new_n406), .B2(new_n407), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(new_n268), .ZN(new_n455));
  INV_X1    g254(.A(G228gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(new_n270), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n453), .B(new_n457), .C1(new_n454), .C2(new_n268), .ZN(new_n460));
  INV_X1    g259(.A(G22gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G78gat), .B(G106gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT31), .B(G50gat), .ZN(new_n464));
  XOR2_X1   g263(.A(new_n463), .B(new_n464), .Z(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n461), .B1(new_n459), .B2(new_n460), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n467), .B1(KEYINPUT83), .B2(new_n469), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n469), .A2(KEYINPUT83), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(KEYINPUT82), .A3(new_n462), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n459), .A2(new_n460), .A3(new_n473), .A4(new_n461), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n474), .A2(new_n465), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n470), .A2(new_n471), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n314), .A2(new_n390), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n326), .A2(new_n413), .A3(new_n329), .ZN(new_n478));
  NAND2_X1  g277(.A1(G227gat), .A2(G233gat), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT34), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT34), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n477), .A2(new_n478), .A3(new_n482), .A4(new_n479), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT71), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT71), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(new_n486), .A3(new_n483), .ZN(new_n487));
  XOR2_X1   g286(.A(G15gat), .B(G43gat), .Z(new_n488));
  XNOR2_X1  g287(.A(G71gat), .B(G99gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n479), .B1(new_n477), .B2(new_n478), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(KEYINPUT33), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT32), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n478), .ZN(new_n496));
  INV_X1    g295(.A(new_n479), .ZN(new_n497));
  AOI221_X4 g296(.A(new_n493), .B1(KEYINPUT33), .B2(new_n490), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n485), .B(new_n487), .C1(new_n495), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT72), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n487), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n486), .B1(new_n481), .B2(new_n483), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n496), .A2(new_n497), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT32), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT33), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n508), .A3(new_n490), .ZN(new_n509));
  INV_X1    g308(.A(new_n498), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n504), .A2(new_n511), .A3(KEYINPUT72), .ZN(new_n512));
  INV_X1    g311(.A(new_n484), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n501), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n476), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n443), .A2(new_n451), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT35), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n470), .A2(new_n471), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n472), .A2(new_n475), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n484), .B1(new_n495), .B2(new_n498), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n514), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(KEYINPUT35), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n450), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT84), .ZN(new_n527));
  INV_X1    g326(.A(new_n341), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n528), .A2(new_n339), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n527), .B1(new_n530), .B2(new_n345), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n342), .A2(new_n346), .A3(KEYINPUT84), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n534), .ZN(new_n535));
  AOI221_X4 g334(.A(new_n442), .B1(new_n342), .B2(new_n346), .C1(new_n449), .C2(new_n436), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT81), .B1(new_n450), .B2(new_n347), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n476), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n344), .B1(new_n343), .B2(KEYINPUT37), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n267), .B1(new_n331), .B2(new_n334), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n336), .A2(new_n268), .A3(new_n337), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(KEYINPUT37), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT38), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(new_n528), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n343), .A2(KEYINPUT37), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT38), .B1(new_n547), .B2(new_n539), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n546), .A2(new_n436), .A3(new_n449), .A4(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT39), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n421), .A2(new_n423), .A3(new_n410), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(KEYINPUT85), .A3(new_n399), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT85), .B1(new_n551), .B2(new_n399), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n551), .A2(new_n399), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT85), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n397), .A2(new_n399), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(new_n550), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n552), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n555), .A2(new_n561), .A3(new_n434), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT40), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n555), .A2(new_n561), .A3(KEYINPUT40), .A4(new_n434), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n446), .A2(new_n435), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n531), .A2(new_n567), .A3(new_n532), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n521), .B(new_n549), .C1(new_n566), .C2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n514), .B1(new_n499), .B2(new_n500), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT72), .B1(new_n504), .B2(new_n511), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT36), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n523), .A2(KEYINPUT36), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n538), .A2(new_n569), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n257), .B1(new_n535), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n578), .A2(KEYINPUT92), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(KEYINPUT92), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT21), .ZN(new_n583));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G71gat), .B(G78gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  OAI21_X1  g387(.A(new_n233), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT94), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n583), .ZN(new_n593));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n596), .B(KEYINPUT20), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n595), .B(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G183gat), .B(G211gat), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n598), .A2(new_n600), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n592), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  INV_X1    g404(.A(new_n591), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n590), .B(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n607), .A3(new_n601), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT7), .ZN(new_n612));
  NOR2_X1   g411(.A1(G85gat), .A2(G92gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(KEYINPUT8), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT95), .ZN(new_n616));
  XNOR2_X1  g415(.A(G99gat), .B(G106gat), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n612), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n616), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n222), .A2(new_n235), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G190gat), .B(G218gat), .Z(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n234), .ZN(new_n624));
  INV_X1    g423(.A(new_n620), .ZN(new_n625));
  AND2_X1   g424(.A1(G232gat), .A2(G233gat), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n624), .A2(new_n625), .B1(KEYINPUT41), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n621), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n623), .B1(new_n621), .B2(new_n627), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n626), .A2(KEYINPUT41), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n631), .A2(new_n634), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n620), .A2(new_n588), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT96), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n620), .A2(new_n588), .ZN(new_n644));
  OAI211_X1 g443(.A(KEYINPUT96), .B(KEYINPUT10), .C1(new_n620), .C2(new_n588), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n643), .ZN(new_n647));
  INV_X1    g446(.A(new_n644), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(new_n640), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  NAND3_X1  g451(.A1(new_n646), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n646), .A2(new_n649), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n658), .A2(new_n652), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n610), .A2(new_n638), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT98), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n450), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n449), .A2(KEYINPUT98), .A3(new_n436), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n582), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g468(.A1(new_n662), .A2(new_n533), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  AND3_X1   g470(.A1(new_n582), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n230), .B1(new_n582), .B2(new_n670), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT42), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(KEYINPUT42), .B2(new_n672), .ZN(G1325gat));
  NAND2_X1  g474(.A1(new_n582), .A2(new_n663), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n575), .A2(KEYINPUT99), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n572), .A2(new_n574), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n523), .A2(G15gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n676), .B2(new_n682), .ZN(G1326gat));
  NOR2_X1   g482(.A1(new_n676), .A2(new_n521), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n684), .B(new_n685), .Z(G1327gat));
  NAND2_X1  g485(.A1(new_n609), .A2(new_n661), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n638), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n582), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n667), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n689), .A2(G29gat), .A3(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(KEYINPUT45), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n680), .A2(new_n538), .A3(new_n569), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n535), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n636), .A2(new_n637), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n535), .A2(new_n577), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n638), .A2(new_n697), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n696), .A2(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n687), .A2(new_n257), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(new_n667), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT100), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n205), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n703), .B2(new_n702), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n691), .A2(KEYINPUT45), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n692), .A2(new_n705), .A3(new_n706), .ZN(G1328gat));
  NOR3_X1   g506(.A1(new_n581), .A2(new_n638), .A3(new_n687), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n533), .A2(G36gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT101), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n709), .B1(new_n708), .B2(new_n710), .ZN(new_n713));
  INV_X1    g512(.A(new_n533), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n700), .A2(new_n714), .A3(new_n701), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(G36gat), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n712), .A2(new_n716), .ZN(G1329gat));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n523), .A2(G43gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n582), .A2(new_n688), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n700), .A2(new_n701), .ZN(new_n721));
  OAI21_X1  g520(.A(G43gat), .B1(new_n721), .B2(new_n680), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n718), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1330gat));
  OAI21_X1  g524(.A(G50gat), .B1(new_n721), .B2(new_n521), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n476), .A2(new_n210), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n689), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT48), .Z(G1331gat));
  NOR2_X1   g528(.A1(new_n695), .A2(new_n609), .ZN(new_n730));
  AND4_X1   g529(.A1(new_n257), .A2(new_n694), .A3(new_n730), .A4(new_n660), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n667), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g532(.A(new_n533), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT103), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1333gat));
  INV_X1    g537(.A(new_n680), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n731), .A2(G71gat), .A3(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n523), .B(KEYINPUT104), .Z(new_n741));
  AND2_X1   g540(.A1(new_n731), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n742), .B2(G71gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n731), .A2(new_n476), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  AND3_X1   g545(.A1(new_n538), .A2(new_n569), .A3(new_n576), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n517), .A2(KEYINPUT35), .B1(new_n533), .B2(new_n526), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n699), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n610), .A2(new_n256), .A3(new_n661), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n638), .B1(new_n535), .B2(new_n693), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(KEYINPUT44), .ZN(new_n752));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n690), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n610), .A2(new_n256), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n694), .A2(KEYINPUT51), .A3(new_n695), .A4(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n694), .A2(new_n695), .A3(new_n754), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n751), .A2(KEYINPUT105), .A3(KEYINPUT51), .A4(new_n754), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n757), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  OR3_X1    g561(.A1(new_n690), .A2(G85gat), .A3(new_n661), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n753), .B1(new_n762), .B2(new_n763), .ZN(G1336gat));
  NAND3_X1  g563(.A1(new_n757), .A2(new_n760), .A3(new_n761), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n533), .A2(new_n661), .A3(G92gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  OAI21_X1  g567(.A(G92gat), .B1(new_n752), .B2(new_n533), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(KEYINPUT107), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(KEYINPUT107), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n759), .A2(KEYINPUT106), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n751), .A2(new_n754), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n751), .B2(new_n754), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n766), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n776), .A2(new_n769), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n771), .A2(new_n772), .B1(new_n768), .B2(new_n777), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n752), .B2(new_n680), .ZN(new_n779));
  OR3_X1    g578(.A1(new_n661), .A2(G99gat), .A3(new_n523), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n762), .B2(new_n780), .ZN(G1338gat));
  NOR3_X1   g580(.A1(new_n661), .A2(new_n521), .A3(G106gat), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n765), .A2(KEYINPUT109), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT109), .B1(new_n765), .B2(new_n782), .ZN(new_n784));
  OAI21_X1  g583(.A(G106gat), .B1(new_n752), .B2(new_n521), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n783), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n789), .B(G106gat), .C1(new_n752), .C2(new_n521), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n782), .B1(new_n774), .B2(new_n775), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n785), .A2(KEYINPUT108), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n786), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT110), .B1(new_n788), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n796));
  INV_X1    g595(.A(new_n782), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n762), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n765), .A2(KEYINPUT109), .A3(new_n782), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n798), .A2(new_n786), .A3(new_n785), .A4(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n793), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n790), .A2(new_n791), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT53), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n800), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n795), .A2(new_n805), .ZN(G1339gat));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n662), .B2(new_n256), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n730), .A2(new_n257), .A3(KEYINPUT111), .A4(new_n661), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n646), .A2(KEYINPUT54), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n652), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n647), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(KEYINPUT54), .A3(new_n646), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n695), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n238), .B1(new_n236), .B2(new_n239), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n243), .A2(new_n244), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n251), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n255), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n816), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n824), .A2(KEYINPUT55), .B1(new_n656), .B2(new_n655), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n819), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n256), .A2(new_n825), .A3(new_n818), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n823), .A2(new_n660), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n695), .B1(new_n830), .B2(KEYINPUT112), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n828), .A2(new_n832), .A3(new_n829), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n827), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n810), .B1(new_n834), .B2(new_n610), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(new_n521), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n667), .A2(new_n533), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n523), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n839), .A2(new_n353), .A3(new_n257), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n835), .A2(new_n516), .A3(new_n667), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n714), .ZN(new_n842));
  AOI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n256), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n840), .A2(new_n843), .ZN(G1340gat));
  NOR3_X1   g643(.A1(new_n839), .A2(new_n351), .A3(new_n661), .ZN(new_n845));
  AOI21_X1  g644(.A(G120gat), .B1(new_n842), .B2(new_n660), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(G1341gat));
  OAI21_X1  g646(.A(G127gat), .B1(new_n839), .B2(new_n609), .ZN(new_n848));
  INV_X1    g647(.A(G127gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n842), .A2(new_n849), .A3(new_n610), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(G1342gat));
  OAI21_X1  g650(.A(G134gat), .B1(new_n839), .B2(new_n638), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT113), .ZN(new_n853));
  NOR4_X1   g652(.A1(new_n841), .A2(G134gat), .A3(new_n714), .A4(new_n638), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT56), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(G1343gat));
  AND2_X1   g655(.A1(new_n808), .A2(new_n809), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n660), .A2(new_n255), .A3(new_n822), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n657), .B1(new_n817), .B2(new_n816), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n254), .B2(new_n255), .ZN(new_n861));
  XNOR2_X1  g660(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n816), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n858), .B1(new_n864), .B2(new_n695), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n256), .A2(new_n825), .A3(new_n863), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n829), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(KEYINPUT115), .A3(new_n638), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n868), .A3(new_n826), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n857), .B1(new_n869), .B2(new_n609), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT57), .B1(new_n870), .B2(new_n521), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n831), .A2(new_n833), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n610), .B1(new_n873), .B2(new_n826), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n872), .B(new_n476), .C1(new_n874), .C2(new_n857), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n739), .A2(new_n837), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n871), .A2(new_n256), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT58), .B1(new_n877), .B2(G141gat), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n680), .A2(new_n476), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT117), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n835), .A2(new_n880), .A3(new_n667), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n835), .A2(new_n880), .A3(KEYINPUT118), .A4(new_n667), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n533), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n257), .A2(G141gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n878), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n877), .A2(KEYINPUT116), .A3(G141gat), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT116), .B1(new_n877), .B2(G141gat), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n881), .A2(new_n714), .A3(new_n887), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT58), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(G1344gat));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  OAI211_X1 g694(.A(KEYINPUT57), .B(new_n476), .C1(new_n874), .C2(new_n857), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n826), .B1(new_n864), .B2(new_n695), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n899), .A2(new_n609), .B1(new_n257), .B2(new_n663), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n872), .B1(new_n900), .B2(new_n521), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n897), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n660), .B(new_n876), .C1(new_n898), .C2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n895), .B1(new_n903), .B2(G148gat), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n871), .A2(new_n660), .A3(new_n875), .A4(new_n876), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n906));
  INV_X1    g705(.A(G148gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(KEYINPUT59), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n906), .B1(new_n905), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n660), .A2(new_n907), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n904), .A2(new_n911), .B1(new_n886), .B2(new_n912), .ZN(G1345gat));
  NAND3_X1  g712(.A1(new_n871), .A2(new_n875), .A3(new_n876), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n914), .A2(new_n369), .A3(new_n609), .ZN(new_n915));
  AND4_X1   g714(.A1(new_n533), .A2(new_n883), .A3(new_n610), .A4(new_n884), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(G155gat), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(G1346gat));
  NAND4_X1  g719(.A1(new_n885), .A2(new_n370), .A3(new_n533), .A4(new_n695), .ZN(new_n921));
  OAI21_X1  g720(.A(G162gat), .B1(new_n914), .B2(new_n638), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1347gat));
  NAND3_X1  g722(.A1(new_n690), .A2(new_n714), .A3(new_n741), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT122), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n836), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n926), .A2(new_n284), .A3(new_n257), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n835), .A2(new_n690), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n533), .A2(new_n515), .A3(new_n476), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n256), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n927), .B1(new_n284), .B2(new_n930), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n926), .B2(new_n661), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n660), .A2(new_n285), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(G1349gat));
  NOR2_X1   g734(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n936));
  AND2_X1   g735(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n937));
  OAI21_X1  g736(.A(G183gat), .B1(new_n926), .B2(new_n609), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n928), .A2(new_n274), .A3(new_n610), .A4(new_n929), .ZN(new_n939));
  AOI211_X1 g738(.A(new_n936), .B(new_n937), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  AND4_X1   g739(.A1(KEYINPUT123), .A2(new_n938), .A3(KEYINPUT60), .A4(new_n939), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(G1350gat));
  OR3_X1    g741(.A1(new_n933), .A2(G190gat), .A3(new_n638), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n835), .A2(new_n521), .A3(new_n695), .A4(new_n925), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G190gat), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n945), .A2(KEYINPUT124), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(KEYINPUT124), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n947), .B1(new_n946), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(G1351gat));
  NAND3_X1  g750(.A1(new_n680), .A2(new_n476), .A3(new_n714), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n928), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g753(.A(KEYINPUT125), .B(G197gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(new_n256), .A3(new_n955), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n898), .A2(new_n902), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n680), .A2(new_n714), .A3(new_n690), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT126), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n957), .A2(new_n256), .A3(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n956), .B1(new_n961), .B2(new_n955), .ZN(G1352gat));
  NAND3_X1  g761(.A1(new_n957), .A2(new_n660), .A3(new_n959), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G204gat), .ZN(new_n964));
  INV_X1    g763(.A(G204gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n954), .A2(new_n965), .A3(new_n660), .ZN(new_n966));
  AND2_X1   g765(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n966), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n964), .A2(new_n968), .A3(new_n970), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n262), .A3(new_n610), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n610), .B(new_n959), .C1(new_n898), .C2(new_n902), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  NAND3_X1  g775(.A1(new_n954), .A2(new_n263), .A3(new_n695), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n957), .A2(new_n695), .A3(new_n959), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n977), .B1(new_n979), .B2(new_n263), .ZN(G1355gat));
endmodule


