

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U556 ( .A1(n527), .A2(n528), .ZN(n885) );
  AND2_X1 U557 ( .A1(n788), .A2(n1012), .ZN(n789) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n727) );
  INV_X1 U559 ( .A(n771), .ZN(n754) );
  INV_X1 U560 ( .A(KEYINPUT28), .ZN(n732) );
  OR2_X1 U561 ( .A1(n770), .A2(n779), .ZN(n776) );
  INV_X1 U562 ( .A(n805), .ZN(n788) );
  NAND2_X1 U563 ( .A1(n728), .A2(n727), .ZN(n771) );
  NAND2_X1 U564 ( .A1(n790), .A2(n789), .ZN(n792) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  NOR2_X1 U566 ( .A1(G651), .A2(n642), .ZN(n662) );
  NOR2_X2 U567 ( .A1(G2105), .A2(n527), .ZN(n881) );
  NOR2_X2 U568 ( .A1(n528), .A2(G2104), .ZN(n886) );
  INV_X1 U569 ( .A(KEYINPUT89), .ZN(n538) );
  XOR2_X1 U570 ( .A(KEYINPUT17), .B(n523), .Z(n882) );
  NAND2_X1 U571 ( .A1(n882), .A2(G137), .ZN(n526) );
  INV_X1 U572 ( .A(G2104), .ZN(n527) );
  NAND2_X1 U573 ( .A1(G101), .A2(n881), .ZN(n524) );
  XOR2_X1 U574 ( .A(KEYINPUT23), .B(n524), .Z(n525) );
  NAND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n532) );
  INV_X1 U576 ( .A(G2105), .ZN(n528) );
  NAND2_X1 U577 ( .A1(G113), .A2(n885), .ZN(n530) );
  NAND2_X1 U578 ( .A1(G125), .A2(n886), .ZN(n529) );
  NAND2_X1 U579 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U580 ( .A1(n532), .A2(n531), .ZN(G160) );
  NAND2_X1 U581 ( .A1(G102), .A2(n881), .ZN(n534) );
  NAND2_X1 U582 ( .A1(G138), .A2(n882), .ZN(n533) );
  NAND2_X1 U583 ( .A1(n534), .A2(n533), .ZN(n541) );
  NAND2_X1 U584 ( .A1(n886), .A2(G126), .ZN(n535) );
  XNOR2_X1 U585 ( .A(n535), .B(KEYINPUT88), .ZN(n537) );
  NAND2_X1 U586 ( .A1(G114), .A2(n885), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n537), .A2(n536), .ZN(n539) );
  XNOR2_X1 U588 ( .A(n539), .B(n538), .ZN(n540) );
  NOR2_X1 U589 ( .A1(n541), .A2(n540), .ZN(G164) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n542) );
  XNOR2_X1 U591 ( .A(KEYINPUT66), .B(n542), .ZN(n642) );
  NAND2_X1 U592 ( .A1(n662), .A2(G51), .ZN(n545) );
  XNOR2_X1 U593 ( .A(G651), .B(KEYINPUT67), .ZN(n548) );
  NOR2_X1 U594 ( .A1(G543), .A2(n548), .ZN(n543) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n543), .Z(n663) );
  NAND2_X1 U596 ( .A1(G63), .A2(n663), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U598 ( .A(KEYINPUT6), .B(n546), .ZN(n554) );
  NOR2_X1 U599 ( .A1(G543), .A2(G651), .ZN(n658) );
  NAND2_X1 U600 ( .A1(n658), .A2(G89), .ZN(n547) );
  XNOR2_X1 U601 ( .A(n547), .B(KEYINPUT4), .ZN(n550) );
  NOR2_X1 U602 ( .A1(n642), .A2(n548), .ZN(n659) );
  NAND2_X1 U603 ( .A1(G76), .A2(n659), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U605 ( .A(KEYINPUT5), .B(n551), .ZN(n552) );
  XNOR2_X1 U606 ( .A(KEYINPUT75), .B(n552), .ZN(n553) );
  NOR2_X1 U607 ( .A1(n554), .A2(n553), .ZN(n557) );
  XNOR2_X1 U608 ( .A(KEYINPUT7), .B(KEYINPUT76), .ZN(n555) );
  XNOR2_X1 U609 ( .A(n555), .B(KEYINPUT77), .ZN(n556) );
  XNOR2_X1 U610 ( .A(n557), .B(n556), .ZN(G168) );
  XOR2_X1 U611 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U612 ( .A1(G85), .A2(n658), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G72), .A2(n659), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U615 ( .A1(n662), .A2(G47), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G60), .A2(n663), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n562) );
  OR2_X1 U618 ( .A1(n563), .A2(n562), .ZN(G290) );
  XOR2_X1 U619 ( .A(G2435), .B(G2454), .Z(n565) );
  XNOR2_X1 U620 ( .A(G2430), .B(G2438), .ZN(n564) );
  XNOR2_X1 U621 ( .A(n565), .B(n564), .ZN(n572) );
  XOR2_X1 U622 ( .A(G2446), .B(KEYINPUT105), .Z(n567) );
  XNOR2_X1 U623 ( .A(G2451), .B(G2443), .ZN(n566) );
  XNOR2_X1 U624 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U625 ( .A(n568), .B(G2427), .Z(n570) );
  XNOR2_X1 U626 ( .A(G1348), .B(G1341), .ZN(n569) );
  XNOR2_X1 U627 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U628 ( .A(n572), .B(n571), .ZN(n573) );
  AND2_X1 U629 ( .A1(n573), .A2(G14), .ZN(G401) );
  NAND2_X1 U630 ( .A1(n662), .A2(G52), .ZN(n574) );
  XNOR2_X1 U631 ( .A(n574), .B(KEYINPUT68), .ZN(n576) );
  NAND2_X1 U632 ( .A1(G64), .A2(n663), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n576), .A2(n575), .ZN(n582) );
  NAND2_X1 U634 ( .A1(G90), .A2(n658), .ZN(n578) );
  NAND2_X1 U635 ( .A1(G77), .A2(n659), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U637 ( .A(KEYINPUT9), .B(n579), .ZN(n580) );
  XNOR2_X1 U638 ( .A(KEYINPUT69), .B(n580), .ZN(n581) );
  NOR2_X1 U639 ( .A1(n582), .A2(n581), .ZN(G171) );
  INV_X1 U640 ( .A(G171), .ZN(G301) );
  AND2_X1 U641 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U642 ( .A(G57), .ZN(G237) );
  INV_X1 U643 ( .A(G108), .ZN(G238) );
  INV_X1 U644 ( .A(G132), .ZN(G219) );
  INV_X1 U645 ( .A(G82), .ZN(G220) );
  NAND2_X1 U646 ( .A1(G75), .A2(n659), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT83), .B(n583), .Z(n585) );
  NAND2_X1 U648 ( .A1(n658), .A2(G88), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT84), .B(n586), .Z(n590) );
  NAND2_X1 U651 ( .A1(n663), .A2(G62), .ZN(n588) );
  NAND2_X1 U652 ( .A1(n662), .A2(G50), .ZN(n587) );
  AND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(G303) );
  NAND2_X1 U655 ( .A1(G7), .A2(G661), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n591), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U657 ( .A(G223), .ZN(n832) );
  NAND2_X1 U658 ( .A1(n832), .A2(G567), .ZN(n592) );
  XOR2_X1 U659 ( .A(KEYINPUT11), .B(n592), .Z(G234) );
  XNOR2_X1 U660 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n598) );
  NAND2_X1 U661 ( .A1(n658), .A2(G81), .ZN(n593) );
  XNOR2_X1 U662 ( .A(n593), .B(KEYINPUT12), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G68), .A2(n659), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U665 ( .A(n596), .B(KEYINPUT13), .ZN(n597) );
  XNOR2_X1 U666 ( .A(n598), .B(n597), .ZN(n602) );
  NAND2_X1 U667 ( .A1(n663), .A2(G56), .ZN(n599) );
  XNOR2_X1 U668 ( .A(n599), .B(KEYINPUT71), .ZN(n600) );
  XNOR2_X1 U669 ( .A(n600), .B(KEYINPUT14), .ZN(n601) );
  NOR2_X1 U670 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U671 ( .A1(n662), .A2(G43), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n604), .A2(n603), .ZN(n1003) );
  INV_X1 U673 ( .A(G860), .ZN(n625) );
  OR2_X1 U674 ( .A1(n1003), .A2(n625), .ZN(G153) );
  NAND2_X1 U675 ( .A1(G868), .A2(G301), .ZN(n614) );
  NAND2_X1 U676 ( .A1(G54), .A2(n662), .ZN(n611) );
  NAND2_X1 U677 ( .A1(n658), .A2(G92), .ZN(n606) );
  NAND2_X1 U678 ( .A1(G66), .A2(n663), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n659), .A2(G79), .ZN(n607) );
  XOR2_X1 U681 ( .A(KEYINPUT74), .B(n607), .Z(n608) );
  NOR2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n612), .B(KEYINPUT15), .ZN(n1008) );
  OR2_X1 U685 ( .A1(n1008), .A2(G868), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(G284) );
  NAND2_X1 U687 ( .A1(G91), .A2(n658), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G78), .A2(n659), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U690 ( .A(KEYINPUT70), .B(n617), .Z(n621) );
  NAND2_X1 U691 ( .A1(n663), .A2(G65), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n662), .A2(G53), .ZN(n618) );
  AND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(G299) );
  INV_X1 U695 ( .A(G868), .ZN(n674) );
  NOR2_X1 U696 ( .A1(G286), .A2(n674), .ZN(n623) );
  NOR2_X1 U697 ( .A1(G868), .A2(G299), .ZN(n622) );
  NOR2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U699 ( .A(KEYINPUT78), .B(n624), .ZN(G297) );
  NAND2_X1 U700 ( .A1(n625), .A2(G559), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n626), .A2(n1008), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n627), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U703 ( .A1(G868), .A2(n1003), .ZN(n630) );
  NAND2_X1 U704 ( .A1(G868), .A2(n1008), .ZN(n628) );
  NOR2_X1 U705 ( .A1(G559), .A2(n628), .ZN(n629) );
  NOR2_X1 U706 ( .A1(n630), .A2(n629), .ZN(G282) );
  NAND2_X1 U707 ( .A1(G111), .A2(n885), .ZN(n637) );
  NAND2_X1 U708 ( .A1(G99), .A2(n881), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G135), .A2(n882), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n886), .A2(G123), .ZN(n633) );
  XOR2_X1 U712 ( .A(KEYINPUT18), .B(n633), .Z(n634) );
  NOR2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U715 ( .A(n638), .B(KEYINPUT79), .ZN(n972) );
  XNOR2_X1 U716 ( .A(n972), .B(G2096), .ZN(n639) );
  XNOR2_X1 U717 ( .A(n639), .B(KEYINPUT80), .ZN(n641) );
  INV_X1 U718 ( .A(G2100), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(G156) );
  NAND2_X1 U720 ( .A1(G49), .A2(n662), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G87), .A2(n642), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U723 ( .A1(n663), .A2(n645), .ZN(n647) );
  NAND2_X1 U724 ( .A1(G651), .A2(G74), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U726 ( .A1(n659), .A2(G73), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n648), .B(KEYINPUT2), .ZN(n655) );
  NAND2_X1 U728 ( .A1(G86), .A2(n658), .ZN(n650) );
  NAND2_X1 U729 ( .A1(G48), .A2(n662), .ZN(n649) );
  NAND2_X1 U730 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n663), .A2(G61), .ZN(n651) );
  XOR2_X1 U732 ( .A(KEYINPUT82), .B(n651), .Z(n652) );
  NOR2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n655), .A2(n654), .ZN(G305) );
  NAND2_X1 U735 ( .A1(n1008), .A2(G559), .ZN(n841) );
  INV_X1 U736 ( .A(G299), .ZN(n1014) );
  XOR2_X1 U737 ( .A(n1003), .B(G288), .Z(n656) );
  XNOR2_X1 U738 ( .A(G290), .B(n656), .ZN(n657) );
  XNOR2_X1 U739 ( .A(KEYINPUT19), .B(n657), .ZN(n670) );
  NAND2_X1 U740 ( .A1(G93), .A2(n658), .ZN(n661) );
  NAND2_X1 U741 ( .A1(G80), .A2(n659), .ZN(n660) );
  NAND2_X1 U742 ( .A1(n661), .A2(n660), .ZN(n667) );
  NAND2_X1 U743 ( .A1(n662), .A2(G55), .ZN(n665) );
  NAND2_X1 U744 ( .A1(G67), .A2(n663), .ZN(n664) );
  NAND2_X1 U745 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U746 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U747 ( .A(KEYINPUT81), .B(n668), .ZN(n843) );
  XOR2_X1 U748 ( .A(G305), .B(n843), .Z(n669) );
  XNOR2_X1 U749 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U750 ( .A(n1014), .B(n671), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n672), .B(G303), .ZN(n906) );
  XNOR2_X1 U752 ( .A(n841), .B(n906), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n673), .A2(G868), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n674), .A2(n843), .ZN(n675) );
  NAND2_X1 U755 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U757 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U760 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XOR2_X1 U761 ( .A(KEYINPUT85), .B(G44), .Z(n681) );
  XNOR2_X1 U762 ( .A(KEYINPUT3), .B(n681), .ZN(G218) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U764 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U765 ( .A1(G218), .A2(n683), .ZN(n684) );
  NAND2_X1 U766 ( .A1(G96), .A2(n684), .ZN(n839) );
  NAND2_X1 U767 ( .A1(n839), .A2(G2106), .ZN(n690) );
  NAND2_X1 U768 ( .A1(G120), .A2(G69), .ZN(n685) );
  NOR2_X1 U769 ( .A1(G237), .A2(n685), .ZN(n686) );
  XOR2_X1 U770 ( .A(KEYINPUT86), .B(n686), .Z(n687) );
  NOR2_X1 U771 ( .A1(G238), .A2(n687), .ZN(n688) );
  XNOR2_X1 U772 ( .A(KEYINPUT87), .B(n688), .ZN(n840) );
  NAND2_X1 U773 ( .A1(n840), .A2(G567), .ZN(n689) );
  NAND2_X1 U774 ( .A1(n690), .A2(n689), .ZN(n918) );
  NAND2_X1 U775 ( .A1(G483), .A2(G661), .ZN(n691) );
  NOR2_X1 U776 ( .A1(n918), .A2(n691), .ZN(n838) );
  NAND2_X1 U777 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U778 ( .A1(n886), .A2(G119), .ZN(n692) );
  XOR2_X1 U779 ( .A(KEYINPUT93), .B(n692), .Z(n694) );
  NAND2_X1 U780 ( .A1(n885), .A2(G107), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U782 ( .A(KEYINPUT94), .B(n695), .Z(n699) );
  NAND2_X1 U783 ( .A1(n881), .A2(G95), .ZN(n697) );
  NAND2_X1 U784 ( .A1(G131), .A2(n882), .ZN(n696) );
  AND2_X1 U785 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n902) );
  NAND2_X1 U787 ( .A1(G1991), .A2(n902), .ZN(n700) );
  XNOR2_X1 U788 ( .A(n700), .B(KEYINPUT95), .ZN(n711) );
  NAND2_X1 U789 ( .A1(G105), .A2(n881), .ZN(n701) );
  XNOR2_X1 U790 ( .A(n701), .B(KEYINPUT38), .ZN(n709) );
  NAND2_X1 U791 ( .A1(G129), .A2(n886), .ZN(n702) );
  XNOR2_X1 U792 ( .A(n702), .B(KEYINPUT96), .ZN(n704) );
  NAND2_X1 U793 ( .A1(n885), .A2(G117), .ZN(n703) );
  NAND2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U795 ( .A1(G141), .A2(n882), .ZN(n705) );
  XNOR2_X1 U796 ( .A(KEYINPUT97), .B(n705), .ZN(n706) );
  NOR2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n897) );
  AND2_X1 U799 ( .A1(G1996), .A2(n897), .ZN(n710) );
  NOR2_X1 U800 ( .A1(n711), .A2(n710), .ZN(n982) );
  NAND2_X1 U801 ( .A1(G160), .A2(G40), .ZN(n726) );
  NOR2_X1 U802 ( .A1(n727), .A2(n726), .ZN(n827) );
  INV_X1 U803 ( .A(n827), .ZN(n712) );
  NOR2_X1 U804 ( .A1(n982), .A2(n712), .ZN(n818) );
  INV_X1 U805 ( .A(n818), .ZN(n724) );
  NAND2_X1 U806 ( .A1(G104), .A2(n881), .ZN(n714) );
  NAND2_X1 U807 ( .A1(G140), .A2(n882), .ZN(n713) );
  NAND2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U809 ( .A(KEYINPUT34), .B(n715), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n886), .A2(G128), .ZN(n716) );
  XOR2_X1 U811 ( .A(KEYINPUT91), .B(n716), .Z(n718) );
  NAND2_X1 U812 ( .A1(n885), .A2(G116), .ZN(n717) );
  NAND2_X1 U813 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U814 ( .A(n719), .B(KEYINPUT35), .Z(n720) );
  NOR2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U816 ( .A(KEYINPUT36), .B(n722), .Z(n723) );
  XOR2_X1 U817 ( .A(KEYINPUT92), .B(n723), .Z(n896) );
  XNOR2_X1 U818 ( .A(G2067), .B(KEYINPUT37), .ZN(n823) );
  NOR2_X1 U819 ( .A1(n896), .A2(n823), .ZN(n974) );
  NAND2_X1 U820 ( .A1(n827), .A2(n974), .ZN(n821) );
  NAND2_X1 U821 ( .A1(n724), .A2(n821), .ZN(n725) );
  XNOR2_X1 U822 ( .A(n725), .B(KEYINPUT98), .ZN(n812) );
  INV_X1 U823 ( .A(G286), .ZN(n770) );
  INV_X1 U824 ( .A(n726), .ZN(n728) );
  XOR2_X1 U825 ( .A(n754), .B(KEYINPUT100), .Z(n756) );
  INV_X1 U826 ( .A(n756), .ZN(n735) );
  NAND2_X1 U827 ( .A1(G2072), .A2(n735), .ZN(n729) );
  XNOR2_X1 U828 ( .A(n729), .B(KEYINPUT27), .ZN(n731) );
  INV_X1 U829 ( .A(G1956), .ZN(n922) );
  NOR2_X1 U830 ( .A1(n735), .A2(n922), .ZN(n730) );
  NOR2_X1 U831 ( .A1(n731), .A2(n730), .ZN(n734) );
  NOR2_X1 U832 ( .A1(n1014), .A2(n734), .ZN(n733) );
  XNOR2_X1 U833 ( .A(n733), .B(n732), .ZN(n752) );
  NAND2_X1 U834 ( .A1(n1014), .A2(n734), .ZN(n750) );
  AND2_X1 U835 ( .A1(n735), .A2(G2067), .ZN(n737) );
  INV_X1 U836 ( .A(G1348), .ZN(n920) );
  NOR2_X1 U837 ( .A1(n754), .A2(n920), .ZN(n736) );
  NOR2_X1 U838 ( .A1(n737), .A2(n736), .ZN(n738) );
  OR2_X1 U839 ( .A1(n1008), .A2(n738), .ZN(n748) );
  NAND2_X1 U840 ( .A1(n1008), .A2(n738), .ZN(n746) );
  INV_X1 U841 ( .A(G1996), .ZN(n946) );
  NOR2_X1 U842 ( .A1(n771), .A2(n946), .ZN(n740) );
  XOR2_X1 U843 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n739) );
  XNOR2_X1 U844 ( .A(n740), .B(n739), .ZN(n742) );
  NAND2_X1 U845 ( .A1(n771), .A2(G1341), .ZN(n741) );
  NAND2_X1 U846 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U847 ( .A1(n1003), .A2(n743), .ZN(n744) );
  XNOR2_X1 U848 ( .A(KEYINPUT65), .B(n744), .ZN(n745) );
  NAND2_X1 U849 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U850 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U851 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U852 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U853 ( .A(n753), .B(KEYINPUT29), .ZN(n760) );
  NOR2_X1 U854 ( .A1(n754), .A2(G1961), .ZN(n755) );
  XOR2_X1 U855 ( .A(KEYINPUT99), .B(n755), .Z(n758) );
  XOR2_X1 U856 ( .A(KEYINPUT25), .B(G2078), .Z(n950) );
  NOR2_X1 U857 ( .A1(n950), .A2(n756), .ZN(n757) );
  NOR2_X1 U858 ( .A1(n758), .A2(n757), .ZN(n764) );
  NOR2_X1 U859 ( .A1(G301), .A2(n764), .ZN(n759) );
  NOR2_X1 U860 ( .A1(n760), .A2(n759), .ZN(n769) );
  NAND2_X1 U861 ( .A1(G8), .A2(n771), .ZN(n805) );
  NOR2_X1 U862 ( .A1(G1966), .A2(n805), .ZN(n780) );
  NOR2_X1 U863 ( .A1(G2084), .A2(n771), .ZN(n781) );
  NOR2_X1 U864 ( .A1(n780), .A2(n781), .ZN(n761) );
  NAND2_X1 U865 ( .A1(G8), .A2(n761), .ZN(n762) );
  XNOR2_X1 U866 ( .A(KEYINPUT30), .B(n762), .ZN(n763) );
  NOR2_X1 U867 ( .A1(G168), .A2(n763), .ZN(n766) );
  AND2_X1 U868 ( .A1(G301), .A2(n764), .ZN(n765) );
  NOR2_X1 U869 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U870 ( .A(n767), .B(KEYINPUT31), .ZN(n768) );
  NOR2_X1 U871 ( .A1(n769), .A2(n768), .ZN(n779) );
  NOR2_X1 U872 ( .A1(G1971), .A2(n805), .ZN(n773) );
  NOR2_X1 U873 ( .A1(G2090), .A2(n771), .ZN(n772) );
  NOR2_X1 U874 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U875 ( .A1(n774), .A2(G303), .ZN(n775) );
  NAND2_X1 U876 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U877 ( .A1(G8), .A2(n777), .ZN(n778) );
  XNOR2_X1 U878 ( .A(n778), .B(KEYINPUT32), .ZN(n786) );
  NOR2_X1 U879 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U880 ( .A1(G8), .A2(n781), .ZN(n782) );
  NAND2_X1 U881 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U882 ( .A(KEYINPUT101), .B(n784), .Z(n785) );
  NAND2_X1 U883 ( .A1(n786), .A2(n785), .ZN(n804) );
  NOR2_X1 U884 ( .A1(G1976), .A2(G288), .ZN(n794) );
  NOR2_X1 U885 ( .A1(G1971), .A2(G303), .ZN(n787) );
  NOR2_X1 U886 ( .A1(n794), .A2(n787), .ZN(n1013) );
  NAND2_X1 U887 ( .A1(n804), .A2(n1013), .ZN(n790) );
  NAND2_X1 U888 ( .A1(G1976), .A2(G288), .ZN(n1012) );
  INV_X1 U889 ( .A(KEYINPUT33), .ZN(n791) );
  NAND2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n799) );
  XOR2_X1 U891 ( .A(G1981), .B(KEYINPUT102), .Z(n793) );
  XNOR2_X1 U892 ( .A(G305), .B(n793), .ZN(n1000) );
  INV_X1 U893 ( .A(n1000), .ZN(n797) );
  NAND2_X1 U894 ( .A1(n794), .A2(KEYINPUT33), .ZN(n795) );
  NOR2_X1 U895 ( .A1(n805), .A2(n795), .ZN(n796) );
  NOR2_X1 U896 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U897 ( .A1(n799), .A2(n798), .ZN(n810) );
  NOR2_X1 U898 ( .A1(G1981), .A2(G305), .ZN(n800) );
  XOR2_X1 U899 ( .A(n800), .B(KEYINPUT24), .Z(n801) );
  OR2_X1 U900 ( .A1(n805), .A2(n801), .ZN(n808) );
  NOR2_X1 U901 ( .A1(G2090), .A2(G303), .ZN(n802) );
  NAND2_X1 U902 ( .A1(G8), .A2(n802), .ZN(n803) );
  NAND2_X1 U903 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U904 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n809) );
  AND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n815) );
  XNOR2_X1 U908 ( .A(KEYINPUT90), .B(G1986), .ZN(n813) );
  XNOR2_X1 U909 ( .A(n813), .B(G290), .ZN(n1005) );
  NAND2_X1 U910 ( .A1(n1005), .A2(n827), .ZN(n814) );
  NAND2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n830) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n897), .ZN(n979) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U914 ( .A1(G1991), .A2(n902), .ZN(n973) );
  NOR2_X1 U915 ( .A1(n816), .A2(n973), .ZN(n817) );
  NOR2_X1 U916 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U917 ( .A1(n979), .A2(n819), .ZN(n820) );
  XNOR2_X1 U918 ( .A(n820), .B(KEYINPUT39), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n825) );
  AND2_X1 U920 ( .A1(n896), .A2(n823), .ZN(n824) );
  XNOR2_X1 U921 ( .A(n824), .B(KEYINPUT103), .ZN(n989) );
  NAND2_X1 U922 ( .A1(n825), .A2(n989), .ZN(n826) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U924 ( .A(KEYINPUT104), .B(n828), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U926 ( .A(KEYINPUT40), .B(n831), .ZN(G329) );
  NAND2_X1 U927 ( .A1(n832), .A2(G2106), .ZN(n833) );
  XNOR2_X1 U928 ( .A(n833), .B(KEYINPUT106), .ZN(G217) );
  NAND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n835) );
  INV_X1 U930 ( .A(G661), .ZN(n834) );
  NOR2_X1 U931 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U932 ( .A(n836), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  INV_X1 U938 ( .A(G69), .ZN(G235) );
  NOR2_X1 U939 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U941 ( .A(n1003), .B(n841), .ZN(n842) );
  NOR2_X1 U942 ( .A1(n842), .A2(G860), .ZN(n844) );
  XOR2_X1 U943 ( .A(n844), .B(n843), .Z(G145) );
  XOR2_X1 U944 ( .A(G2100), .B(G2096), .Z(n846) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(G2090), .Z(n848) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U950 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U951 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U953 ( .A(KEYINPUT108), .B(G1991), .Z(n854) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1981), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U956 ( .A(n855), .B(KEYINPUT41), .Z(n857) );
  XNOR2_X1 U957 ( .A(G1971), .B(G1976), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U959 ( .A(G1986), .B(G1956), .Z(n859) );
  XNOR2_X1 U960 ( .A(G1966), .B(G1961), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U962 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U963 ( .A(G2474), .B(KEYINPUT109), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U965 ( .A1(G124), .A2(n886), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n864), .B(KEYINPUT44), .ZN(n865) );
  XNOR2_X1 U967 ( .A(KEYINPUT110), .B(n865), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G136), .A2(n882), .ZN(n866) );
  XOR2_X1 U969 ( .A(KEYINPUT111), .B(n866), .Z(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G100), .A2(n881), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G112), .A2(n885), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U974 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U975 ( .A1(G118), .A2(n885), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G130), .A2(n886), .ZN(n873) );
  NAND2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G106), .A2(n881), .ZN(n876) );
  NAND2_X1 U979 ( .A1(G142), .A2(n882), .ZN(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U981 ( .A(KEYINPUT45), .B(n877), .Z(n878) );
  NOR2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U983 ( .A(n880), .B(KEYINPUT48), .Z(n894) );
  NAND2_X1 U984 ( .A1(G103), .A2(n881), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n892) );
  NAND2_X1 U987 ( .A1(G115), .A2(n885), .ZN(n888) );
  NAND2_X1 U988 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U990 ( .A(KEYINPUT112), .B(n889), .Z(n890) );
  XNOR2_X1 U991 ( .A(KEYINPUT47), .B(n890), .ZN(n891) );
  NOR2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n983) );
  XNOR2_X1 U993 ( .A(n983), .B(KEYINPUT46), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n901) );
  XOR2_X1 U996 ( .A(G162), .B(n972), .Z(n899) );
  XOR2_X1 U997 ( .A(G160), .B(n897), .Z(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n902), .B(G164), .Z(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1003 ( .A(n1008), .B(G286), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n908), .B(G301), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n909), .ZN(G397) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n918), .ZN(n910) );
  XOR2_X1 U1008 ( .A(KEYINPUT113), .B(n910), .Z(n914) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n911) );
  XOR2_X1 U1010 ( .A(KEYINPUT49), .B(n911), .Z(n912) );
  XNOR2_X1 U1011 ( .A(KEYINPUT114), .B(n912), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(KEYINPUT115), .B(n915), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G303), .ZN(G166) );
  INV_X1 U1018 ( .A(n918), .ZN(G319) );
  XNOR2_X1 U1019 ( .A(G21), .B(G1966), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(n919), .B(KEYINPUT125), .ZN(n942) );
  XOR2_X1 U1021 ( .A(G1961), .B(G5), .Z(n932) );
  XNOR2_X1 U1022 ( .A(KEYINPUT59), .B(G4), .ZN(n921) );
  XNOR2_X1 U1023 ( .A(n921), .B(n920), .ZN(n929) );
  XOR2_X1 U1024 ( .A(G1341), .B(G19), .Z(n924) );
  XNOR2_X1 U1025 ( .A(n922), .B(G20), .ZN(n923) );
  NAND2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(G6), .B(G1981), .ZN(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1029 ( .A(KEYINPUT124), .B(n927), .Z(n928) );
  NOR2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(n930), .B(KEYINPUT60), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(G1971), .B(G22), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(G23), .B(G1976), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n937) );
  XOR2_X1 U1036 ( .A(G1986), .B(KEYINPUT126), .Z(n935) );
  XNOR2_X1 U1037 ( .A(G24), .B(n935), .ZN(n936) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(KEYINPUT58), .B(n938), .ZN(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1042 ( .A(n943), .B(KEYINPUT127), .Z(n944) );
  XNOR2_X1 U1043 ( .A(KEYINPUT61), .B(n944), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(G16), .A2(n945), .ZN(n970) );
  XNOR2_X1 U1045 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n994) );
  XNOR2_X1 U1046 ( .A(G32), .B(n946), .ZN(n947) );
  NAND2_X1 U1047 ( .A1(n947), .A2(G28), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(G2072), .B(G33), .ZN(n949) );
  XNOR2_X1 U1049 ( .A(G1991), .B(G25), .ZN(n948) );
  NOR2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(n950), .B(G27), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n951) );
  NOR2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1056 ( .A(KEYINPUT118), .B(n957), .Z(n958) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n958), .ZN(n964) );
  XOR2_X1 U1058 ( .A(G34), .B(KEYINPUT119), .Z(n960) );
  XNOR2_X1 U1059 ( .A(G2084), .B(KEYINPUT54), .ZN(n959) );
  XNOR2_X1 U1060 ( .A(n960), .B(n959), .ZN(n962) );
  XNOR2_X1 U1061 ( .A(G35), .B(G2090), .ZN(n961) );
  NOR2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1064 ( .A(n994), .B(n965), .ZN(n967) );
  INV_X1 U1065 ( .A(G29), .ZN(n966) );
  NAND2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1067 ( .A1(G11), .A2(n968), .ZN(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n998) );
  XOR2_X1 U1069 ( .A(G2084), .B(G160), .Z(n971) );
  NOR2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(KEYINPUT116), .B(n977), .ZN(n992) );
  XOR2_X1 U1074 ( .A(G2090), .B(G162), .Z(n978) );
  NOR2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1076 ( .A(KEYINPUT51), .B(n980), .Z(n981) );
  NAND2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n988) );
  XOR2_X1 U1078 ( .A(G2072), .B(n983), .Z(n985) );
  XOR2_X1 U1079 ( .A(G164), .B(G2078), .Z(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1081 ( .A(KEYINPUT50), .B(n986), .Z(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(KEYINPUT52), .B(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(n996), .A2(G29), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1028) );
  XOR2_X1 U1089 ( .A(G16), .B(KEYINPUT56), .Z(n1026) );
  XNOR2_X1 U1090 ( .A(G1966), .B(KEYINPUT120), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(n999), .B(G168), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1002), .B(KEYINPUT57), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G1341), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1023) );
  XNOR2_X1 U1097 ( .A(n1008), .B(G1348), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G171), .B(G1961), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(n1011), .B(KEYINPUT121), .ZN(n1021) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(n1014), .B(G1956), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(G1971), .A2(G303), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(n1019), .B(KEYINPUT122), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1109 ( .A(KEYINPUT123), .B(n1024), .Z(n1025) );
  NOR2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(n1029), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

