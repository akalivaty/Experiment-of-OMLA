

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U557 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X2 U558 ( .A1(n563), .A2(n562), .ZN(G160) );
  NOR2_X1 U559 ( .A1(G164), .A2(G1384), .ZN(n794) );
  NOR2_X2 U560 ( .A1(n527), .A2(G2105), .ZN(n876) );
  NOR2_X2 U561 ( .A1(n711), .A2(n1020), .ZN(n714) );
  NOR2_X1 U562 ( .A1(n743), .A2(n742), .ZN(n759) );
  INV_X1 U563 ( .A(KEYINPUT67), .ZN(n555) );
  INV_X1 U564 ( .A(KEYINPUT94), .ZN(n712) );
  NOR2_X1 U565 ( .A1(n724), .A2(n1009), .ZN(n725) );
  NOR2_X1 U566 ( .A1(n759), .A2(n758), .ZN(n760) );
  INV_X1 U567 ( .A(KEYINPUT95), .ZN(n762) );
  XNOR2_X1 U568 ( .A(n763), .B(n762), .ZN(n764) );
  INV_X1 U569 ( .A(KEYINPUT97), .ZN(n779) );
  NAND2_X1 U570 ( .A1(G160), .A2(G40), .ZN(n793) );
  XOR2_X1 U571 ( .A(KEYINPUT64), .B(G2104), .Z(n527) );
  NAND2_X1 U572 ( .A1(n833), .A2(n824), .ZN(n825) );
  NOR2_X1 U573 ( .A1(G651), .A2(n645), .ZN(n660) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XOR2_X1 U575 ( .A(KEYINPUT17), .B(n522), .Z(n875) );
  NAND2_X1 U576 ( .A1(G138), .A2(n875), .ZN(n525) );
  NAND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X2 U578 ( .A(KEYINPUT66), .B(n523), .Z(n872) );
  NAND2_X1 U579 ( .A1(G114), .A2(n872), .ZN(n524) );
  NAND2_X1 U580 ( .A1(n525), .A2(n524), .ZN(n531) );
  NAND2_X1 U581 ( .A1(G2105), .A2(n527), .ZN(n526) );
  XNOR2_X2 U582 ( .A(n526), .B(KEYINPUT65), .ZN(n871) );
  NAND2_X1 U583 ( .A1(n871), .A2(G126), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n876), .A2(G102), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U586 ( .A1(n531), .A2(n530), .ZN(G164) );
  XOR2_X1 U587 ( .A(KEYINPUT102), .B(G2443), .Z(n533) );
  XNOR2_X1 U588 ( .A(G2451), .B(G2427), .ZN(n532) );
  XNOR2_X1 U589 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U590 ( .A(n534), .B(G2430), .Z(n536) );
  XNOR2_X1 U591 ( .A(G1341), .B(G1348), .ZN(n535) );
  XNOR2_X1 U592 ( .A(n536), .B(n535), .ZN(n540) );
  XOR2_X1 U593 ( .A(KEYINPUT103), .B(G2435), .Z(n538) );
  XNOR2_X1 U594 ( .A(G2438), .B(G2454), .ZN(n537) );
  XNOR2_X1 U595 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U596 ( .A(n540), .B(n539), .Z(n542) );
  XNOR2_X1 U597 ( .A(G2446), .B(KEYINPUT101), .ZN(n541) );
  XNOR2_X1 U598 ( .A(n542), .B(n541), .ZN(n543) );
  AND2_X1 U599 ( .A1(n543), .A2(G14), .ZN(G401) );
  INV_X1 U600 ( .A(G651), .ZN(n546) );
  NOR2_X1 U601 ( .A1(G543), .A2(n546), .ZN(n544) );
  XOR2_X1 U602 ( .A(KEYINPUT1), .B(n544), .Z(n659) );
  NAND2_X1 U603 ( .A1(G64), .A2(n659), .ZN(n545) );
  XNOR2_X1 U604 ( .A(n545), .B(KEYINPUT69), .ZN(n554) );
  NOR2_X1 U605 ( .A1(G651), .A2(G543), .ZN(n657) );
  NAND2_X1 U606 ( .A1(G90), .A2(n657), .ZN(n549) );
  XOR2_X1 U607 ( .A(KEYINPUT0), .B(G543), .Z(n645) );
  OR2_X1 U608 ( .A1(n546), .A2(n645), .ZN(n547) );
  XOR2_X1 U609 ( .A(KEYINPUT68), .B(n547), .Z(n663) );
  NAND2_X1 U610 ( .A1(G77), .A2(n663), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U612 ( .A(n550), .B(KEYINPUT9), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G52), .A2(n660), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U615 ( .A1(n554), .A2(n553), .ZN(G171) );
  AND2_X1 U616 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U617 ( .A(G120), .ZN(G236) );
  INV_X1 U618 ( .A(G69), .ZN(G235) );
  INV_X1 U619 ( .A(G57), .ZN(G237) );
  INV_X1 U620 ( .A(G132), .ZN(G219) );
  INV_X1 U621 ( .A(G82), .ZN(G220) );
  NAND2_X1 U622 ( .A1(n872), .A2(G113), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n559) );
  NAND2_X1 U624 ( .A1(G101), .A2(n876), .ZN(n557) );
  XOR2_X1 U625 ( .A(KEYINPUT23), .B(n557), .Z(n558) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G137), .A2(n875), .ZN(n561) );
  NAND2_X1 U628 ( .A1(G125), .A2(n871), .ZN(n560) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U630 ( .A1(G63), .A2(n659), .ZN(n565) );
  NAND2_X1 U631 ( .A1(G51), .A2(n660), .ZN(n564) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(KEYINPUT6), .B(n566), .ZN(n573) );
  NAND2_X1 U634 ( .A1(G89), .A2(n657), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT4), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(KEYINPUT74), .ZN(n570) );
  NAND2_X1 U637 ( .A1(G76), .A2(n663), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U639 ( .A(n571), .B(KEYINPUT5), .Z(n572) );
  NOR2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U641 ( .A(KEYINPUT7), .B(n574), .Z(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT75), .B(n575), .Z(G168) );
  XOR2_X1 U643 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U644 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U645 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U646 ( .A(G567), .ZN(n692) );
  NOR2_X1 U647 ( .A1(n692), .A2(G223), .ZN(n577) );
  XNOR2_X1 U648 ( .A(n577), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U649 ( .A1(n657), .A2(G81), .ZN(n578) );
  XNOR2_X1 U650 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U651 ( .A1(G68), .A2(n663), .ZN(n579) );
  NAND2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U653 ( .A(KEYINPUT13), .B(n581), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n659), .A2(G56), .ZN(n582) );
  XNOR2_X1 U655 ( .A(KEYINPUT14), .B(n582), .ZN(n583) );
  NAND2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U657 ( .A(KEYINPUT71), .B(n585), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n660), .A2(G43), .ZN(n586) );
  XNOR2_X1 U659 ( .A(KEYINPUT72), .B(n586), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n1020) );
  INV_X1 U661 ( .A(n1020), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n589), .A2(G860), .ZN(G153) );
  NAND2_X1 U663 ( .A1(G868), .A2(G171), .ZN(n598) );
  NAND2_X1 U664 ( .A1(G92), .A2(n657), .ZN(n591) );
  NAND2_X1 U665 ( .A1(G79), .A2(n663), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U667 ( .A1(G66), .A2(n659), .ZN(n593) );
  NAND2_X1 U668 ( .A1(G54), .A2(n660), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U671 ( .A(KEYINPUT15), .B(n596), .Z(n1006) );
  INV_X1 U672 ( .A(G868), .ZN(n678) );
  NAND2_X1 U673 ( .A1(n1006), .A2(n678), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U675 ( .A(n599), .B(KEYINPUT73), .ZN(G284) );
  NAND2_X1 U676 ( .A1(G91), .A2(n657), .ZN(n601) );
  NAND2_X1 U677 ( .A1(G78), .A2(n663), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U679 ( .A(KEYINPUT70), .B(n602), .Z(n606) );
  NAND2_X1 U680 ( .A1(G65), .A2(n659), .ZN(n604) );
  NAND2_X1 U681 ( .A1(G53), .A2(n660), .ZN(n603) );
  AND2_X1 U682 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U683 ( .A1(n606), .A2(n605), .ZN(G299) );
  NOR2_X1 U684 ( .A1(G868), .A2(G299), .ZN(n607) );
  XNOR2_X1 U685 ( .A(n607), .B(KEYINPUT76), .ZN(n609) );
  NOR2_X1 U686 ( .A1(n678), .A2(G286), .ZN(n608) );
  NOR2_X1 U687 ( .A1(n609), .A2(n608), .ZN(G297) );
  INV_X1 U688 ( .A(G559), .ZN(n610) );
  NOR2_X1 U689 ( .A1(G860), .A2(n610), .ZN(n611) );
  XNOR2_X1 U690 ( .A(KEYINPUT77), .B(n611), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n612), .A2(n1006), .ZN(n613) );
  XNOR2_X1 U692 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U693 ( .A1(G868), .A2(n1020), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G868), .A2(n1006), .ZN(n614) );
  NOR2_X1 U695 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U696 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U697 ( .A1(G135), .A2(n875), .ZN(n618) );
  NAND2_X1 U698 ( .A1(G111), .A2(n872), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G123), .A2(n871), .ZN(n619) );
  XNOR2_X1 U701 ( .A(n619), .B(KEYINPUT18), .ZN(n622) );
  NAND2_X1 U702 ( .A1(G99), .A2(n876), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n620), .B(KEYINPUT78), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n929) );
  XNOR2_X1 U706 ( .A(G2096), .B(n929), .ZN(n626) );
  INV_X1 U707 ( .A(G2100), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(G156) );
  NAND2_X1 U709 ( .A1(n1006), .A2(G559), .ZN(n676) );
  XNOR2_X1 U710 ( .A(n1020), .B(n676), .ZN(n627) );
  NOR2_X1 U711 ( .A1(n627), .A2(G860), .ZN(n635) );
  NAND2_X1 U712 ( .A1(G67), .A2(n659), .ZN(n629) );
  NAND2_X1 U713 ( .A1(G55), .A2(n660), .ZN(n628) );
  NAND2_X1 U714 ( .A1(n629), .A2(n628), .ZN(n634) );
  NAND2_X1 U715 ( .A1(G93), .A2(n657), .ZN(n631) );
  NAND2_X1 U716 ( .A1(G80), .A2(n663), .ZN(n630) );
  NAND2_X1 U717 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U718 ( .A(KEYINPUT79), .B(n632), .Z(n633) );
  OR2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n679) );
  XOR2_X1 U720 ( .A(n635), .B(n679), .Z(G145) );
  NAND2_X1 U721 ( .A1(n663), .A2(G73), .ZN(n636) );
  XNOR2_X1 U722 ( .A(n636), .B(KEYINPUT2), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G86), .A2(n657), .ZN(n638) );
  NAND2_X1 U724 ( .A1(G48), .A2(n660), .ZN(n637) );
  NAND2_X1 U725 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U726 ( .A1(G61), .A2(n659), .ZN(n639) );
  XNOR2_X1 U727 ( .A(KEYINPUT81), .B(n639), .ZN(n640) );
  NOR2_X1 U728 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U730 ( .A1(G49), .A2(n660), .ZN(n644) );
  XNOR2_X1 U731 ( .A(n644), .B(KEYINPUT80), .ZN(n650) );
  NAND2_X1 U732 ( .A1(G87), .A2(n645), .ZN(n647) );
  NAND2_X1 U733 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U734 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U735 ( .A1(n659), .A2(n648), .ZN(n649) );
  NAND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(G288) );
  AND2_X1 U737 ( .A1(G72), .A2(n663), .ZN(n654) );
  NAND2_X1 U738 ( .A1(G85), .A2(n657), .ZN(n652) );
  NAND2_X1 U739 ( .A1(G47), .A2(n660), .ZN(n651) );
  NAND2_X1 U740 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U741 ( .A1(n654), .A2(n653), .ZN(n656) );
  NAND2_X1 U742 ( .A1(n659), .A2(G60), .ZN(n655) );
  NAND2_X1 U743 ( .A1(n656), .A2(n655), .ZN(G290) );
  NAND2_X1 U744 ( .A1(G88), .A2(n657), .ZN(n658) );
  XNOR2_X1 U745 ( .A(n658), .B(KEYINPUT82), .ZN(n668) );
  NAND2_X1 U746 ( .A1(G62), .A2(n659), .ZN(n662) );
  NAND2_X1 U747 ( .A1(G50), .A2(n660), .ZN(n661) );
  NAND2_X1 U748 ( .A1(n662), .A2(n661), .ZN(n666) );
  NAND2_X1 U749 ( .A1(G75), .A2(n663), .ZN(n664) );
  XNOR2_X1 U750 ( .A(KEYINPUT83), .B(n664), .ZN(n665) );
  NOR2_X1 U751 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U752 ( .A1(n668), .A2(n667), .ZN(G303) );
  INV_X1 U753 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U754 ( .A(KEYINPUT84), .B(G305), .ZN(n669) );
  XNOR2_X1 U755 ( .A(n669), .B(G288), .ZN(n670) );
  XNOR2_X1 U756 ( .A(KEYINPUT19), .B(n670), .ZN(n672) );
  XNOR2_X1 U757 ( .A(G290), .B(G166), .ZN(n671) );
  XNOR2_X1 U758 ( .A(n672), .B(n671), .ZN(n673) );
  XOR2_X1 U759 ( .A(n679), .B(n673), .Z(n675) );
  INV_X1 U760 ( .A(G299), .ZN(n1009) );
  XNOR2_X1 U761 ( .A(n1020), .B(n1009), .ZN(n674) );
  XNOR2_X1 U762 ( .A(n675), .B(n674), .ZN(n893) );
  XNOR2_X1 U763 ( .A(n893), .B(n676), .ZN(n677) );
  NOR2_X1 U764 ( .A1(n678), .A2(n677), .ZN(n681) );
  NOR2_X1 U765 ( .A1(G868), .A2(n679), .ZN(n680) );
  NOR2_X1 U766 ( .A1(n681), .A2(n680), .ZN(G295) );
  NAND2_X1 U767 ( .A1(G2078), .A2(G2084), .ZN(n682) );
  XOR2_X1 U768 ( .A(KEYINPUT20), .B(n682), .Z(n683) );
  NAND2_X1 U769 ( .A1(G2090), .A2(n683), .ZN(n684) );
  XNOR2_X1 U770 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U772 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U773 ( .A1(G220), .A2(G219), .ZN(n686) );
  XOR2_X1 U774 ( .A(KEYINPUT22), .B(n686), .Z(n687) );
  NOR2_X1 U775 ( .A1(G218), .A2(n687), .ZN(n688) );
  NAND2_X1 U776 ( .A1(G96), .A2(n688), .ZN(n848) );
  NAND2_X1 U777 ( .A1(G2106), .A2(n848), .ZN(n689) );
  XNOR2_X1 U778 ( .A(n689), .B(KEYINPUT85), .ZN(n694) );
  NOR2_X1 U779 ( .A1(G235), .A2(G236), .ZN(n690) );
  NAND2_X1 U780 ( .A1(G108), .A2(n690), .ZN(n691) );
  NOR2_X1 U781 ( .A1(G237), .A2(n691), .ZN(n847) );
  NOR2_X1 U782 ( .A1(n692), .A2(n847), .ZN(n693) );
  NOR2_X1 U783 ( .A1(n694), .A2(n693), .ZN(G319) );
  INV_X1 U784 ( .A(G319), .ZN(n917) );
  NAND2_X1 U785 ( .A1(G661), .A2(G483), .ZN(n695) );
  XNOR2_X1 U786 ( .A(KEYINPUT86), .B(n695), .ZN(n696) );
  NOR2_X1 U787 ( .A1(n917), .A2(n696), .ZN(n846) );
  NAND2_X1 U788 ( .A1(n846), .A2(G36), .ZN(G176) );
  INV_X1 U789 ( .A(G171), .ZN(G301) );
  INV_X1 U790 ( .A(n794), .ZN(n698) );
  NOR2_X4 U791 ( .A1(n793), .A2(n698), .ZN(n730) );
  INV_X1 U792 ( .A(KEYINPUT92), .ZN(n699) );
  XNOR2_X1 U793 ( .A(n730), .B(n699), .ZN(n729) );
  INV_X1 U794 ( .A(n729), .ZN(n715) );
  NAND2_X1 U795 ( .A1(G2072), .A2(n715), .ZN(n700) );
  XNOR2_X1 U796 ( .A(n700), .B(KEYINPUT27), .ZN(n702) );
  AND2_X1 U797 ( .A1(n729), .A2(G1956), .ZN(n701) );
  NOR2_X1 U798 ( .A1(n702), .A2(n701), .ZN(n724) );
  NAND2_X1 U799 ( .A1(n1009), .A2(n724), .ZN(n723) );
  NAND2_X1 U800 ( .A1(G1996), .A2(n730), .ZN(n703) );
  XNOR2_X1 U801 ( .A(n703), .B(KEYINPUT26), .ZN(n705) );
  INV_X1 U802 ( .A(G1341), .ZN(n951) );
  NOR2_X1 U803 ( .A1(n730), .A2(n951), .ZN(n704) );
  NAND2_X1 U804 ( .A1(KEYINPUT26), .A2(n704), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n705), .A2(n708), .ZN(n707) );
  INV_X1 U806 ( .A(KEYINPUT93), .ZN(n706) );
  NAND2_X1 U807 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U808 ( .A1(n708), .A2(KEYINPUT93), .ZN(n709) );
  NAND2_X1 U809 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U810 ( .A1(n1006), .A2(n714), .ZN(n713) );
  XNOR2_X1 U811 ( .A(n713), .B(n712), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n1006), .A2(n714), .ZN(n719) );
  NAND2_X1 U813 ( .A1(G2067), .A2(n715), .ZN(n717) );
  INV_X1 U814 ( .A(n730), .ZN(n746) );
  NAND2_X1 U815 ( .A1(G1348), .A2(n746), .ZN(n716) );
  NAND2_X1 U816 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U817 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U818 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U819 ( .A1(n723), .A2(n722), .ZN(n727) );
  XOR2_X1 U820 ( .A(n725), .B(KEYINPUT28), .Z(n726) );
  NAND2_X1 U821 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U822 ( .A(n728), .B(KEYINPUT29), .ZN(n734) );
  XOR2_X1 U823 ( .A(G2078), .B(KEYINPUT25), .Z(n984) );
  NOR2_X1 U824 ( .A1(n984), .A2(n729), .ZN(n732) );
  NOR2_X1 U825 ( .A1(n730), .A2(G1961), .ZN(n731) );
  NOR2_X1 U826 ( .A1(n732), .A2(n731), .ZN(n738) );
  NOR2_X1 U827 ( .A1(G301), .A2(n738), .ZN(n733) );
  NOR2_X1 U828 ( .A1(n734), .A2(n733), .ZN(n743) );
  NAND2_X1 U829 ( .A1(G8), .A2(n746), .ZN(n790) );
  NOR2_X1 U830 ( .A1(G1966), .A2(n790), .ZN(n758) );
  NOR2_X1 U831 ( .A1(G2084), .A2(n746), .ZN(n756) );
  NOR2_X1 U832 ( .A1(n758), .A2(n756), .ZN(n735) );
  NAND2_X1 U833 ( .A1(G8), .A2(n735), .ZN(n736) );
  XNOR2_X1 U834 ( .A(KEYINPUT30), .B(n736), .ZN(n737) );
  NOR2_X1 U835 ( .A1(G168), .A2(n737), .ZN(n740) );
  AND2_X1 U836 ( .A1(G301), .A2(n738), .ZN(n739) );
  NOR2_X1 U837 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U838 ( .A(n741), .B(KEYINPUT31), .ZN(n742) );
  INV_X1 U839 ( .A(n759), .ZN(n745) );
  AND2_X1 U840 ( .A1(G286), .A2(G8), .ZN(n744) );
  NAND2_X1 U841 ( .A1(n745), .A2(n744), .ZN(n754) );
  INV_X1 U842 ( .A(G8), .ZN(n752) );
  NOR2_X1 U843 ( .A1(G1971), .A2(n790), .ZN(n748) );
  NOR2_X1 U844 ( .A1(G2090), .A2(n746), .ZN(n747) );
  NOR2_X1 U845 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U846 ( .A1(n749), .A2(G303), .ZN(n750) );
  XNOR2_X1 U847 ( .A(n750), .B(KEYINPUT96), .ZN(n751) );
  OR2_X1 U848 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U849 ( .A(KEYINPUT32), .B(n755), .ZN(n765) );
  NAND2_X1 U850 ( .A1(G8), .A2(n756), .ZN(n757) );
  XOR2_X1 U851 ( .A(KEYINPUT91), .B(n757), .Z(n761) );
  NAND2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n783) );
  NOR2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n1011) );
  NOR2_X1 U855 ( .A1(G1971), .A2(G303), .ZN(n766) );
  NOR2_X1 U856 ( .A1(n1011), .A2(n766), .ZN(n768) );
  INV_X1 U857 ( .A(KEYINPUT33), .ZN(n767) );
  AND2_X1 U858 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n783), .A2(n769), .ZN(n773) );
  INV_X1 U860 ( .A(n790), .ZN(n770) );
  NAND2_X1 U861 ( .A1(G1976), .A2(G288), .ZN(n1012) );
  AND2_X1 U862 ( .A1(n770), .A2(n1012), .ZN(n771) );
  OR2_X1 U863 ( .A1(KEYINPUT33), .A2(n771), .ZN(n772) );
  AND2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n1011), .A2(KEYINPUT33), .ZN(n774) );
  NOR2_X1 U866 ( .A1(n774), .A2(n790), .ZN(n776) );
  XOR2_X1 U867 ( .A(G1981), .B(G305), .Z(n1003) );
  INV_X1 U868 ( .A(n1003), .ZN(n775) );
  NOR2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n780) );
  XNOR2_X1 U871 ( .A(n780), .B(n779), .ZN(n787) );
  NOR2_X1 U872 ( .A1(G2090), .A2(G303), .ZN(n781) );
  NAND2_X1 U873 ( .A1(G8), .A2(n781), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n784), .A2(n790), .ZN(n785) );
  XNOR2_X1 U876 ( .A(n785), .B(KEYINPUT98), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n792) );
  NOR2_X1 U878 ( .A1(G1981), .A2(G305), .ZN(n788) );
  XOR2_X1 U879 ( .A(n788), .B(KEYINPUT24), .Z(n789) );
  NOR2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n826) );
  NOR2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n838) );
  NAND2_X1 U883 ( .A1(G140), .A2(n875), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G104), .A2(n876), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U886 ( .A(KEYINPUT34), .B(n797), .ZN(n803) );
  NAND2_X1 U887 ( .A1(n871), .A2(G128), .ZN(n799) );
  NAND2_X1 U888 ( .A1(G116), .A2(n872), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U890 ( .A(KEYINPUT87), .B(n800), .ZN(n801) );
  XNOR2_X1 U891 ( .A(KEYINPUT35), .B(n801), .ZN(n802) );
  NOR2_X1 U892 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U893 ( .A(n804), .B(KEYINPUT36), .ZN(n805) );
  XNOR2_X1 U894 ( .A(n805), .B(KEYINPUT88), .ZN(n886) );
  XNOR2_X1 U895 ( .A(KEYINPUT37), .B(G2067), .ZN(n835) );
  NOR2_X1 U896 ( .A1(n886), .A2(n835), .ZN(n944) );
  NAND2_X1 U897 ( .A1(n838), .A2(n944), .ZN(n833) );
  NAND2_X1 U898 ( .A1(G107), .A2(n872), .ZN(n808) );
  NAND2_X1 U899 ( .A1(G131), .A2(n875), .ZN(n806) );
  XOR2_X1 U900 ( .A(KEYINPUT89), .B(n806), .Z(n807) );
  NAND2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U902 ( .A1(G95), .A2(n876), .ZN(n810) );
  NAND2_X1 U903 ( .A1(G119), .A2(n871), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n861) );
  INV_X1 U906 ( .A(G1991), .ZN(n980) );
  NOR2_X1 U907 ( .A1(n861), .A2(n980), .ZN(n822) );
  NAND2_X1 U908 ( .A1(G141), .A2(n875), .ZN(n814) );
  NAND2_X1 U909 ( .A1(G117), .A2(n872), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n876), .A2(G105), .ZN(n815) );
  XOR2_X1 U912 ( .A(KEYINPUT38), .B(n815), .Z(n816) );
  NOR2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n871), .A2(G129), .ZN(n818) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n862) );
  NAND2_X1 U916 ( .A1(G1996), .A2(n862), .ZN(n820) );
  XOR2_X1 U917 ( .A(KEYINPUT90), .B(n820), .Z(n821) );
  NOR2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n931) );
  XOR2_X1 U919 ( .A(G1986), .B(G290), .Z(n1007) );
  NAND2_X1 U920 ( .A1(n931), .A2(n1007), .ZN(n823) );
  NAND2_X1 U921 ( .A1(n823), .A2(n838), .ZN(n824) );
  OR2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n841) );
  NOR2_X1 U923 ( .A1(G1996), .A2(n862), .ZN(n924) );
  AND2_X1 U924 ( .A1(n980), .A2(n861), .ZN(n933) );
  NOR2_X1 U925 ( .A1(G1986), .A2(G290), .ZN(n827) );
  XOR2_X1 U926 ( .A(n827), .B(KEYINPUT99), .Z(n828) );
  NOR2_X1 U927 ( .A1(n933), .A2(n828), .ZN(n830) );
  INV_X1 U928 ( .A(n931), .ZN(n829) );
  NOR2_X1 U929 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U930 ( .A1(n924), .A2(n831), .ZN(n832) );
  XNOR2_X1 U931 ( .A(KEYINPUT39), .B(n832), .ZN(n834) );
  NAND2_X1 U932 ( .A1(n834), .A2(n833), .ZN(n836) );
  NAND2_X1 U933 ( .A1(n886), .A2(n835), .ZN(n943) );
  NAND2_X1 U934 ( .A1(n836), .A2(n943), .ZN(n837) );
  XNOR2_X1 U935 ( .A(KEYINPUT100), .B(n837), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n839), .A2(n838), .ZN(n840) );
  NAND2_X1 U937 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U938 ( .A(n842), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U939 ( .A(G223), .ZN(n843) );
  NAND2_X1 U940 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U942 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U944 ( .A1(n846), .A2(n845), .ZN(G188) );
  XOR2_X1 U945 ( .A(G108), .B(KEYINPUT112), .Z(G238) );
  INV_X1 U947 ( .A(n847), .ZN(n849) );
  NOR2_X1 U948 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U949 ( .A(KEYINPUT104), .B(n850), .ZN(G325) );
  XNOR2_X1 U950 ( .A(KEYINPUT105), .B(G325), .ZN(G261) );
  INV_X1 U951 ( .A(G96), .ZN(G221) );
  NAND2_X1 U952 ( .A1(n876), .A2(G100), .ZN(n852) );
  NAND2_X1 U953 ( .A1(G112), .A2(n872), .ZN(n851) );
  NAND2_X1 U954 ( .A1(n852), .A2(n851), .ZN(n857) );
  NAND2_X1 U955 ( .A1(G124), .A2(n871), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n875), .A2(G136), .ZN(n854) );
  NAND2_X1 U958 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U959 ( .A1(n857), .A2(n856), .ZN(G162) );
  XOR2_X1 U960 ( .A(KEYINPUT48), .B(KEYINPUT108), .Z(n859) );
  XNOR2_X1 U961 ( .A(G164), .B(KEYINPUT46), .ZN(n858) );
  XNOR2_X1 U962 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n890) );
  NAND2_X1 U965 ( .A1(G139), .A2(n875), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G103), .A2(n876), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n871), .A2(G127), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G115), .A2(n872), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n868), .Z(n869) );
  NOR2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n936) );
  XNOR2_X1 U973 ( .A(G160), .B(n936), .ZN(n884) );
  NAND2_X1 U974 ( .A1(n871), .A2(G130), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G118), .A2(n872), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G142), .A2(n875), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G106), .A2(n876), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U980 ( .A(KEYINPUT107), .B(n879), .ZN(n880) );
  XNOR2_X1 U981 ( .A(KEYINPUT45), .B(n880), .ZN(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U984 ( .A(n885), .B(n929), .Z(n888) );
  XNOR2_X1 U985 ( .A(n886), .B(G162), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U987 ( .A(n890), .B(n889), .Z(n891) );
  NOR2_X1 U988 ( .A1(G37), .A2(n891), .ZN(n892) );
  XOR2_X1 U989 ( .A(KEYINPUT109), .B(n892), .Z(G395) );
  XOR2_X1 U990 ( .A(n893), .B(G286), .Z(n895) );
  XNOR2_X1 U991 ( .A(G171), .B(n1006), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U993 ( .A1(G37), .A2(n896), .ZN(G397) );
  XOR2_X1 U994 ( .A(G2096), .B(KEYINPUT43), .Z(n898) );
  XNOR2_X1 U995 ( .A(G2090), .B(KEYINPUT42), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U997 ( .A(n899), .B(G2678), .Z(n901) );
  XNOR2_X1 U998 ( .A(G2067), .B(G2072), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U1000 ( .A(KEYINPUT106), .B(G2100), .Z(n903) );
  XNOR2_X1 U1001 ( .A(G2078), .B(G2084), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(G227) );
  XOR2_X1 U1004 ( .A(G1976), .B(G1971), .Z(n907) );
  XNOR2_X1 U1005 ( .A(G1986), .B(G1966), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1007 ( .A(n908), .B(G2474), .Z(n910) );
  XNOR2_X1 U1008 ( .A(G1996), .B(G1991), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n910), .B(n909), .ZN(n914) );
  XOR2_X1 U1010 ( .A(KEYINPUT41), .B(G1956), .Z(n912) );
  XNOR2_X1 U1011 ( .A(G1981), .B(G1961), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(G229) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(G397), .A2(n916), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G401), .A2(n917), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT110), .ZN(n919) );
  NAND2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(G395), .A2(n921), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(KEYINPUT111), .B(n922), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1025 ( .A(KEYINPUT51), .B(n925), .Z(n926) );
  XNOR2_X1 U1026 ( .A(KEYINPUT114), .B(n926), .ZN(n935) );
  XNOR2_X1 U1027 ( .A(G2084), .B(G160), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(KEYINPUT113), .B(n927), .ZN(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(G2072), .B(n936), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(G164), .B(G2078), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1036 ( .A(KEYINPUT115), .B(n939), .Z(n940) );
  XNOR2_X1 U1037 ( .A(KEYINPUT50), .B(n940), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n947) );
  INV_X1 U1039 ( .A(n943), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(KEYINPUT116), .B(n948), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(n949), .B(KEYINPUT52), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n950), .A2(G29), .ZN(n1002) );
  XOR2_X1 U1045 ( .A(G1961), .B(G5), .Z(n961) );
  XNOR2_X1 U1046 ( .A(G19), .B(n951), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(G1981), .B(G6), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(G1956), .B(G20), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1051 ( .A(KEYINPUT59), .B(G1348), .Z(n956) );
  XNOR2_X1 U1052 ( .A(G4), .B(n956), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(KEYINPUT60), .B(n959), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n972) );
  XOR2_X1 U1056 ( .A(G1966), .B(G21), .Z(n970) );
  XOR2_X1 U1057 ( .A(G1986), .B(G24), .Z(n964) );
  XOR2_X1 U1058 ( .A(G22), .B(KEYINPUT126), .Z(n962) );
  XNOR2_X1 U1059 ( .A(n962), .B(G1971), .ZN(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n967) );
  XOR2_X1 U1061 ( .A(KEYINPUT127), .B(G1976), .Z(n965) );
  XNOR2_X1 U1062 ( .A(G23), .B(n965), .ZN(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(n968), .B(KEYINPUT58), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n973), .B(KEYINPUT61), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G16), .B(KEYINPUT125), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(G11), .A2(n976), .ZN(n1000) );
  XOR2_X1 U1071 ( .A(G34), .B(KEYINPUT119), .Z(n978) );
  XNOR2_X1 U1072 ( .A(G2084), .B(KEYINPUT54), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(n978), .B(n977), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(KEYINPUT118), .B(n979), .ZN(n996) );
  XNOR2_X1 U1075 ( .A(G2090), .B(G35), .ZN(n993) );
  XNOR2_X1 U1076 ( .A(G25), .B(n980), .ZN(n981) );
  NAND2_X1 U1077 ( .A1(n981), .A2(G28), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(G2067), .B(G26), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(G33), .B(G2072), .ZN(n982) );
  NOR2_X1 U1080 ( .A1(n983), .A2(n982), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(G1996), .B(G32), .ZN(n986) );
  XNOR2_X1 U1082 ( .A(G27), .B(n984), .ZN(n985) );
  NOR2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1086 ( .A(KEYINPUT53), .B(n991), .ZN(n992) );
  NOR2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1088 ( .A(KEYINPUT117), .B(n994), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(G29), .A2(n997), .ZN(n998) );
  XOR2_X1 U1091 ( .A(KEYINPUT55), .B(n998), .Z(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1033) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G168), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1096 ( .A(KEYINPUT57), .B(n1005), .Z(n1029) );
  XNOR2_X1 U1097 ( .A(n1006), .B(G1348), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1026) );
  XNOR2_X1 U1099 ( .A(G1956), .B(n1009), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(KEYINPUT120), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(KEYINPUT121), .B(n1011), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(G1971), .B(G166), .Z(n1014) );
  XNOR2_X1 U1104 ( .A(KEYINPUT122), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(KEYINPUT123), .B(n1019), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(G301), .B(G1961), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(n1020), .B(G1341), .ZN(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1113 ( .A(KEYINPUT124), .B(n1027), .Z(n1028) );
  NOR2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(G16), .B(KEYINPUT56), .Z(n1030) );
  NOR2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1118 ( .A(n1034), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

