//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n555, new_n556, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(new_n454), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT68), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT69), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT69), .B1(new_n463), .B2(new_n465), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  XOR2_X1   g045(.A(new_n470), .B(KEYINPUT70), .Z(new_n471));
  AOI21_X1  g046(.A(new_n461), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n462), .A2(G2105), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT72), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NOR3_X1   g050(.A1(new_n464), .A2(KEYINPUT71), .A3(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT71), .B1(new_n464), .B2(G2104), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n478), .A2(G137), .A3(new_n461), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n472), .A2(new_n481), .ZN(G160));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(new_n462), .A3(KEYINPUT3), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n479), .A2(new_n484), .A3(new_n465), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT73), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n485), .B(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n487), .A2(new_n461), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(G136), .B2(new_n493), .ZN(G162));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n495), .A2(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n461), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  OAI22_X1  g075(.A1(new_n498), .A2(new_n499), .B1(new_n485), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n478), .A2(KEYINPUT75), .A3(new_n479), .A4(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n479), .A2(new_n484), .A3(new_n465), .A4(new_n503), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT75), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n504), .A2(KEYINPUT4), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n509), .B(new_n503), .C1(new_n467), .C2(new_n468), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n501), .B1(new_n508), .B2(new_n510), .ZN(G164));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT76), .B1(new_n512), .B2(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT76), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(G543), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n517), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G88), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n515), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n521), .A2(new_n527), .A3(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND3_X1  g106(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n526), .A2(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n520), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(new_n526), .A2(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n520), .A2(G52), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n515), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  NAND2_X1  g121(.A1(new_n526), .A2(G81), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n520), .A2(G43), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n515), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n519), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n525), .A2(KEYINPUT78), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n517), .A2(new_n563), .A3(new_n518), .A4(new_n524), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(G91), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n524), .A2(G65), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT79), .Z(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n561), .A2(new_n565), .A3(new_n569), .ZN(G299));
  OR2_X1    g145(.A1(new_n524), .A2(G74), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n520), .A2(G49), .B1(G651), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n562), .A2(G87), .A3(new_n564), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(new_n524), .A2(G61), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n519), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n562), .A2(G86), .A3(new_n564), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT80), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n562), .A2(new_n583), .A3(G86), .A4(new_n564), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n580), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(new_n526), .A2(G85), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n520), .A2(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n587), .B(new_n588), .C1(new_n515), .C2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n562), .A2(G92), .A3(new_n564), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G54), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n524), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n595), .A2(new_n519), .B1(new_n596), .B2(new_n515), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n592), .A2(new_n593), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n594), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n591), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n591), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G299), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  NOR2_X1   g185(.A1(new_n552), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n602), .A2(new_n609), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT82), .Z(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g190(.A(new_n474), .B1(new_n467), .B2(new_n468), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n493), .A2(G135), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n488), .A2(G123), .ZN(new_n621));
  OR2_X1    g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n622), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(G2096), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n619), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT83), .ZN(G156));
  XOR2_X1   g203(.A(G2451), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT84), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n636), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n633), .B(new_n639), .Z(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(G14), .A3(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(G401));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT86), .Z(new_n647));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT17), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n647), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT87), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n650), .A2(new_n646), .A3(new_n648), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n650), .B1(new_n647), .B2(new_n649), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n647), .B2(new_n648), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n653), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2096), .B(G2100), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT88), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n669), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n670), .A2(KEYINPUT20), .A3(new_n669), .ZN(new_n675));
  OAI221_X1 g250(.A(new_n671), .B1(new_n669), .B2(new_n667), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G229));
  INV_X1    g257(.A(G29), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G32), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n474), .A2(G105), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT95), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT26), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n493), .A2(G141), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n488), .A2(G129), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n693), .A2(KEYINPUT94), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(KEYINPUT94), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n692), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n684), .B1(new_n696), .B2(new_n683), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT27), .B(G1996), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G20), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT23), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n606), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1956), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n683), .A2(G26), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT28), .Z(new_n706));
  OR2_X1    g281(.A1(G104), .A2(G2105), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n707), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT91), .Z(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n488), .B2(G128), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n493), .A2(G140), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(G29), .ZN(new_n713));
  INV_X1    g288(.A(G2067), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n699), .A2(new_n704), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G27), .A2(G29), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G164), .B2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT98), .ZN(new_n719));
  INV_X1    g294(.A(G2078), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(G4), .A2(G16), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT90), .Z(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n601), .B2(new_n700), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1348), .ZN(new_n726));
  NAND2_X1  g301(.A1(G286), .A2(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n700), .A2(G21), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G1966), .ZN(new_n730));
  NOR2_X1   g305(.A1(G16), .A2(G19), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n552), .B2(G16), .ZN(new_n732));
  OAI22_X1  g307(.A1(new_n729), .A2(new_n730), .B1(G1341), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n730), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT31), .B(G11), .ZN(new_n735));
  INV_X1    g310(.A(G28), .ZN(new_n736));
  AOI21_X1  g311(.A(G29), .B1(new_n736), .B2(KEYINPUT30), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(KEYINPUT96), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(KEYINPUT96), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(KEYINPUT30), .B2(new_n736), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n734), .B(new_n735), .C1(new_n738), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n700), .A2(G5), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G171), .B2(new_n700), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1961), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n732), .A2(G1341), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n683), .B2(new_n624), .ZN(new_n746));
  OR4_X1    g321(.A1(new_n733), .A2(new_n741), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n683), .A2(G33), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n493), .A2(G139), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT25), .ZN(new_n751));
  OAI21_X1  g326(.A(G127), .B1(new_n467), .B2(new_n468), .ZN(new_n752));
  INV_X1    g327(.A(G115), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n462), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n751), .B1(new_n754), .B2(G2105), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n748), .B1(new_n757), .B2(new_n683), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(G2072), .Z(new_n759));
  AND2_X1   g334(.A1(KEYINPUT24), .A2(G34), .ZN(new_n760));
  NOR2_X1   g335(.A1(KEYINPUT24), .A2(G34), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n683), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT92), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G160), .B2(G29), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G2084), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT93), .Z(new_n766));
  NOR2_X1   g341(.A1(new_n764), .A2(G2084), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT97), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n759), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G29), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT29), .B(G2090), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n747), .A2(new_n769), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n722), .A2(new_n726), .A3(new_n774), .ZN(new_n775));
  MUX2_X1   g350(.A(G24), .B(G290), .S(G16), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1986), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n493), .A2(G131), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n488), .A2(G119), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n461), .A2(G107), .ZN(new_n780));
  OAI21_X1  g355(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n778), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G29), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G25), .B2(G29), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT35), .B(G1991), .Z(new_n787));
  AOI21_X1  g362(.A(new_n777), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n700), .A2(G6), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n585), .B2(new_n700), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT32), .B(G1981), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n700), .A2(G23), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G288), .B2(G16), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT33), .B(G1976), .Z(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n794), .A2(new_n796), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n700), .A2(G22), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G303), .B2(G16), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1971), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n792), .A2(new_n797), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n791), .B2(new_n790), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n788), .B(new_n805), .C1(new_n786), .C2(new_n787), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n803), .A2(new_n804), .ZN(new_n807));
  OR3_X1    g382(.A1(new_n806), .A2(KEYINPUT36), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT36), .B1(new_n806), .B2(new_n807), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n775), .B1(new_n808), .B2(new_n809), .ZN(G311));
  INV_X1    g385(.A(G311), .ZN(G150));
  NAND2_X1  g386(.A1(new_n602), .A2(G559), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT99), .B(G55), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n520), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n526), .A2(G93), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n815), .B(new_n816), .C1(new_n515), .C2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(new_n551), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n551), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n813), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n823));
  AOI21_X1  g398(.A(G860), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n823), .B2(new_n822), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n818), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT101), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT101), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n825), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(G145));
  INV_X1    g408(.A(new_n507), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT4), .B1(new_n505), .B2(new_n506), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n510), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n501), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n712), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n710), .A2(G164), .A3(new_n711), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n694), .A2(new_n695), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n839), .B(new_n840), .C1(new_n841), .C2(new_n692), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(new_n696), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n757), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n842), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n756), .A2(KEYINPUT102), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n842), .A2(new_n848), .A3(new_n844), .A4(new_n846), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  INV_X1    g428(.A(G118), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n853), .B1(new_n854), .B2(G2105), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(new_n493), .B2(G142), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(new_n488), .B2(G130), .ZN(new_n858));
  AND4_X1   g433(.A1(new_n857), .A2(new_n487), .A3(G130), .A4(G2105), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n617), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n784), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n852), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n624), .B(G160), .Z(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(G162), .Z(new_n866));
  NAND3_X1  g441(.A1(new_n850), .A2(new_n862), .A3(new_n851), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n864), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n866), .B1(new_n864), .B2(new_n867), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT40), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n868), .A2(new_n869), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n874), .A2(new_n875), .A3(new_n871), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n873), .A2(new_n876), .ZN(G395));
  XNOR2_X1  g452(.A(new_n585), .B(G290), .ZN(new_n878));
  XOR2_X1   g453(.A(G288), .B(G303), .Z(new_n879));
  OR2_X1    g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n880), .B(new_n881), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(KEYINPUT105), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(KEYINPUT105), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n821), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n612), .B(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n606), .A2(new_n599), .A3(new_n594), .A4(new_n600), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n601), .A2(G299), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n892), .A2(KEYINPUT41), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(new_n890), .B2(new_n891), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n894), .B1(new_n898), .B2(new_n889), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n887), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n898), .A2(new_n889), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n885), .B(new_n886), .C1(new_n902), .C2(new_n894), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n901), .B1(new_n900), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g480(.A(G868), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G868), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n818), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(G295));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n908), .ZN(G331));
  XOR2_X1   g485(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n911));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  NAND2_X1  g487(.A1(G168), .A2(G171), .ZN(new_n913));
  NAND2_X1  g488(.A1(G286), .A2(G301), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n821), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n913), .A2(new_n819), .A3(new_n820), .A4(new_n914), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(KEYINPUT108), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n915), .A2(new_n821), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n892), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n916), .A2(KEYINPUT107), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n915), .A2(new_n821), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n917), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(new_n895), .B2(new_n897), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n880), .A2(new_n881), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n921), .A2(new_n922), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n923), .A2(new_n928), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n931), .A2(new_n869), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n929), .B(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n923), .A2(new_n928), .A3(new_n930), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n912), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n927), .A2(new_n892), .ZN(new_n939));
  INV_X1    g514(.A(new_n895), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n941));
  INV_X1    g516(.A(new_n897), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n918), .A2(new_n920), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(KEYINPUT111), .B2(new_n897), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n939), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n931), .B(new_n869), .C1(new_n946), .C2(new_n934), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n911), .B1(new_n938), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n932), .A2(new_n912), .A3(new_n937), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(G397));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(G164), .B2(G1384), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n475), .A2(new_n480), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n469), .A2(new_n471), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n956), .B(G40), .C1(new_n957), .C2(new_n461), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n696), .B(G1996), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n712), .B(new_n714), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n784), .A2(new_n787), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n782), .B(KEYINPUT89), .ZN(new_n964));
  INV_X1    g539(.A(new_n787), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n959), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(G290), .A2(G1986), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT112), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n959), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n959), .A2(G1986), .A3(G290), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n973), .A2(KEYINPUT113), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(KEYINPUT113), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n968), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n976), .B(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n572), .A2(new_n573), .A3(G1976), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n503), .A2(new_n509), .ZN(new_n982));
  INV_X1    g557(.A(new_n468), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n983), .B2(new_n466), .ZN(new_n984));
  AND4_X1   g559(.A1(new_n465), .A2(new_n479), .A3(new_n484), .A4(new_n503), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n509), .B1(new_n985), .B2(KEYINPUT75), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n986), .B2(new_n507), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n981), .B1(new_n987), .B2(new_n501), .ZN(new_n988));
  OAI211_X1 g563(.A(G8), .B(new_n980), .C1(new_n988), .C2(new_n958), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT52), .ZN(new_n990));
  INV_X1    g565(.A(G8), .ZN(new_n991));
  INV_X1    g566(.A(G40), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n472), .A2(new_n481), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(G1384), .B1(new_n836), .B2(new_n837), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1976), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(G288), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n980), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n990), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n585), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n526), .A2(G86), .ZN(new_n1002));
  OAI21_X1  g577(.A(G1981), .B1(new_n580), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(KEYINPUT49), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n995), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n999), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n958), .B1(new_n988), .B2(new_n954), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n954), .A2(G1384), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(G164), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT115), .B(new_n1012), .C1(new_n987), .C2(new_n501), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1971), .B1(new_n1010), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2090), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1020), .B(new_n981), .C1(new_n987), .C2(new_n501), .ZN(new_n1021));
  AND4_X1   g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n993), .A4(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(G8), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G303), .A2(G8), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n1024), .B(KEYINPUT55), .Z(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(G8), .B(new_n1025), .C1(new_n1017), .C2(new_n1022), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n838), .A2(new_n1012), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n955), .A2(new_n1029), .A3(new_n993), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n730), .ZN(new_n1031));
  INV_X1    g606(.A(G2084), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1019), .A2(new_n1021), .A3(new_n1032), .A4(new_n993), .ZN(new_n1033));
  AOI211_X1 g608(.A(new_n991), .B(G286), .C1(new_n1031), .C2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1009), .A2(new_n1027), .A3(new_n1028), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT63), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1038), .A2(new_n1004), .A3(new_n995), .ZN(new_n1039));
  INV_X1    g614(.A(new_n999), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1028), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1041), .A2(KEYINPUT63), .A3(new_n1027), .A4(new_n1034), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1037), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1001), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G288), .A2(G1976), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1040), .A2(new_n1039), .ZN(new_n1047));
  OAI22_X1  g622(.A1(new_n1046), .A2(new_n1005), .B1(new_n1047), .B2(new_n1028), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n979), .B1(new_n1043), .B2(new_n1049), .ZN(new_n1050));
  AOI211_X1 g625(.A(KEYINPUT116), .B(new_n1048), .C1(new_n1037), .C2(new_n1042), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G168), .A2(new_n991), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n1053), .B2(KEYINPUT123), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1019), .A2(new_n993), .A3(new_n1021), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1057), .A2(new_n1032), .B1(new_n1030), .B2(new_n730), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1054), .B(new_n1056), .C1(new_n1058), .C2(new_n991), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1056), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1061));
  OAI211_X1 g636(.A(G8), .B(new_n1060), .C1(new_n1061), .C2(G286), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1053), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1059), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1064), .A2(KEYINPUT62), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(KEYINPUT62), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1041), .A2(new_n1027), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1010), .A2(new_n1016), .A3(new_n720), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  INV_X1    g644(.A(G1961), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1019), .A2(new_n1021), .A3(new_n993), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1068), .A2(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1010), .A2(KEYINPUT124), .A3(new_n720), .A4(new_n1029), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n955), .A2(new_n1029), .A3(new_n720), .A4(new_n993), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1076), .A3(KEYINPUT53), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1072), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G171), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1080), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1082));
  NAND2_X1  g657(.A1(G299), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT119), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n606), .A2(KEYINPUT57), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n1086));
  NAND3_X1  g661(.A1(G299), .A2(new_n1086), .A3(new_n1082), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT56), .B(G2072), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1010), .A2(new_n1016), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1956), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT117), .B1(new_n1071), .B2(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1071), .A2(KEYINPUT117), .A3(new_n1091), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1088), .B(new_n1090), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G1348), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n988), .A2(new_n958), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1071), .A2(new_n1096), .B1(new_n1097), .B2(new_n714), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(new_n601), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT120), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1090), .B1(new_n1093), .B2(new_n1092), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1088), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1095), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(KEYINPUT61), .A3(new_n1094), .ZN(new_n1105));
  INV_X1    g680(.A(G1996), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1010), .A2(new_n1016), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n993), .A2(new_n994), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT121), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1112), .A3(new_n1109), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1107), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n552), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT59), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1117), .A3(new_n552), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1105), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1103), .A2(new_n1094), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1097), .A2(new_n714), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1057), .B2(G1348), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n601), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1098), .A2(new_n1127), .A3(KEYINPUT60), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(new_n1098), .B2(KEYINPUT60), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT122), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n602), .B1(new_n1098), .B2(KEYINPUT60), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1098), .A2(new_n1127), .A3(KEYINPUT60), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1121), .A2(new_n1122), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1104), .B1(new_n1120), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1071), .A2(new_n1070), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1010), .A2(new_n1016), .A3(KEYINPUT53), .A4(new_n720), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1137), .A2(G301), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT125), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1072), .A2(new_n1142), .A3(G301), .A4(new_n1139), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1079), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1064), .A2(new_n1027), .A3(new_n1041), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1072), .A2(new_n1139), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1145), .B1(new_n1148), .B2(G171), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(G171), .B2(new_n1078), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1081), .B1(new_n1136), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n978), .B1(new_n1052), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n962), .A2(new_n963), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n712), .A2(G2067), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n959), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n961), .A2(new_n696), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n959), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n959), .A2(new_n1106), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT46), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT47), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1163));
  XNOR2_X1  g738(.A(new_n971), .B(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n968), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1156), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT127), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1153), .A2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g743(.A1(new_n938), .A2(new_n948), .ZN(new_n1170));
  NAND3_X1  g744(.A1(new_n661), .A2(new_n644), .A3(G319), .ZN(new_n1171));
  NOR2_X1   g745(.A1(G229), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g746(.A(new_n1172), .B1(new_n874), .B2(new_n871), .ZN(new_n1173));
  NOR2_X1   g747(.A1(new_n1170), .A2(new_n1173), .ZN(G308));
  OAI221_X1 g748(.A(new_n1172), .B1(new_n871), .B2(new_n874), .C1(new_n938), .C2(new_n948), .ZN(G225));
endmodule


