

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771;

  XNOR2_X1 U371 ( .A(n364), .B(n453), .ZN(n577) );
  XNOR2_X1 U372 ( .A(n462), .B(n461), .ZN(n669) );
  XNOR2_X2 U373 ( .A(G116), .B(G107), .ZN(n518) );
  XNOR2_X2 U374 ( .A(n443), .B(KEYINPUT66), .ZN(n696) );
  XNOR2_X2 U375 ( .A(n476), .B(n444), .ZN(n754) );
  XNOR2_X2 U376 ( .A(n520), .B(KEYINPUT4), .ZN(n476) );
  OR2_X2 U377 ( .A1(n640), .A2(G902), .ZN(n364) );
  AND2_X1 U378 ( .A1(n616), .A2(n615), .ZN(n620) );
  NOR2_X1 U379 ( .A1(n704), .A2(n584), .ZN(n585) );
  INV_X1 U380 ( .A(KEYINPUT0), .ZN(n349) );
  NOR2_X1 U381 ( .A1(n660), .A2(n674), .ZN(n661) );
  NOR2_X1 U382 ( .A1(n650), .A2(n674), .ZN(n651) );
  NOR2_X1 U383 ( .A1(n643), .A2(n674), .ZN(n646) );
  BUF_X1 U384 ( .A(n652), .Z(n668) );
  NOR2_X1 U385 ( .A1(n620), .A2(n422), .ZN(n421) );
  NOR2_X1 U386 ( .A1(n620), .A2(n623), .ZN(n418) );
  XNOR2_X1 U387 ( .A(n560), .B(KEYINPUT81), .ZN(n561) );
  AND2_X1 U388 ( .A1(n637), .A2(n636), .ZN(n541) );
  NAND2_X1 U389 ( .A1(n351), .A2(n407), .ZN(n637) );
  BUF_X1 U390 ( .A(n636), .Z(n350) );
  XNOR2_X1 U391 ( .A(n410), .B(n536), .ZN(n636) );
  NAND2_X1 U392 ( .A1(n404), .A2(n402), .ZN(n594) );
  AND2_X1 U393 ( .A1(n406), .A2(n405), .ZN(n404) );
  OR2_X1 U394 ( .A1(n553), .A2(n552), .ZN(n583) );
  INV_X1 U395 ( .A(n580), .ZN(n347) );
  XNOR2_X1 U396 ( .A(n440), .B(n439), .ZN(n567) );
  XNOR2_X1 U397 ( .A(n426), .B(G119), .ZN(n470) );
  XNOR2_X1 U398 ( .A(KEYINPUT69), .B(KEYINPUT3), .ZN(n445) );
  XNOR2_X2 U399 ( .A(n496), .B(n349), .ZN(n348) );
  NAND2_X1 U400 ( .A1(n421), .A2(n417), .ZN(n420) );
  XNOR2_X2 U401 ( .A(n465), .B(n464), .ZN(n545) );
  NOR2_X2 U402 ( .A1(G902), .A2(n669), .ZN(n465) );
  INV_X1 U403 ( .A(n768), .ZN(n378) );
  XNOR2_X1 U404 ( .A(G146), .B(G125), .ZN(n479) );
  NAND2_X1 U405 ( .A1(n572), .A2(n688), .ZN(n607) );
  XNOR2_X1 U406 ( .A(n582), .B(n401), .ZN(n605) );
  INV_X1 U407 ( .A(KEYINPUT39), .ZN(n401) );
  NAND2_X1 U408 ( .A1(n533), .A2(n413), .ZN(n409) );
  NOR2_X1 U409 ( .A1(n610), .A2(n414), .ZN(n413) );
  XNOR2_X1 U410 ( .A(KEYINPUT5), .B(G119), .ZN(n447) );
  XOR2_X1 U411 ( .A(G116), .B(G137), .Z(n448) );
  NAND2_X1 U412 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U413 ( .A1(n375), .A2(n374), .ZN(n370) );
  NOR2_X1 U414 ( .A1(n378), .A2(n377), .ZN(n374) );
  XNOR2_X1 U415 ( .A(G113), .B(G101), .ZN(n446) );
  INV_X1 U416 ( .A(G110), .ZN(n426) );
  XNOR2_X1 U417 ( .A(G122), .B(G104), .ZN(n506) );
  NOR2_X1 U418 ( .A1(G953), .A2(G237), .ZN(n501) );
  XNOR2_X1 U419 ( .A(G131), .B(G143), .ZN(n507) );
  XNOR2_X1 U420 ( .A(KEYINPUT67), .B(KEYINPUT10), .ZN(n435) );
  INV_X1 U421 ( .A(KEYINPUT40), .ZN(n398) );
  NOR2_X1 U422 ( .A1(n583), .A2(n398), .ZN(n394) );
  NAND2_X1 U423 ( .A1(n389), .A2(n358), .ZN(n388) );
  XNOR2_X1 U424 ( .A(n607), .B(KEYINPUT103), .ZN(n389) );
  INV_X1 U425 ( .A(KEYINPUT36), .ZN(n387) );
  NOR2_X1 U426 ( .A1(n696), .A2(n390), .ZN(n578) );
  XNOR2_X1 U427 ( .A(n391), .B(KEYINPUT30), .ZN(n390) );
  NAND2_X1 U428 ( .A1(n363), .A2(n362), .ZN(n391) );
  INV_X1 U429 ( .A(KEYINPUT97), .ZN(n414) );
  NOR2_X1 U430 ( .A1(n354), .A2(n412), .ZN(n411) );
  NOR2_X1 U431 ( .A1(n695), .A2(KEYINPUT97), .ZN(n412) );
  NAND2_X1 U432 ( .A1(n348), .A2(n353), .ZN(n532) );
  XNOR2_X1 U433 ( .A(KEYINPUT18), .B(KEYINPUT76), .ZN(n474) );
  XNOR2_X1 U434 ( .A(KEYINPUT84), .B(KEYINPUT75), .ZN(n473) );
  NAND2_X1 U435 ( .A1(n419), .A2(KEYINPUT79), .ZN(n415) );
  NOR2_X1 U436 ( .A1(n579), .A2(n567), .ZN(n568) );
  INV_X1 U437 ( .A(n577), .ZN(n363) );
  XNOR2_X1 U438 ( .A(n463), .B(KEYINPUT68), .ZN(n464) );
  XNOR2_X1 U439 ( .A(n462), .B(n452), .ZN(n640) );
  AND2_X1 U440 ( .A1(n638), .A2(n614), .ZN(n368) );
  XNOR2_X1 U441 ( .A(G128), .B(KEYINPUT90), .ZN(n427) );
  XNOR2_X1 U442 ( .A(KEYINPUT89), .B(KEYINPUT74), .ZN(n428) );
  XNOR2_X1 U443 ( .A(G134), .B(G122), .ZN(n519) );
  XNOR2_X1 U444 ( .A(G101), .B(G110), .ZN(n455) );
  XOR2_X1 U445 ( .A(G104), .B(G107), .Z(n456) );
  XOR2_X1 U446 ( .A(G137), .B(G140), .Z(n458) );
  INV_X1 U447 ( .A(n347), .ZN(n613) );
  XNOR2_X1 U448 ( .A(n589), .B(n400), .ZN(n694) );
  INV_X1 U449 ( .A(KEYINPUT41), .ZN(n400) );
  NAND2_X1 U450 ( .A1(n347), .A2(n403), .ZN(n402) );
  AND2_X1 U451 ( .A1(n348), .A2(n466), .ZN(n548) );
  BUF_X1 U452 ( .A(n577), .Z(n704) );
  BUF_X1 U453 ( .A(n567), .Z(n555) );
  XNOR2_X1 U454 ( .A(n512), .B(n511), .ZN(n647) );
  XNOR2_X1 U455 ( .A(n510), .B(n509), .ZN(n511) );
  NOR2_X1 U456 ( .A1(n761), .A2(G952), .ZN(n674) );
  XNOR2_X1 U457 ( .A(n399), .B(KEYINPUT42), .ZN(n766) );
  NOR2_X1 U458 ( .A1(n694), .A2(n596), .ZN(n399) );
  NAND2_X1 U459 ( .A1(n395), .A2(n393), .ZN(n771) );
  AND2_X1 U460 ( .A1(n397), .A2(n396), .ZN(n395) );
  NAND2_X1 U461 ( .A1(n392), .A2(n394), .ZN(n393) );
  XNOR2_X1 U462 ( .A(n576), .B(KEYINPUT104), .ZN(n768) );
  XNOR2_X1 U463 ( .A(n388), .B(n387), .ZN(n575) );
  AND2_X1 U464 ( .A1(n365), .A2(n357), .ZN(n686) );
  XNOR2_X1 U465 ( .A(n367), .B(n366), .ZN(n365) );
  INV_X1 U466 ( .A(KEYINPUT102), .ZN(n366) );
  NAND2_X1 U467 ( .A1(n408), .A2(n414), .ZN(n407) );
  AND2_X1 U468 ( .A1(n409), .A2(n411), .ZN(n351) );
  NOR2_X1 U469 ( .A1(n704), .A2(n695), .ZN(n352) );
  AND2_X1 U470 ( .A1(n715), .A2(n698), .ZN(n353) );
  NOR2_X1 U471 ( .A1(n624), .A2(n618), .ZN(n619) );
  NAND2_X1 U472 ( .A1(n704), .A2(n699), .ZN(n354) );
  AND2_X1 U473 ( .A1(n569), .A2(n535), .ZN(n355) );
  AND2_X1 U474 ( .A1(n569), .A2(n556), .ZN(n356) );
  NOR2_X1 U475 ( .A1(n553), .A2(n551), .ZN(n357) );
  AND2_X1 U476 ( .A1(n347), .A2(n362), .ZN(n358) );
  AND2_X1 U477 ( .A1(n347), .A2(n593), .ZN(n359) );
  XOR2_X1 U478 ( .A(n531), .B(KEYINPUT22), .Z(n360) );
  INV_X1 U479 ( .A(n623), .ZN(n419) );
  INV_X1 U480 ( .A(KEYINPUT79), .ZN(n422) );
  NOR2_X1 U481 ( .A1(n714), .A2(n713), .ZN(n718) );
  INV_X1 U482 ( .A(n713), .ZN(n362) );
  NAND2_X1 U483 ( .A1(n713), .A2(KEYINPUT19), .ZN(n405) );
  NOR2_X1 U484 ( .A1(n713), .A2(KEYINPUT19), .ZN(n403) );
  NAND2_X1 U485 ( .A1(n361), .A2(n420), .ZN(n423) );
  NAND2_X1 U486 ( .A1(n416), .A2(n415), .ZN(n361) );
  NAND2_X1 U487 ( .A1(n369), .A2(n368), .ZN(n759) );
  NOR2_X1 U488 ( .A1(n771), .A2(n766), .ZN(n590) );
  XNOR2_X2 U489 ( .A(n379), .B(n485), .ZN(n580) );
  AND2_X2 U490 ( .A1(n424), .A2(n423), .ZN(n652) );
  NAND2_X1 U491 ( .A1(n592), .A2(n359), .ZN(n367) );
  XNOR2_X1 U492 ( .A(n612), .B(KEYINPUT101), .ZN(n373) );
  NAND2_X1 U493 ( .A1(n373), .A2(n613), .ZN(n638) );
  NAND2_X1 U494 ( .A1(n371), .A2(n370), .ZN(n369) );
  AND2_X1 U495 ( .A1(n372), .A2(n376), .ZN(n371) );
  NAND2_X1 U496 ( .A1(n383), .A2(n377), .ZN(n372) );
  INV_X1 U497 ( .A(n383), .ZN(n375) );
  INV_X1 U498 ( .A(KEYINPUT48), .ZN(n377) );
  NAND2_X1 U499 ( .A1(n594), .A2(n495), .ZN(n496) );
  OR2_X2 U500 ( .A1(n653), .A2(n621), .ZN(n379) );
  XNOR2_X1 U501 ( .A(n380), .B(n744), .ZN(n653) );
  XNOR2_X1 U502 ( .A(n482), .B(n481), .ZN(n380) );
  XNOR2_X1 U503 ( .A(n472), .B(n471), .ZN(n744) );
  NAND2_X1 U504 ( .A1(n541), .A2(n663), .ZN(n537) );
  NAND2_X1 U505 ( .A1(n533), .A2(n355), .ZN(n410) );
  NAND2_X1 U506 ( .A1(n533), .A2(n356), .ZN(n630) );
  XNOR2_X2 U507 ( .A(n532), .B(n360), .ZN(n533) );
  NAND2_X1 U508 ( .A1(n466), .A2(n381), .ZN(n467) );
  NOR2_X1 U509 ( .A1(n382), .A2(n569), .ZN(n381) );
  INV_X1 U510 ( .A(n610), .ZN(n382) );
  XNOR2_X2 U511 ( .A(n545), .B(KEYINPUT1), .ZN(n610) );
  NAND2_X1 U512 ( .A1(n384), .A2(n591), .ZN(n383) );
  AND2_X1 U513 ( .A1(n604), .A2(n385), .ZN(n384) );
  XNOR2_X1 U514 ( .A(n686), .B(n386), .ZN(n385) );
  INV_X1 U515 ( .A(KEYINPUT78), .ZN(n386) );
  INV_X1 U516 ( .A(n605), .ZN(n392) );
  NAND2_X1 U517 ( .A1(n583), .A2(n398), .ZN(n396) );
  NAND2_X1 U518 ( .A1(n605), .A2(n398), .ZN(n397) );
  XNOR2_X1 U519 ( .A(n434), .B(n433), .ZN(n436) );
  NAND2_X1 U520 ( .A1(n580), .A2(KEYINPUT19), .ZN(n406) );
  INV_X1 U521 ( .A(n533), .ZN(n408) );
  INV_X1 U522 ( .A(n693), .ZN(n424) );
  NAND2_X1 U523 ( .A1(n418), .A2(n417), .ZN(n416) );
  INV_X1 U524 ( .A(n619), .ZN(n417) );
  AND2_X1 U525 ( .A1(G217), .A2(n441), .ZN(n425) );
  INV_X1 U526 ( .A(KEYINPUT99), .ZN(n570) );
  BUF_X1 U527 ( .A(n653), .Z(n657) );
  INV_X1 U528 ( .A(n674), .ZN(n628) );
  XNOR2_X1 U529 ( .A(n470), .B(n427), .ZN(n431) );
  XOR2_X1 U530 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n429) );
  XNOR2_X1 U531 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U532 ( .A(n431), .B(n430), .ZN(n434) );
  INV_X2 U533 ( .A(G953), .ZN(n761) );
  NAND2_X1 U534 ( .A1(G234), .A2(n761), .ZN(n432) );
  XOR2_X1 U535 ( .A(KEYINPUT8), .B(n432), .Z(n515) );
  NAND2_X1 U536 ( .A1(G221), .A2(n515), .ZN(n433) );
  XNOR2_X1 U537 ( .A(n435), .B(n479), .ZN(n509) );
  XNOR2_X1 U538 ( .A(n509), .B(n458), .ZN(n751) );
  XNOR2_X1 U539 ( .A(n436), .B(n751), .ZN(n626) );
  INV_X1 U540 ( .A(G902), .ZN(n525) );
  NAND2_X1 U541 ( .A1(n626), .A2(n525), .ZN(n440) );
  XOR2_X1 U542 ( .A(KEYINPUT25), .B(KEYINPUT91), .Z(n438) );
  XNOR2_X1 U543 ( .A(G902), .B(KEYINPUT15), .ZN(n483) );
  NAND2_X1 U544 ( .A1(n483), .A2(G234), .ZN(n437) );
  XNOR2_X1 U545 ( .A(n437), .B(KEYINPUT20), .ZN(n441) );
  XNOR2_X1 U546 ( .A(n438), .B(n425), .ZN(n439) );
  AND2_X1 U547 ( .A1(n441), .A2(G221), .ZN(n442) );
  XNOR2_X1 U548 ( .A(n442), .B(KEYINPUT21), .ZN(n698) );
  NAND2_X1 U549 ( .A1(n567), .A2(n698), .ZN(n443) );
  INV_X1 U550 ( .A(n696), .ZN(n466) );
  XNOR2_X2 U551 ( .A(G143), .B(G128), .ZN(n520) );
  XNOR2_X1 U552 ( .A(G131), .B(G134), .ZN(n444) );
  XNOR2_X2 U553 ( .A(n754), .B(G146), .ZN(n462) );
  XNOR2_X1 U554 ( .A(n446), .B(n445), .ZN(n469) );
  XNOR2_X1 U555 ( .A(n448), .B(n447), .ZN(n450) );
  NAND2_X1 U556 ( .A1(n501), .A2(G210), .ZN(n449) );
  XNOR2_X1 U557 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U558 ( .A(n469), .B(n451), .ZN(n452) );
  INV_X1 U559 ( .A(G472), .ZN(n453) );
  INV_X1 U560 ( .A(KEYINPUT6), .ZN(n454) );
  XNOR2_X1 U561 ( .A(n577), .B(n454), .ZN(n569) );
  XNOR2_X1 U562 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U563 ( .A(n458), .B(n457), .ZN(n460) );
  AND2_X1 U564 ( .A1(G227), .A2(n761), .ZN(n459) );
  XNOR2_X1 U565 ( .A(n460), .B(n459), .ZN(n461) );
  INV_X1 U566 ( .A(G469), .ZN(n463) );
  XNOR2_X2 U567 ( .A(n467), .B(KEYINPUT33), .ZN(n729) );
  XNOR2_X1 U568 ( .A(n518), .B(KEYINPUT16), .ZN(n468) );
  XNOR2_X1 U569 ( .A(n469), .B(n468), .ZN(n472) );
  XNOR2_X1 U570 ( .A(n470), .B(n506), .ZN(n471) );
  XNOR2_X1 U571 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U572 ( .A(n476), .B(n475), .ZN(n482) );
  NAND2_X1 U573 ( .A1(n761), .A2(G224), .ZN(n478) );
  XNOR2_X1 U574 ( .A(KEYINPUT87), .B(KEYINPUT17), .ZN(n477) );
  XNOR2_X1 U575 ( .A(n478), .B(n477), .ZN(n480) );
  XNOR2_X1 U576 ( .A(n480), .B(n479), .ZN(n481) );
  INV_X1 U577 ( .A(n483), .ZN(n621) );
  INV_X1 U578 ( .A(G237), .ZN(n484) );
  NAND2_X1 U579 ( .A1(n525), .A2(n484), .ZN(n486) );
  NAND2_X1 U580 ( .A1(n486), .A2(G210), .ZN(n485) );
  NAND2_X1 U581 ( .A1(n486), .A2(G214), .ZN(n488) );
  INV_X1 U582 ( .A(KEYINPUT88), .ZN(n487) );
  XNOR2_X1 U583 ( .A(n488), .B(n487), .ZN(n713) );
  NAND2_X1 U584 ( .A1(G234), .A2(G237), .ZN(n489) );
  XNOR2_X1 U585 ( .A(n489), .B(KEYINPUT14), .ZN(n490) );
  XNOR2_X1 U586 ( .A(KEYINPUT72), .B(n490), .ZN(n491) );
  NAND2_X1 U587 ( .A1(G952), .A2(n491), .ZN(n727) );
  NOR2_X1 U588 ( .A1(n727), .A2(G953), .ZN(n566) );
  INV_X1 U589 ( .A(n566), .ZN(n494) );
  AND2_X1 U590 ( .A1(n491), .A2(G953), .ZN(n492) );
  NAND2_X1 U591 ( .A1(G902), .A2(n492), .ZN(n564) );
  OR2_X1 U592 ( .A1(n564), .A2(G898), .ZN(n493) );
  NAND2_X1 U593 ( .A1(n494), .A2(n493), .ZN(n495) );
  NAND2_X1 U594 ( .A1(n729), .A2(n348), .ZN(n498) );
  INV_X1 U595 ( .A(KEYINPUT34), .ZN(n497) );
  XNOR2_X1 U596 ( .A(n498), .B(n497), .ZN(n528) );
  XOR2_X1 U597 ( .A(KEYINPUT94), .B(KEYINPUT11), .Z(n500) );
  XNOR2_X1 U598 ( .A(G113), .B(G140), .ZN(n499) );
  XNOR2_X1 U599 ( .A(n500), .B(n499), .ZN(n505) );
  NAND2_X1 U600 ( .A1(G214), .A2(n501), .ZN(n503) );
  XOR2_X1 U601 ( .A(KEYINPUT95), .B(KEYINPUT12), .Z(n502) );
  XNOR2_X1 U602 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U603 ( .A(n505), .B(n504), .Z(n512) );
  INV_X1 U604 ( .A(n506), .ZN(n508) );
  XNOR2_X1 U605 ( .A(n508), .B(n507), .ZN(n510) );
  NAND2_X1 U606 ( .A1(n647), .A2(n525), .ZN(n514) );
  XNOR2_X1 U607 ( .A(KEYINPUT13), .B(G475), .ZN(n513) );
  XNOR2_X1 U608 ( .A(n514), .B(n513), .ZN(n553) );
  XOR2_X1 U609 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n517) );
  NAND2_X1 U610 ( .A1(G217), .A2(n515), .ZN(n516) );
  XNOR2_X1 U611 ( .A(n517), .B(n516), .ZN(n524) );
  XNOR2_X1 U612 ( .A(n518), .B(n519), .ZN(n522) );
  XNOR2_X1 U613 ( .A(n520), .B(KEYINPUT96), .ZN(n521) );
  XNOR2_X1 U614 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U615 ( .A(n524), .B(n523), .ZN(n664) );
  NAND2_X1 U616 ( .A1(n664), .A2(n525), .ZN(n527) );
  INV_X1 U617 ( .A(G478), .ZN(n526) );
  XNOR2_X1 U618 ( .A(n527), .B(n526), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n528), .A2(n357), .ZN(n530) );
  INV_X1 U620 ( .A(KEYINPUT35), .ZN(n529) );
  XNOR2_X2 U621 ( .A(n530), .B(n529), .ZN(n663) );
  AND2_X1 U622 ( .A1(n553), .A2(n551), .ZN(n715) );
  INV_X1 U623 ( .A(KEYINPUT71), .ZN(n531) );
  INV_X1 U624 ( .A(n610), .ZN(n695) );
  INV_X1 U625 ( .A(n555), .ZN(n699) );
  INV_X1 U626 ( .A(KEYINPUT86), .ZN(n534) );
  XNOR2_X1 U627 ( .A(n610), .B(n534), .ZN(n573) );
  NOR2_X1 U628 ( .A1(n555), .A2(n573), .ZN(n535) );
  XNOR2_X1 U629 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n536) );
  XNOR2_X1 U630 ( .A(n537), .B(KEYINPUT70), .ZN(n539) );
  INV_X1 U631 ( .A(KEYINPUT44), .ZN(n538) );
  NAND2_X1 U632 ( .A1(n539), .A2(n538), .ZN(n543) );
  AND2_X1 U633 ( .A1(KEYINPUT70), .A2(KEYINPUT44), .ZN(n540) );
  NAND2_X1 U634 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U635 ( .A1(n543), .A2(n542), .ZN(n562) );
  INV_X1 U636 ( .A(n663), .ZN(n544) );
  NAND2_X1 U637 ( .A1(n544), .A2(KEYINPUT44), .ZN(n559) );
  BUF_X1 U638 ( .A(n545), .Z(n586) );
  AND2_X1 U639 ( .A1(n704), .A2(n586), .ZN(n546) );
  NAND2_X1 U640 ( .A1(n548), .A2(n546), .ZN(n547) );
  XNOR2_X1 U641 ( .A(n547), .B(KEYINPUT92), .ZN(n676) );
  NAND2_X1 U642 ( .A1(n548), .A2(n352), .ZN(n550) );
  XNOR2_X1 U643 ( .A(KEYINPUT93), .B(KEYINPUT31), .ZN(n549) );
  XNOR2_X1 U644 ( .A(n550), .B(n549), .ZN(n634) );
  NAND2_X1 U645 ( .A1(n676), .A2(n634), .ZN(n554) );
  INV_X1 U646 ( .A(n551), .ZN(n552) );
  NAND2_X1 U647 ( .A1(n553), .A2(n552), .ZN(n680) );
  NAND2_X1 U648 ( .A1(n680), .A2(n583), .ZN(n717) );
  NAND2_X1 U649 ( .A1(n554), .A2(n717), .ZN(n557) );
  AND2_X1 U650 ( .A1(n555), .A2(n695), .ZN(n556) );
  AND2_X1 U651 ( .A1(n557), .A2(n630), .ZN(n558) );
  NAND2_X1 U652 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U653 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X2 U654 ( .A(n563), .B(KEYINPUT45), .ZN(n738) );
  NAND2_X1 U655 ( .A1(n738), .A2(n621), .ZN(n616) );
  NOR2_X1 U656 ( .A1(G900), .A2(n564), .ZN(n565) );
  NOR2_X1 U657 ( .A1(n566), .A2(n565), .ZN(n579) );
  NAND2_X1 U658 ( .A1(n568), .A2(n698), .ZN(n584) );
  NOR2_X1 U659 ( .A1(n569), .A2(n584), .ZN(n571) );
  XNOR2_X1 U660 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U661 ( .A(n583), .B(KEYINPUT98), .ZN(n687) );
  INV_X1 U662 ( .A(n573), .ZN(n574) );
  NAND2_X1 U663 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U664 ( .A1(n578), .A2(n586), .ZN(n592) );
  INV_X1 U665 ( .A(n579), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n613), .B(KEYINPUT38), .ZN(n588) );
  AND2_X1 U667 ( .A1(n593), .A2(n588), .ZN(n581) );
  NAND2_X1 U668 ( .A1(n592), .A2(n581), .ZN(n582) );
  XNOR2_X1 U669 ( .A(n585), .B(KEYINPUT28), .ZN(n587) );
  NAND2_X1 U670 ( .A1(n587), .A2(n586), .ZN(n596) );
  INV_X1 U671 ( .A(n588), .ZN(n714) );
  NAND2_X1 U672 ( .A1(n718), .A2(n715), .ZN(n589) );
  XNOR2_X1 U673 ( .A(n590), .B(KEYINPUT46), .ZN(n591) );
  INV_X1 U674 ( .A(n594), .ZN(n595) );
  NOR2_X1 U675 ( .A1(n596), .A2(n595), .ZN(n689) );
  INV_X1 U676 ( .A(KEYINPUT47), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n689), .A2(n601), .ZN(n597) );
  XNOR2_X1 U678 ( .A(n597), .B(KEYINPUT77), .ZN(n600) );
  AND2_X1 U679 ( .A1(n717), .A2(n601), .ZN(n598) );
  NAND2_X1 U680 ( .A1(n689), .A2(n598), .ZN(n599) );
  NAND2_X1 U681 ( .A1(n600), .A2(n599), .ZN(n603) );
  NOR2_X1 U682 ( .A1(n601), .A2(n717), .ZN(n602) );
  NOR2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n604) );
  OR2_X1 U684 ( .A1(n680), .A2(n605), .ZN(n606) );
  XNOR2_X1 U685 ( .A(n606), .B(KEYINPUT105), .ZN(n767) );
  INV_X1 U686 ( .A(n767), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n713), .A2(n607), .ZN(n608) );
  XOR2_X1 U688 ( .A(KEYINPUT100), .B(n608), .Z(n609) );
  NOR2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U690 ( .A(KEYINPUT43), .B(n611), .ZN(n612) );
  NOR2_X1 U691 ( .A1(n759), .A2(KEYINPUT80), .ZN(n615) );
  INV_X1 U692 ( .A(n759), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n617), .A2(n738), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n621), .A2(KEYINPUT80), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n621), .A2(KEYINPUT2), .ZN(n622) );
  XNOR2_X1 U696 ( .A(n622), .B(KEYINPUT65), .ZN(n623) );
  INV_X1 U697 ( .A(n624), .ZN(n691) );
  NAND2_X1 U698 ( .A1(n691), .A2(KEYINPUT2), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n625), .B(KEYINPUT73), .ZN(n693) );
  NAND2_X1 U700 ( .A1(n668), .A2(G217), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(n626), .ZN(n629) );
  AND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(G66) );
  XNOR2_X1 U703 ( .A(n630), .B(G101), .ZN(G3) );
  NOR2_X1 U704 ( .A1(n634), .A2(n680), .ZN(n632) );
  XNOR2_X1 U705 ( .A(G116), .B(KEYINPUT109), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n632), .B(n631), .ZN(G18) );
  NOR2_X1 U707 ( .A1(n676), .A2(n687), .ZN(n633) );
  XOR2_X1 U708 ( .A(G104), .B(n633), .Z(G6) );
  NOR2_X1 U709 ( .A1(n634), .A2(n687), .ZN(n635) );
  XOR2_X1 U710 ( .A(G113), .B(n635), .Z(G15) );
  XNOR2_X1 U711 ( .A(n350), .B(G119), .ZN(G21) );
  XNOR2_X1 U712 ( .A(n637), .B(G110), .ZN(G12) );
  XNOR2_X1 U713 ( .A(n638), .B(G140), .ZN(G42) );
  NAND2_X1 U714 ( .A1(n652), .A2(G472), .ZN(n642) );
  XOR2_X1 U715 ( .A(KEYINPUT85), .B(KEYINPUT62), .Z(n639) );
  XNOR2_X1 U716 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U718 ( .A(KEYINPUT106), .B(KEYINPUT63), .ZN(n644) );
  XOR2_X1 U719 ( .A(n644), .B(KEYINPUT82), .Z(n645) );
  XNOR2_X1 U720 ( .A(n646), .B(n645), .ZN(G57) );
  NAND2_X1 U721 ( .A1(n652), .A2(G475), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n647), .B(KEYINPUT59), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n651), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U725 ( .A1(n652), .A2(G210), .ZN(n659) );
  XOR2_X1 U726 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n655) );
  XNOR2_X1 U727 ( .A(KEYINPUT55), .B(KEYINPUT83), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U732 ( .A(G122), .B(KEYINPUT125), .Z(n662) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(G24) );
  NAND2_X1 U734 ( .A1(n668), .A2(G478), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n664), .B(KEYINPUT119), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n666), .B(n665), .ZN(n667) );
  NOR2_X1 U737 ( .A1(n667), .A2(n674), .ZN(G63) );
  NAND2_X1 U738 ( .A1(n668), .A2(G469), .ZN(n673) );
  XOR2_X1 U739 ( .A(KEYINPUT118), .B(KEYINPUT57), .Z(n670) );
  XNOR2_X1 U740 ( .A(n670), .B(KEYINPUT58), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n669), .B(n671), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n673), .B(n672), .ZN(n675) );
  NOR2_X1 U743 ( .A1(n675), .A2(n674), .ZN(G54) );
  NOR2_X1 U744 ( .A1(n676), .A2(n680), .ZN(n678) );
  XNOR2_X1 U745 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U747 ( .A(G107), .B(n679), .ZN(G9) );
  XOR2_X1 U748 ( .A(KEYINPUT108), .B(KEYINPUT29), .Z(n683) );
  INV_X1 U749 ( .A(n680), .ZN(n681) );
  NAND2_X1 U750 ( .A1(n689), .A2(n681), .ZN(n682) );
  XNOR2_X1 U751 ( .A(n683), .B(n682), .ZN(n685) );
  XOR2_X1 U752 ( .A(G128), .B(KEYINPUT107), .Z(n684) );
  XNOR2_X1 U753 ( .A(n685), .B(n684), .ZN(G30) );
  XOR2_X1 U754 ( .A(G143), .B(n686), .Z(G45) );
  INV_X1 U755 ( .A(n687), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U757 ( .A(n690), .B(G146), .ZN(G48) );
  NOR2_X1 U758 ( .A1(n691), .A2(KEYINPUT2), .ZN(n692) );
  NOR2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n736) );
  INV_X1 U760 ( .A(n694), .ZN(n728) );
  NAND2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U762 ( .A(KEYINPUT50), .B(n697), .ZN(n708) );
  INV_X1 U763 ( .A(n698), .ZN(n700) );
  NAND2_X1 U764 ( .A1(n700), .A2(n699), .ZN(n703) );
  XNOR2_X1 U765 ( .A(KEYINPUT49), .B(KEYINPUT112), .ZN(n701) );
  XNOR2_X1 U766 ( .A(n701), .B(KEYINPUT111), .ZN(n702) );
  XNOR2_X1 U767 ( .A(n703), .B(n702), .ZN(n705) );
  NAND2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U769 ( .A(KEYINPUT113), .B(n706), .ZN(n707) );
  NAND2_X1 U770 ( .A1(n708), .A2(n707), .ZN(n710) );
  NAND2_X1 U771 ( .A1(n352), .A2(n466), .ZN(n709) );
  NAND2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U773 ( .A(KEYINPUT51), .B(n711), .Z(n712) );
  NAND2_X1 U774 ( .A1(n728), .A2(n712), .ZN(n724) );
  NAND2_X1 U775 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U776 ( .A1(n716), .A2(n715), .ZN(n721) );
  NAND2_X1 U777 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U778 ( .A(KEYINPUT114), .B(n719), .ZN(n720) );
  NAND2_X1 U779 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U780 ( .A1(n729), .A2(n722), .ZN(n723) );
  NAND2_X1 U781 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U782 ( .A(KEYINPUT52), .B(n725), .Z(n726) );
  NOR2_X1 U783 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U784 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U785 ( .A(KEYINPUT115), .B(n730), .Z(n731) );
  NOR2_X1 U786 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U787 ( .A(n733), .B(KEYINPUT116), .ZN(n734) );
  NAND2_X1 U788 ( .A1(n734), .A2(n761), .ZN(n735) );
  NOR2_X1 U789 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U790 ( .A(KEYINPUT53), .B(n737), .ZN(G75) );
  INV_X1 U791 ( .A(n738), .ZN(n739) );
  NOR2_X1 U792 ( .A1(n739), .A2(G953), .ZN(n743) );
  INV_X1 U793 ( .A(G898), .ZN(n745) );
  NAND2_X1 U794 ( .A1(G953), .A2(G224), .ZN(n740) );
  XOR2_X1 U795 ( .A(KEYINPUT61), .B(n740), .Z(n741) );
  NOR2_X1 U796 ( .A1(n745), .A2(n741), .ZN(n742) );
  NOR2_X1 U797 ( .A1(n743), .A2(n742), .ZN(n750) );
  INV_X1 U798 ( .A(n744), .ZN(n747) );
  NAND2_X1 U799 ( .A1(n745), .A2(G953), .ZN(n746) );
  NAND2_X1 U800 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n748), .B(KEYINPUT120), .ZN(n749) );
  XNOR2_X1 U802 ( .A(n750), .B(n749), .ZN(G69) );
  XOR2_X1 U803 ( .A(n751), .B(KEYINPUT121), .Z(n752) );
  XNOR2_X1 U804 ( .A(KEYINPUT122), .B(n752), .ZN(n753) );
  XNOR2_X1 U805 ( .A(n754), .B(n753), .ZN(n758) );
  XOR2_X1 U806 ( .A(G227), .B(n758), .Z(n755) );
  NAND2_X1 U807 ( .A1(n755), .A2(G900), .ZN(n756) );
  NAND2_X1 U808 ( .A1(G953), .A2(n756), .ZN(n757) );
  XNOR2_X1 U809 ( .A(n757), .B(KEYINPUT124), .ZN(n764) );
  XNOR2_X1 U810 ( .A(KEYINPUT123), .B(n758), .ZN(n760) );
  XNOR2_X1 U811 ( .A(n760), .B(n759), .ZN(n762) );
  NAND2_X1 U812 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U813 ( .A1(n764), .A2(n763), .ZN(G72) );
  XOR2_X1 U814 ( .A(G137), .B(KEYINPUT126), .Z(n765) );
  XNOR2_X1 U815 ( .A(n766), .B(n765), .ZN(G39) );
  XOR2_X1 U816 ( .A(G134), .B(n767), .Z(G36) );
  XOR2_X1 U817 ( .A(KEYINPUT110), .B(KEYINPUT37), .Z(n770) );
  XNOR2_X1 U818 ( .A(G125), .B(n768), .ZN(n769) );
  XNOR2_X1 U819 ( .A(n770), .B(n769), .ZN(G27) );
  XOR2_X1 U820 ( .A(n771), .B(G131), .Z(G33) );
endmodule

