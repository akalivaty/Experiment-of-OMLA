//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n191), .A2(G143), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n195), .A2(new_n196), .B1(KEYINPUT1), .B2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  OR2_X1    g016(.A1(KEYINPUT74), .A2(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT74), .A2(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT0), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(new_n196), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n195), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n199), .B1(new_n209), .B2(new_n196), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(new_n205), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G224), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n214), .B(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT2), .B(G113), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT64), .B(G119), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G116), .ZN(new_n221));
  INV_X1    g035(.A(G119), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT65), .B1(new_n222), .B2(G116), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  INV_X1    g038(.A(G116), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n219), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n221), .A2(new_n227), .A3(new_n219), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G107), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT83), .B1(new_n232), .B2(G104), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT83), .ZN(new_n234));
  INV_X1    g048(.A(G104), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(G107), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n235), .A2(KEYINPUT3), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n232), .A2(KEYINPUT82), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G107), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n232), .A2(G104), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT3), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n237), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(G101), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n231), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G101), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n237), .A2(new_n242), .A3(new_n249), .A4(new_n244), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT84), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT3), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(G104), .B2(new_n232), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT82), .B(G107), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(new_n238), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT84), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n255), .A2(new_n256), .A3(new_n249), .A4(new_n237), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n246), .B1(new_n245), .B2(G101), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n258), .A2(KEYINPUT85), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT85), .B1(new_n258), .B2(new_n259), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n248), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n243), .B1(new_n254), .B2(G104), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n251), .A2(new_n257), .B1(G101), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n221), .A2(KEYINPUT5), .A3(new_n227), .ZN(new_n266));
  OAI21_X1  g080(.A(G113), .B1(new_n221), .B2(KEYINPUT5), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n230), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(G110), .B(G122), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n270), .A2(new_n272), .B1(KEYINPUT90), .B2(KEYINPUT6), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT90), .A2(KEYINPUT6), .ZN(new_n274));
  AOI211_X1 g088(.A(new_n271), .B(new_n274), .C1(new_n262), .C2(new_n269), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n262), .A2(new_n269), .A3(new_n271), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT91), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n262), .A2(new_n269), .A3(new_n279), .A4(new_n271), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(KEYINPUT6), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n217), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(new_n280), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n216), .A2(KEYINPUT7), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n206), .B1(KEYINPUT93), .B2(new_n213), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n206), .A2(KEYINPUT93), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n207), .A2(KEYINPUT7), .A3(new_n216), .A4(new_n213), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n264), .B(new_n268), .Z(new_n290));
  XNOR2_X1  g104(.A(new_n271), .B(KEYINPUT92), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(KEYINPUT8), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n190), .B1(new_n282), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n217), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n278), .A2(KEYINPUT6), .A3(new_n280), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n265), .A2(new_n268), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n258), .A2(new_n259), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT85), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n258), .A2(KEYINPUT85), .A3(new_n259), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n300), .B1(new_n305), .B2(new_n248), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n274), .B1(new_n306), .B2(new_n271), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n270), .A2(KEYINPUT90), .A3(KEYINPUT6), .A4(new_n272), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n298), .B1(new_n299), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(G902), .B1(new_n283), .B2(new_n293), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n189), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n188), .B1(new_n297), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n315), .B(KEYINPUT80), .Z(new_n316));
  OR2_X1    g130(.A1(new_n316), .A2(G902), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G221), .ZN(new_n318));
  XOR2_X1   g132(.A(new_n318), .B(KEYINPUT81), .Z(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G469), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n211), .A2(new_n212), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n247), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n260), .B2(new_n261), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT11), .ZN(new_n325));
  INV_X1    g139(.A(G134), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(G137), .ZN(new_n327));
  INV_X1    g141(.A(G137), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(KEYINPUT11), .A3(G134), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(G137), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G131), .ZN(new_n332));
  INV_X1    g146(.A(G131), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n327), .A2(new_n329), .A3(new_n333), .A4(new_n330), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n263), .A2(G101), .ZN(new_n337));
  OAI22_X1  g151(.A1(new_n199), .A2(G128), .B1(new_n200), .B2(new_n194), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT86), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI221_X1 g154(.A(KEYINPUT86), .B1(new_n200), .B2(new_n194), .C1(new_n199), .C2(G128), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n201), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n258), .A2(new_n337), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n344));
  INV_X1    g158(.A(new_n202), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(new_n344), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n343), .A2(new_n344), .B1(new_n264), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n324), .A2(new_n336), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G110), .B(G140), .ZN(new_n349));
  INV_X1    g163(.A(G227), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(G953), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n349), .B(new_n351), .Z(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n336), .B1(new_n324), .B2(new_n347), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n258), .A2(new_n337), .A3(new_n342), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n202), .B1(new_n258), .B2(new_n337), .ZN(new_n357));
  OAI211_X1 g171(.A(KEYINPUT12), .B(new_n335), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n343), .B1(new_n202), .B2(new_n264), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT12), .B1(new_n360), .B2(new_n335), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n348), .B(KEYINPUT87), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n352), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n335), .B1(new_n356), .B2(new_n357), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT12), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n358), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT87), .B1(new_n368), .B2(new_n348), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n355), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n321), .B1(new_n370), .B2(new_n295), .ZN(new_n371));
  INV_X1    g185(.A(new_n348), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n363), .B1(new_n372), .B2(new_n354), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n368), .A2(new_n348), .A3(new_n352), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT88), .B(G469), .Z(new_n376));
  AND3_X1   g190(.A1(new_n375), .A2(new_n295), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n320), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT89), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(G902), .B1(new_n373), .B2(new_n374), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n376), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n348), .B1(new_n359), .B2(new_n361), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT87), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n362), .A3(new_n363), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n386), .B2(new_n355), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n382), .B1(new_n387), .B2(new_n321), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(KEYINPUT89), .A3(new_n320), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n314), .B1(new_n380), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G217), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(G234), .B2(new_n295), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G125), .B(G140), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n191), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G110), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n397), .A2(KEYINPUT24), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(KEYINPUT24), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT73), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT24), .B(G110), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT73), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT72), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(new_n220), .B2(G128), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT64), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G119), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n407), .A2(new_n409), .A3(new_n405), .A4(G128), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT71), .B1(new_n222), .B2(G128), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT71), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n196), .A3(G119), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n404), .B1(new_n406), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(KEYINPUT23), .B2(new_n196), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n196), .A2(KEYINPUT23), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n220), .B2(new_n419), .ZN(new_n420));
  XOR2_X1   g234(.A(KEYINPUT77), .B(G110), .Z(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n396), .B1(new_n423), .B2(KEYINPUT78), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n203), .A2(KEYINPUT75), .A3(G140), .A4(new_n204), .ZN(new_n425));
  AND2_X1   g239(.A1(KEYINPUT74), .A2(G125), .ZN(new_n426));
  NOR2_X1   g240(.A1(KEYINPUT74), .A2(G125), .ZN(new_n427));
  INV_X1    g241(.A(G140), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G125), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G140), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT75), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(KEYINPUT16), .B(new_n425), .C1(new_n429), .C2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT76), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI22_X1  g250(.A1(new_n205), .A2(new_n428), .B1(new_n432), .B2(new_n431), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n437), .A2(KEYINPUT76), .A3(KEYINPUT16), .A4(new_n425), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n205), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n440), .A2(KEYINPUT16), .A3(G140), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(G146), .A3(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n424), .B(new_n443), .C1(KEYINPUT78), .C2(new_n423), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n404), .A2(new_n415), .A3(new_n406), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n420), .A2(new_n397), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(G146), .B1(new_n439), .B2(new_n442), .ZN(new_n448));
  AOI211_X1 g262(.A(new_n191), .B(new_n441), .C1(new_n436), .C2(new_n438), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT22), .B(G137), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n454), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n444), .A2(new_n450), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(G902), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT25), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n393), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n444), .A2(new_n450), .A3(new_n456), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n456), .B1(new_n444), .B2(new_n450), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n295), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT25), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n455), .A2(new_n457), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n392), .A2(G902), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT79), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n326), .A2(G137), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n328), .A2(G134), .ZN(new_n473));
  OAI21_X1  g287(.A(G131), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n334), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n201), .B2(new_n198), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n332), .A2(new_n334), .B1(new_n211), .B2(new_n212), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT30), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n335), .A2(new_n322), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n334), .A2(new_n474), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n202), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT30), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n231), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT68), .ZN(new_n486));
  XOR2_X1   g300(.A(KEYINPUT66), .B(KEYINPUT27), .Z(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT67), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT26), .B(G101), .ZN(new_n489));
  NOR2_X1   g303(.A1(G237), .A2(G953), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G210), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n489), .B(new_n491), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n488), .B(new_n492), .Z(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n229), .A2(new_n230), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n479), .A3(new_n481), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n485), .A2(new_n486), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT31), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n495), .B1(new_n478), .B2(new_n483), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n231), .A2(new_n476), .A3(new_n477), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n499), .A2(new_n493), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT31), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n486), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT28), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n231), .B1(new_n476), .B2(new_n477), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(new_n496), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n500), .A2(KEYINPUT28), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n493), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n498), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G472), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n509), .A2(KEYINPUT32), .A3(new_n510), .A4(new_n295), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n511), .A2(new_n512), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n508), .B1(new_n497), .B2(KEYINPUT31), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n502), .B1(new_n501), .B2(new_n486), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n510), .B(new_n295), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT32), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n513), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n506), .A2(new_n507), .A3(new_n493), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(KEYINPUT29), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n499), .A2(new_n500), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(new_n494), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT69), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT69), .B1(new_n523), .B2(new_n494), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(G902), .B1(new_n521), .B2(KEYINPUT29), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n510), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n471), .B1(new_n520), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n439), .A2(new_n442), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n191), .ZN(new_n534));
  AOI21_X1  g348(.A(G143), .B1(new_n490), .B2(G214), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n490), .A2(G143), .A3(G214), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT94), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n490), .A2(KEYINPUT94), .A3(G143), .A4(G214), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n540), .A2(new_n541), .A3(new_n333), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n539), .ZN(new_n543));
  INV_X1    g357(.A(new_n535), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n333), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI211_X1 g359(.A(G131), .B(new_n535), .C1(new_n538), .C2(new_n539), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n542), .B1(new_n547), .B2(new_n541), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n534), .A2(new_n443), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(G113), .B(G122), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(new_n235), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n437), .A2(new_n425), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G146), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n554), .A3(new_n395), .ZN(new_n555));
  AND2_X1   g369(.A1(KEYINPUT18), .A2(G131), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n540), .B(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n191), .B1(new_n437), .B2(new_n425), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT95), .B1(new_n558), .B2(new_n396), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n549), .A2(new_n551), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n552), .A2(KEYINPUT19), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT19), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n394), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT96), .B1(new_n394), .B2(new_n563), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n562), .A2(new_n191), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n545), .B2(new_n546), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n560), .B1(new_n570), .B2(new_n449), .ZN(new_n571));
  INV_X1    g385(.A(new_n551), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n561), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT97), .ZN(new_n575));
  NOR2_X1   g389(.A1(G475), .A2(G902), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n561), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n576), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT20), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n579), .A2(KEYINPUT20), .B1(new_n574), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n549), .A2(new_n560), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n572), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n561), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n295), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G475), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n225), .A2(G122), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n225), .A2(G122), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n589), .B1(new_n590), .B2(KEYINPUT14), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(KEYINPUT14), .B2(new_n589), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n592), .A2(KEYINPUT98), .A3(G107), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT98), .B1(new_n592), .B2(G107), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G122), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G116), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n597), .A2(new_n589), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n254), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n193), .A2(G128), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n193), .A2(G128), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n326), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n326), .B1(new_n601), .B2(new_n602), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n599), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n595), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n598), .B(new_n254), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT13), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n602), .B1(new_n600), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n609), .B2(new_n602), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G134), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n608), .A2(new_n612), .A3(new_n603), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n316), .A2(new_n391), .A3(G953), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n607), .A2(new_n613), .A3(new_n615), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n295), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT15), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n621), .A2(KEYINPUT15), .ZN(new_n624));
  OAI21_X1  g438(.A(G478), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n620), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(G234), .A2(G237), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n628), .A2(G952), .A3(new_n215), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n628), .A2(G902), .A3(G953), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT21), .B(G898), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR4_X1   g446(.A1(new_n582), .A2(new_n588), .A3(new_n627), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n390), .A2(new_n532), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G101), .ZN(G3));
  OAI21_X1  g449(.A(new_n295), .B1(new_n515), .B2(new_n516), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n510), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n509), .B(new_n295), .C1(new_n637), .C2(new_n510), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI211_X1 g455(.A(new_n470), .B(new_n641), .C1(new_n380), .C2(new_n389), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n574), .A2(new_n581), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n561), .A2(new_n573), .A3(new_n577), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n577), .B1(new_n561), .B2(new_n573), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n644), .A2(new_n645), .A3(new_n580), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT20), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n587), .ZN(new_n649));
  AOI211_X1 g463(.A(G478), .B(G902), .C1(new_n617), .C2(new_n618), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n614), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT33), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n619), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n652), .A2(new_n617), .A3(KEYINPUT33), .A4(new_n618), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n295), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n650), .B1(new_n656), .B2(G478), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n649), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n632), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n313), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n642), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  NAND2_X1  g479(.A1(new_n575), .A2(new_n578), .ZN(new_n666));
  INV_X1    g480(.A(new_n581), .ZN(new_n667));
  OAI22_X1  g481(.A1(new_n646), .A2(new_n647), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n627), .A2(new_n587), .ZN(new_n670));
  NOR4_X1   g484(.A1(new_n314), .A2(new_n632), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n642), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  NOR2_X1   g488(.A1(new_n456), .A2(KEYINPUT36), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n451), .B(new_n675), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n460), .A2(new_n464), .B1(new_n468), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n641), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n390), .A2(new_n633), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT37), .B(G110), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  NAND3_X1  g495(.A1(new_n519), .A2(new_n512), .A3(new_n511), .ZN(new_n682));
  INV_X1    g496(.A(new_n636), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n510), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n530), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n630), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n629), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n668), .A2(new_n587), .A3(new_n627), .A4(new_n689), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n685), .A2(new_n690), .A3(new_n677), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n390), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  AND2_X1   g507(.A1(new_n649), .A2(new_n627), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n682), .A2(new_n684), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n494), .B1(new_n496), .B2(new_n505), .ZN(new_n696));
  OR3_X1    g510(.A1(new_n696), .A2(new_n501), .A3(KEYINPUT102), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT102), .B1(new_n696), .B2(new_n501), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n295), .A3(new_n698), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n699), .A2(KEYINPUT103), .A3(G472), .ZN(new_n700));
  AOI21_X1  g514(.A(KEYINPUT103), .B1(new_n699), .B2(G472), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n695), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n694), .A2(new_n703), .A3(new_n187), .A4(new_n677), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n297), .A2(new_n312), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n705), .B(KEYINPUT38), .Z(new_n706));
  NAND2_X1  g520(.A1(new_n380), .A2(new_n389), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n689), .B(KEYINPUT39), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI211_X1 g523(.A(new_n704), .B(new_n706), .C1(KEYINPUT40), .C2(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  OAI211_X1 g527(.A(new_n657), .B(new_n689), .C1(new_n582), .C2(new_n588), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n685), .A2(new_n714), .A3(new_n677), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n390), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  NOR2_X1   g531(.A1(new_n381), .A2(new_n321), .ZN(new_n718));
  INV_X1    g532(.A(new_n318), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n377), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n661), .A2(new_n531), .A3(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT41), .B(G113), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NOR2_X1   g538(.A1(new_n531), .A2(new_n721), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n671), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  INV_X1    g541(.A(new_n685), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n676), .A2(new_n468), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n392), .B1(new_n463), .B2(KEYINPUT25), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n459), .B1(new_n466), .B2(new_n295), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n633), .A2(new_n313), .A3(new_n720), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n222), .ZN(G21));
  NAND2_X1  g550(.A1(new_n694), .A2(new_n313), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n636), .A2(G472), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n738), .A2(new_n517), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n720), .A2(new_n471), .A3(new_n660), .A4(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n596), .ZN(G24));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n738), .A2(new_n517), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n677), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(new_n649), .A3(new_n657), .A4(new_n689), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n313), .A2(new_n720), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n739), .A2(new_n732), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n714), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(KEYINPUT104), .A3(new_n313), .A4(new_n720), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  NAND3_X1  g567(.A1(new_n297), .A2(new_n312), .A3(new_n187), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n297), .A2(new_n312), .A3(KEYINPUT106), .A4(new_n187), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n318), .B1(new_n371), .B2(new_n377), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(KEYINPUT105), .B(new_n318), .C1(new_n371), .C2(new_n377), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n511), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n530), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n470), .B1(new_n766), .B2(new_n519), .ZN(new_n767));
  INV_X1    g581(.A(new_n714), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n768), .A3(KEYINPUT42), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n758), .A2(new_n532), .A3(new_n768), .A4(new_n763), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT42), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n772), .B2(new_n773), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n771), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G131), .ZN(G33));
  INV_X1    g592(.A(new_n690), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n758), .A2(new_n532), .A3(new_n779), .A4(new_n763), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n355), .B(new_n782), .C1(new_n364), .C2(new_n369), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n782), .B1(new_n386), .B2(new_n355), .ZN(new_n785));
  OAI21_X1  g599(.A(G469), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(G469), .A2(G902), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(KEYINPUT46), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n370), .A2(KEYINPUT45), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n783), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n789), .B(G469), .C1(new_n791), .C2(G902), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n788), .A2(new_n792), .A3(new_n382), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n793), .A2(new_n318), .A3(new_n708), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n648), .A2(new_n587), .A3(new_n657), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT43), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n732), .A2(new_n641), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT108), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT43), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n648), .A2(new_n587), .A3(new_n657), .A4(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT108), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n732), .A2(new_n641), .A3(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n796), .A2(new_n798), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT44), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n732), .A2(new_n641), .A3(new_n801), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n801), .B1(new_n732), .B2(new_n641), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n808), .A3(new_n796), .A4(new_n800), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n794), .A2(new_n810), .A3(new_n758), .ZN(new_n811));
  XOR2_X1   g625(.A(KEYINPUT109), .B(G137), .Z(new_n812));
  XNOR2_X1  g626(.A(new_n811), .B(new_n812), .ZN(G39));
  NAND2_X1  g627(.A1(new_n793), .A2(new_n318), .ZN(new_n814));
  XOR2_X1   g628(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n815), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n793), .A2(new_n318), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n756), .A2(new_n757), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n819), .A2(new_n471), .A3(new_n728), .A4(new_n714), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G140), .ZN(G42));
  NAND3_X1  g636(.A1(new_n471), .A2(new_n320), .A3(new_n187), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT111), .Z(new_n824));
  NOR2_X1   g638(.A1(new_n377), .A2(new_n718), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n795), .B1(new_n826), .B2(KEYINPUT49), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT112), .Z(new_n829));
  INV_X1    g643(.A(new_n703), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n826), .A2(KEYINPUT49), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n829), .A2(new_n706), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT113), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n819), .A2(new_n688), .A3(new_n721), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n471), .A3(new_n830), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n835), .A2(KEYINPUT117), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(KEYINPUT117), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n659), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n796), .A2(new_n800), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n470), .A2(new_n688), .A3(new_n744), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n747), .ZN(new_n842));
  INV_X1    g656(.A(G952), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n842), .A2(new_n843), .A3(G953), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n838), .A2(KEYINPUT118), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT118), .B1(new_n838), .B2(new_n844), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n834), .A2(new_n839), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n767), .ZN(new_n848));
  NOR2_X1   g662(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n847), .B(new_n767), .C1(KEYINPUT119), .C2(KEYINPUT48), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n850), .A2(new_n851), .B1(KEYINPUT119), .B2(KEYINPUT48), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n845), .A2(new_n846), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n649), .A2(new_n657), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n836), .A2(new_n837), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n721), .A2(new_n187), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n706), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT50), .ZN(new_n858));
  OR3_X1    g672(.A1(new_n857), .A2(new_n858), .A3(new_n841), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n858), .B1(new_n857), .B2(new_n841), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n859), .A2(new_n860), .B1(new_n745), .B2(new_n847), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n855), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n855), .A2(new_n861), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n816), .A2(new_n818), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n825), .A2(new_n319), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n819), .B(new_n841), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n863), .B(new_n864), .C1(new_n866), .C2(new_n869), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n853), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n707), .B(new_n313), .C1(new_n691), .C2(new_n715), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n729), .B(new_n689), .C1(new_n730), .C2(new_n731), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT115), .B1(new_n759), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n877));
  INV_X1    g691(.A(new_n875), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n388), .A2(new_n877), .A3(new_n878), .A4(new_n318), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n694), .A2(new_n313), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n881), .A3(new_n703), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n752), .A2(new_n874), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT52), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n752), .A2(new_n874), .A3(new_n882), .A4(KEYINPUT52), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n648), .A2(new_n587), .A3(new_n627), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n658), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n889), .A2(new_n632), .A3(new_n314), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n890), .A2(new_n642), .B1(new_n671), .B2(new_n725), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n733), .A2(new_n734), .B1(new_n737), .B2(new_n740), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n722), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n390), .B(new_n633), .C1(new_n532), .C2(new_n678), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n758), .A2(new_n750), .A3(new_n763), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n780), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n627), .B1(new_n688), .B2(new_n687), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(new_n587), .A3(new_n668), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n707), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n728), .A2(new_n756), .A3(new_n732), .A4(new_n757), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT114), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n902), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT114), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n899), .B1(new_n380), .B2(new_n389), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n897), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n887), .A2(new_n777), .A3(new_n895), .A4(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n907), .A2(new_n903), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n913), .A3(new_n897), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(KEYINPUT53), .A3(new_n777), .A4(new_n887), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n911), .A2(new_n915), .A3(KEYINPUT54), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n873), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(G952), .A2(G953), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n833), .B1(new_n920), .B2(new_n921), .ZN(G75));
  NAND3_X1  g736(.A1(new_n916), .A2(G210), .A3(G902), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT56), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n299), .A2(new_n309), .A3(new_n298), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n282), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n928), .B1(new_n923), .B2(new_n924), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n215), .A2(G952), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(G51));
  XOR2_X1   g747(.A(new_n787), .B(KEYINPUT57), .Z(new_n934));
  NAND3_X1  g748(.A1(new_n918), .A2(new_n919), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n375), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n916), .A2(G469), .A3(G902), .A4(new_n791), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(G54));
  INV_X1    g752(.A(new_n932), .ZN(new_n939));
  NAND2_X1  g753(.A1(KEYINPUT58), .A2(G475), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n295), .B(new_n940), .C1(new_n911), .C2(new_n915), .ZN(new_n941));
  INV_X1    g755(.A(new_n666), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n944), .A2(new_n666), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT120), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n932), .B1(new_n944), .B2(new_n666), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT120), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n941), .A2(new_n942), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n950), .ZN(G60));
  NAND2_X1  g765(.A1(G478), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT59), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n918), .A2(new_n919), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n654), .A2(new_n655), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n939), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n954), .A2(new_n955), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(G63));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT60), .Z(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n911), .B2(new_n915), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n963), .A2(new_n466), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n932), .B1(new_n963), .B2(new_n676), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT121), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(new_n963), .B2(new_n676), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n964), .B(new_n965), .C1(new_n968), .C2(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(G66));
  NAND2_X1  g786(.A1(G224), .A2(G953), .ZN(new_n973));
  OAI22_X1  g787(.A1(new_n912), .A2(G953), .B1(new_n631), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT122), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n276), .B(new_n281), .C1(G898), .C2(new_n215), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  NAND2_X1  g791(.A1(new_n562), .A2(new_n568), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n484), .B(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT125), .ZN(new_n981));
  INV_X1    g795(.A(new_n762), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT105), .B1(new_n388), .B2(new_n318), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR4_X1   g798(.A1(new_n984), .A2(new_n819), .A3(new_n531), .A4(new_n714), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT42), .B1(new_n985), .B2(KEYINPUT107), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n772), .A2(new_n773), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n770), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n780), .A2(new_n752), .A3(new_n874), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n694), .A2(new_n767), .A3(new_n313), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n990), .A2(new_n318), .A3(new_n793), .A4(new_n708), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n989), .A2(new_n811), .A3(new_n821), .A4(new_n991), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n988), .A2(new_n992), .A3(KEYINPUT124), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT124), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n821), .A2(new_n811), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n991), .A2(new_n780), .A3(new_n752), .A4(new_n874), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n994), .B1(new_n997), .B2(new_n777), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n215), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n215), .A2(G900), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n981), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(KEYINPUT124), .B1(new_n988), .B2(new_n992), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n821), .A2(new_n811), .ZN(new_n1004));
  INV_X1    g818(.A(new_n996), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n777), .A2(new_n1004), .A3(new_n994), .A4(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(G953), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n1007), .A2(KEYINPUT125), .A3(new_n1000), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n980), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n889), .B(KEYINPUT123), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n1010), .A2(new_n531), .A3(new_n819), .ZN(new_n1011));
  INV_X1    g825(.A(new_n709), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n995), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n752), .A2(new_n874), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n712), .A2(KEYINPUT62), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(KEYINPUT62), .B1(new_n712), .B2(new_n1014), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n980), .B1(new_n1017), .B2(new_n215), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(G953), .B1(new_n350), .B2(new_n686), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT126), .Z(new_n1021));
  NAND3_X1  g835(.A1(new_n1009), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1021), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n999), .A2(new_n981), .A3(new_n1001), .ZN(new_n1024));
  OAI21_X1  g838(.A(KEYINPUT125), .B1(new_n1007), .B2(new_n1000), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n979), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1023), .B1(new_n1026), .B2(new_n1018), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1022), .A2(new_n1027), .ZN(G72));
  NAND2_X1  g842(.A1(G472), .A2(G902), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT63), .Z(new_n1030));
  OAI21_X1  g844(.A(new_n1030), .B1(new_n1017), .B2(new_n912), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n523), .A2(new_n493), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n932), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1003), .A2(new_n895), .A3(new_n1006), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(new_n1030), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1035), .A2(new_n493), .A3(new_n523), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n526), .A2(new_n527), .ZN(new_n1037));
  OAI211_X1 g851(.A(new_n916), .B(new_n1030), .C1(new_n1037), .C2(new_n501), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1033), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(KEYINPUT127), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT127), .ZN(new_n1041));
  NAND4_X1  g855(.A1(new_n1033), .A2(new_n1036), .A3(new_n1038), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1040), .A2(new_n1042), .ZN(G57));
endmodule


