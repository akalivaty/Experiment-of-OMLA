//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1226, new_n1227, new_n1228, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n207), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n210), .B(new_n216), .C1(new_n223), .C2(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(G226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT67), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G68), .Z(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(new_n213), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(KEYINPUT8), .B(G58), .Z(new_n247));
  NAND2_X1  g0047(.A1(new_n214), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n247), .A2(new_n249), .B1(G150), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n204), .A2(G20), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n246), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT68), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(new_n214), .B2(G1), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(KEYINPUT68), .A3(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G50), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n246), .A2(new_n260), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n259), .A2(new_n261), .B1(G50), .B2(new_n260), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT9), .ZN(new_n263));
  OR3_X1    g0063(.A1(new_n253), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G200), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n270), .A3(G274), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n268), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(G226), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G222), .A2(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G223), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n280), .B(new_n273), .C1(G77), .C2(new_n276), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n265), .B1(new_n275), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n263), .B1(new_n253), .B2(new_n262), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n275), .A2(G190), .A3(new_n281), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n264), .A2(new_n283), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT10), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n275), .A2(new_n281), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n282), .B1(new_n289), .B2(G190), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT10), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(new_n264), .A4(new_n284), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n253), .A2(new_n262), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n295), .B(new_n296), .C1(G179), .C2(new_n288), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n276), .A2(G238), .A3(G1698), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n276), .A2(G232), .A3(new_n278), .ZN(new_n301));
  INV_X1    g0101(.A(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT3), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT3), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G107), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n300), .A2(new_n301), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n273), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n272), .B1(G244), .B2(new_n274), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT69), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT69), .B1(new_n309), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n299), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n309), .A2(new_n310), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT69), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n317), .A2(new_n294), .A3(new_n311), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n247), .A2(new_n250), .B1(G20), .B2(G77), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT15), .B(G87), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n249), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n245), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n258), .A2(G77), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n325), .A2(new_n261), .B1(G77), .B2(new_n260), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n314), .A2(new_n318), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n298), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(G190), .B1(new_n312), .B2(new_n313), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n317), .A2(G200), .A3(new_n311), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT70), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n324), .B2(new_n327), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n246), .B1(new_n319), .B2(new_n322), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n336), .A2(new_n326), .A3(KEYINPUT70), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n332), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n260), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n203), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n342), .A2(KEYINPUT12), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(KEYINPUT12), .ZN(new_n344));
  INV_X1    g0144(.A(new_n258), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n203), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n341), .A2(new_n245), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n343), .A2(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n250), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n349));
  INV_X1    g0149(.A(G77), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n248), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n245), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT11), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(KEYINPUT11), .A3(new_n245), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n348), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT73), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n348), .A2(new_n354), .A3(KEYINPUT73), .A4(new_n355), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT14), .ZN(new_n362));
  INV_X1    g0162(.A(G226), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n278), .ZN(new_n364));
  INV_X1    g0164(.A(G232), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G1698), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n303), .A2(new_n364), .A3(new_n305), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G97), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT71), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT71), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(new_n371), .A3(new_n368), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n372), .A3(new_n273), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n270), .A2(G238), .A3(new_n374), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n271), .A2(new_n375), .A3(KEYINPUT72), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT72), .B1(new_n271), .B2(new_n375), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT13), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n373), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n379), .B1(new_n373), .B2(new_n378), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n362), .B(G169), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n373), .A2(new_n378), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT13), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n373), .A2(new_n378), .A3(new_n379), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(G179), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n385), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n362), .B1(new_n388), .B2(G169), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n361), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(G200), .B1(new_n380), .B2(new_n381), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n384), .A2(G190), .A3(new_n385), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n360), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n247), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(new_n345), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(new_n347), .B1(new_n341), .B2(new_n395), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(G58), .B(G68), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G20), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n250), .A2(G159), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n304), .A2(G33), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n302), .A2(KEYINPUT3), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n214), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n203), .B1(new_n405), .B2(KEYINPUT7), .ZN(new_n406));
  AOI21_X1  g0206(.A(G20), .B1(new_n303), .B2(new_n305), .ZN(new_n407));
  AND2_X1   g0207(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n408));
  NOR2_X1   g0208(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n402), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n246), .B1(new_n412), .B2(KEYINPUT16), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT75), .B1(new_n304), .B2(G33), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT75), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(new_n302), .A3(KEYINPUT3), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n417), .A3(new_n305), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT7), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(G20), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n410), .B1(new_n276), .B2(G20), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n203), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n414), .B1(new_n423), .B2(new_n402), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n398), .B1(new_n413), .B2(new_n424), .ZN(new_n425));
  OR2_X1    g0225(.A1(G223), .A2(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n363), .A2(G1698), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n303), .A2(new_n426), .A3(new_n305), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G87), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n273), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n270), .A2(G232), .A3(new_n374), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n271), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n294), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n270), .B1(new_n428), .B2(new_n429), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n271), .A2(new_n432), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n435), .A2(new_n436), .A3(new_n299), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT18), .B1(new_n425), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n421), .A2(new_n422), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G68), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n399), .A2(G20), .B1(G159), .B2(new_n250), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT16), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(G68), .B1(new_n407), .B2(new_n419), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n306), .A2(new_n410), .A3(new_n214), .ZN(new_n445));
  OAI211_X1 g0245(.A(KEYINPUT16), .B(new_n442), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n245), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n397), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT18), .ZN(new_n449));
  INV_X1    g0249(.A(new_n438), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n265), .B1(new_n431), .B2(new_n433), .ZN(new_n453));
  INV_X1    g0253(.A(G190), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n435), .A2(new_n436), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n452), .B1(new_n425), .B2(new_n456), .ZN(new_n457));
  XOR2_X1   g0257(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n424), .A2(new_n245), .A3(new_n446), .ZN(new_n460));
  AND4_X1   g0260(.A1(new_n459), .A2(new_n460), .A3(new_n397), .A4(new_n456), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n439), .B(new_n451), .C1(new_n457), .C2(new_n461), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n340), .A2(new_n394), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n303), .A2(new_n305), .A3(G244), .A4(G1698), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n303), .A2(new_n305), .A3(G238), .A4(new_n278), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G116), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n273), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n267), .A2(G1), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n270), .A2(G274), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n256), .A2(G45), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n270), .A2(G250), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n468), .A2(new_n299), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n473), .B1(new_n273), .B2(new_n467), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(G169), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n321), .A2(new_n260), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n256), .A2(G33), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n246), .A2(new_n260), .A3(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n303), .A2(new_n305), .A3(new_n214), .A4(G68), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT19), .ZN(new_n484));
  INV_X1    g0284(.A(G97), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n484), .B1(new_n248), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n214), .B1(new_n368), .B2(new_n484), .ZN(new_n488));
  INV_X1    g0288(.A(G87), .ZN(new_n489));
  INV_X1    g0289(.A(G107), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT78), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n488), .A2(KEYINPUT78), .A3(new_n491), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI221_X1 g0295(.A(new_n480), .B1(new_n320), .B2(new_n482), .C1(new_n495), .C2(new_n246), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n468), .A2(G190), .A3(new_n474), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n265), .B1(new_n468), .B2(new_n474), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n482), .A2(new_n489), .ZN(new_n500));
  INV_X1    g0300(.A(new_n494), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n483), .B(new_n486), .C1(new_n501), .C2(new_n492), .ZN(new_n502));
  AOI211_X1 g0302(.A(new_n479), .B(new_n500), .C1(new_n502), .C2(new_n245), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n478), .A2(new_n496), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n303), .A2(new_n305), .A3(G244), .A4(new_n278), .ZN(new_n505));
  NOR2_X1   g0305(.A1(KEYINPUT77), .A2(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n506), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n276), .A2(G244), .A3(new_n278), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n507), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n273), .ZN(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT5), .B(G41), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n514), .A2(G274), .A3(new_n270), .A4(new_n469), .ZN(new_n515));
  NAND2_X1  g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(KEYINPUT5), .A2(G41), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n469), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n270), .ZN(new_n520));
  INV_X1    g0320(.A(G257), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n513), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n294), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n490), .B1(new_n421), .B2(new_n422), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n250), .A2(G77), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT6), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n528), .A2(new_n485), .A3(G107), .ZN(new_n529));
  XNOR2_X1  g0329(.A(G97), .B(G107), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n529), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n527), .B1(new_n531), .B2(new_n214), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n245), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n260), .A2(G97), .ZN(new_n534));
  INV_X1    g0334(.A(new_n482), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n534), .B1(new_n535), .B2(G97), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n522), .B1(new_n512), .B2(new_n273), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n299), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n525), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n533), .A2(new_n536), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n524), .A2(G190), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n538), .A2(G200), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n504), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n303), .A2(new_n305), .A3(new_n214), .A4(G87), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT22), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT22), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n276), .A2(new_n548), .A3(new_n214), .A4(G87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT24), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n466), .A2(G20), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT23), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n214), .B2(G107), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n490), .A2(KEYINPUT23), .A3(G20), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n550), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n551), .B1(new_n550), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n245), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n260), .A2(G107), .ZN(new_n560));
  XNOR2_X1  g0360(.A(KEYINPUT80), .B(KEYINPUT25), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n560), .B(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(G107), .B2(new_n535), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n303), .A2(new_n305), .A3(G257), .A4(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n303), .A2(new_n305), .A3(G250), .A4(new_n278), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G294), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n273), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n273), .B1(new_n469), .B2(new_n514), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G264), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n571), .A3(new_n515), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n294), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n568), .A2(new_n273), .B1(new_n570), .B2(G264), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(new_n299), .A3(new_n515), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n564), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(G190), .A3(new_n515), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n572), .A2(G200), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n559), .A2(new_n563), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n519), .A2(G270), .A3(new_n270), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n581), .A2(new_n515), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n303), .A2(new_n305), .A3(G264), .A4(G1698), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n303), .A2(new_n305), .A3(G257), .A4(new_n278), .ZN(new_n584));
  XOR2_X1   g0384(.A(KEYINPUT79), .B(G303), .Z(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n276), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n273), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n347), .A2(G116), .A3(new_n481), .ZN(new_n589));
  INV_X1    g0389(.A(G116), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n341), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n244), .A2(new_n213), .B1(G20), .B2(new_n590), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n510), .B(new_n214), .C1(G33), .C2(new_n485), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n592), .A2(KEYINPUT20), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT20), .B1(new_n592), .B2(new_n593), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n589), .B(new_n591), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n588), .A2(KEYINPUT21), .A3(new_n596), .A4(G169), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n581), .A2(new_n515), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n273), .B2(new_n586), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(G179), .A3(new_n596), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n588), .A2(G169), .A3(new_n596), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n596), .B1(new_n588), .B2(G200), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n454), .B2(new_n588), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n601), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n545), .A2(new_n580), .A3(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n463), .A2(new_n608), .ZN(G372));
  NOR2_X1   g0409(.A1(new_n457), .A2(new_n461), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n330), .A2(new_n393), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n610), .B1(new_n390), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT82), .ZN(new_n613));
  AOI211_X1 g0413(.A(KEYINPUT18), .B(new_n438), .C1(new_n460), .C2(new_n397), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n449), .B1(new_n448), .B2(new_n450), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n439), .A2(KEYINPUT82), .A3(new_n451), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n293), .B1(new_n612), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT83), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n620), .A2(new_n621), .A3(new_n297), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n620), .B2(new_n297), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n478), .A2(new_n496), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n504), .A2(new_n544), .A3(new_n540), .A4(new_n579), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n573), .A2(new_n575), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n559), .B2(new_n563), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n604), .A2(new_n600), .A3(new_n597), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n625), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n525), .A2(new_n537), .A3(new_n539), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT26), .B1(new_n504), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n482), .A2(new_n320), .ZN(new_n634));
  AOI211_X1 g0434(.A(new_n479), .B(new_n634), .C1(new_n502), .C2(new_n245), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n468), .A2(G190), .A3(new_n474), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n265), .B2(new_n476), .ZN(new_n637));
  INV_X1    g0437(.A(new_n500), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n638), .B(new_n480), .C1(new_n495), .C2(new_n246), .ZN(new_n639));
  OAI22_X1  g0439(.A1(new_n635), .A2(new_n477), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  XOR2_X1   g0440(.A(KEYINPUT81), .B(KEYINPUT26), .Z(new_n641));
  NOR3_X1   g0441(.A1(new_n640), .A2(new_n540), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n633), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n463), .B1(new_n631), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n624), .A2(new_n644), .ZN(G369));
  NAND3_X1  g0445(.A1(new_n256), .A2(new_n214), .A3(G13), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(G343), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n596), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n629), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n607), .B2(new_n652), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G330), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n651), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n559), .B2(new_n563), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n580), .A2(new_n659), .B1(new_n576), .B2(new_n658), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n579), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n628), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n651), .B1(new_n601), .B2(new_n604), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n576), .B2(new_n651), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n661), .A2(new_n666), .ZN(G399));
  INV_X1    g0467(.A(new_n208), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n491), .A2(G116), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G1), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n211), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  AOI21_X1  g0474(.A(G179), .B1(new_n582), .B2(new_n587), .ZN(new_n675));
  INV_X1    g0475(.A(new_n476), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n524), .A2(new_n675), .A3(new_n676), .A4(new_n572), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT84), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n599), .A2(G179), .A3(new_n476), .A4(new_n574), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n524), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n513), .A2(new_n523), .B1(new_n574), .B2(new_n515), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT84), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n676), .A4(new_n675), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n588), .A2(new_n299), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n574), .A2(new_n476), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT30), .A4(new_n538), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n678), .A2(new_n681), .A3(new_n684), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n651), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT31), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT85), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT85), .ZN(new_n692));
  AOI211_X1 g0492(.A(new_n692), .B(KEYINPUT31), .C1(new_n688), .C2(new_n651), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n651), .A2(KEYINPUT31), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n681), .A2(new_n687), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n677), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n608), .B2(new_n658), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n656), .B1(new_n694), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n658), .B1(new_n631), .B2(new_n643), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n504), .A2(new_n632), .ZN(new_n703));
  INV_X1    g0503(.A(new_n641), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(KEYINPUT26), .B2(new_n703), .ZN(new_n706));
  OAI211_X1 g0506(.A(KEYINPUT29), .B(new_n658), .C1(new_n706), .C2(new_n631), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n699), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n674), .B1(new_n708), .B2(G1), .ZN(G364));
  AND2_X1   g0509(.A1(new_n214), .A2(G13), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n256), .B1(new_n710), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n669), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n657), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(G330), .B2(new_n654), .ZN(new_n715));
  INV_X1    g0515(.A(new_n713), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n213), .B1(G20), .B2(new_n294), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n299), .A2(new_n265), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT90), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n214), .A2(G190), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G159), .ZN(new_n724));
  XOR2_X1   g0524(.A(KEYINPUT91), .B(KEYINPUT32), .Z(new_n725));
  XNOR2_X1  g0525(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(G20), .B1(new_n720), .B2(new_n454), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n485), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n214), .A2(new_n454), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n299), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT89), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n733), .A2(new_n734), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G58), .ZN(new_n740));
  NAND3_X1  g0540(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G190), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n741), .A2(new_n454), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n743), .A2(new_n203), .B1(new_n745), .B2(new_n201), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n732), .A2(new_n721), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n265), .A2(G179), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n721), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n747), .A2(new_n350), .B1(new_n749), .B2(new_n490), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n731), .A2(new_n748), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n276), .B1(new_n751), .B2(new_n489), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n746), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n726), .A2(new_n730), .A3(new_n740), .A4(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n751), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n276), .B1(new_n755), .B2(G303), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT92), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n739), .B2(G322), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n723), .A2(G329), .B1(new_n756), .B2(new_n757), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n727), .A2(G294), .ZN(new_n761));
  INV_X1    g0561(.A(G326), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n745), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  INV_X1    g0564(.A(G283), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n747), .A2(new_n764), .B1(new_n749), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT33), .B(G317), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n763), .B(new_n766), .C1(new_n742), .C2(new_n767), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n759), .A2(new_n760), .A3(new_n761), .A4(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n718), .B1(new_n754), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n717), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n668), .A2(new_n306), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT86), .ZN(new_n776));
  XOR2_X1   g0576(.A(G355), .B(KEYINPUT87), .Z(new_n777));
  AOI22_X1  g0577(.A1(new_n776), .A2(new_n777), .B1(new_n590), .B2(new_n668), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n668), .A2(new_n276), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n212), .B2(new_n267), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT88), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n267), .B2(new_n242), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n781), .A2(new_n782), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n778), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n716), .B(new_n770), .C1(new_n774), .C2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n773), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n654), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n715), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G396));
  NAND2_X1  g0591(.A1(new_n328), .A2(new_n651), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n339), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n329), .ZN(new_n794));
  AND4_X1   g0594(.A1(new_n328), .A2(new_n314), .A3(new_n318), .A4(new_n658), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n700), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n795), .B1(new_n329), .B2(new_n793), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n658), .B(new_n799), .C1(new_n631), .C2(new_n643), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n699), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n670), .B2(new_n711), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n699), .A2(new_n798), .A3(new_n800), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n718), .A2(new_n772), .ZN(new_n805));
  INV_X1    g0605(.A(new_n747), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n806), .A2(G159), .B1(G137), .B2(new_n744), .ZN(new_n807));
  INV_X1    g0607(.A(G150), .ZN(new_n808));
  INV_X1    g0608(.A(G143), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n808), .B2(new_n743), .C1(new_n738), .C2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT34), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n751), .A2(new_n201), .B1(new_n749), .B2(new_n203), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT94), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n306), .B1(new_n723), .B2(G132), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n202), .C2(new_n728), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n749), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n723), .A2(G311), .B1(G87), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT93), .ZN(new_n819));
  INV_X1    g0619(.A(G294), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n738), .A2(new_n820), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n306), .B1(new_n747), .B2(new_n590), .C1(new_n490), .C2(new_n751), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n744), .A2(G303), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n743), .B2(new_n765), .ZN(new_n824));
  NOR4_X1   g0624(.A1(new_n729), .A2(new_n821), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n811), .A2(new_n816), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n713), .B1(G77), .B2(new_n805), .C1(new_n826), .C2(new_n718), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n771), .B2(new_n797), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT95), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n804), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G384));
  NAND2_X1  g0631(.A1(new_n530), .A2(new_n528), .ZN(new_n832));
  INV_X1    g0632(.A(new_n529), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n834), .A2(KEYINPUT35), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(KEYINPUT35), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n835), .A2(G116), .A3(new_n215), .A4(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(KEYINPUT96), .B(KEYINPUT36), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n837), .B(new_n838), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n350), .B(new_n211), .C1(G58), .C2(G68), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT97), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n840), .A2(new_n841), .B1(new_n201), .B2(G68), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n256), .B(G13), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(G169), .B1(new_n380), .B2(new_n381), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT14), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(new_n386), .A3(new_n382), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(new_n361), .A3(new_n658), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT99), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  INV_X1    g0652(.A(new_n649), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n448), .A2(new_n853), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n457), .A2(new_n461), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n854), .B1(new_n618), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n448), .A2(new_n450), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n460), .A2(new_n397), .A3(new_n456), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n857), .A2(new_n854), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n852), .B1(new_n856), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT98), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT98), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n868), .B(new_n442), .C1(new_n444), .C2(new_n445), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n414), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n398), .B1(new_n870), .B2(new_n413), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n858), .B1(new_n871), .B2(new_n649), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n871), .A2(new_n438), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT37), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n871), .A2(new_n649), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n874), .A2(new_n862), .B1(new_n462), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT39), .B1(new_n876), .B2(KEYINPUT38), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n865), .A2(new_n877), .A3(KEYINPUT100), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n874), .A2(new_n862), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n462), .A2(new_n875), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n879), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT39), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT100), .B1(new_n865), .B2(new_n877), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n851), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n618), .A2(new_n853), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n800), .A2(new_n796), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n361), .A2(new_n651), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n390), .A2(new_n393), .A3(new_n890), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n360), .A2(new_n391), .A3(new_n392), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n361), .B(new_n651), .C1(new_n848), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n881), .A2(new_n882), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n888), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n886), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT101), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n886), .A2(KEYINPUT101), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n463), .A2(new_n702), .A3(new_n707), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n624), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n903), .B(new_n905), .Z(new_n906));
  INV_X1    g0706(.A(KEYINPUT40), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n504), .A2(new_n540), .A3(new_n544), .ZN(new_n908));
  INV_X1    g0708(.A(new_n607), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n908), .A2(new_n909), .A3(new_n663), .A4(new_n658), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n689), .A2(new_n690), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n688), .A2(KEYINPUT31), .A3(new_n651), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n797), .B1(new_n891), .B2(new_n893), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n913), .B(new_n914), .C1(new_n881), .C2(new_n882), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n914), .A2(KEYINPUT40), .A3(new_n913), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n439), .A2(KEYINPUT82), .A3(new_n451), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT82), .B1(new_n439), .B2(new_n451), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n855), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n854), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n920), .A2(new_n921), .B1(new_n862), .B2(new_n860), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n917), .B1(new_n922), .B2(KEYINPUT38), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n907), .A2(new_n915), .B1(new_n916), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n924), .A2(new_n463), .A3(new_n913), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n924), .B1(new_n463), .B2(new_n913), .ZN(new_n926));
  OR3_X1    g0726(.A1(new_n925), .A2(new_n926), .A3(new_n656), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n906), .A2(new_n927), .B1(new_n256), .B2(new_n710), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT102), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n906), .A2(new_n927), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n928), .A2(KEYINPUT102), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n845), .B1(new_n931), .B2(new_n932), .ZN(G367));
  OAI211_X1 g0733(.A(new_n544), .B(new_n540), .C1(new_n541), .C2(new_n658), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n632), .A2(new_n651), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n661), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT103), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n639), .A2(new_n651), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n504), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n625), .B2(new_n940), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n939), .B(new_n943), .Z(new_n944));
  NOR2_X1   g0744(.A1(new_n936), .A2(new_n665), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT42), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n540), .B1(new_n934), .B2(new_n576), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n946), .A2(KEYINPUT42), .B1(new_n658), .B2(new_n948), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n947), .A2(new_n949), .B1(KEYINPUT43), .B2(new_n942), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n944), .B(new_n950), .Z(new_n951));
  XOR2_X1   g0751(.A(new_n669), .B(KEYINPUT41), .Z(new_n952));
  NAND2_X1  g0752(.A1(new_n666), .A2(new_n936), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT44), .Z(new_n954));
  NOR2_X1   g0754(.A1(new_n666), .A2(new_n936), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT45), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(new_n661), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n665), .B1(new_n660), .B2(new_n664), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(new_n657), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n708), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n952), .B1(new_n962), .B2(new_n708), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n951), .B1(new_n963), .B2(new_n712), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n774), .B1(new_n208), .B2(new_n320), .C1(new_n235), .C2(new_n780), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(new_n713), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n739), .A2(G150), .B1(new_n723), .B2(G137), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n727), .A2(G68), .ZN(new_n968));
  INV_X1    g0768(.A(G159), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n743), .A2(new_n969), .B1(new_n745), .B2(new_n809), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n747), .A2(new_n201), .B1(new_n749), .B2(new_n350), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n276), .B1(new_n751), .B2(new_n202), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n967), .A2(new_n968), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n723), .A2(G317), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n306), .B1(new_n747), .B2(new_n765), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G97), .B2(new_n817), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n975), .B(new_n977), .C1(new_n585), .C2(new_n738), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n751), .A2(new_n590), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n979), .A2(KEYINPUT46), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(G311), .B2(new_n744), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n979), .A2(KEYINPUT46), .B1(G294), .B2(new_n742), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(new_n490), .C2(new_n728), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n974), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT47), .Z(new_n985));
  OAI221_X1 g0785(.A(new_n966), .B1(new_n788), .B2(new_n942), .C1(new_n985), .C2(new_n718), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n964), .A2(new_n986), .ZN(G387));
  NAND2_X1  g0787(.A1(new_n960), .A2(new_n712), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n660), .A2(new_n788), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n780), .B1(new_n230), .B2(G45), .ZN(new_n990));
  INV_X1    g0790(.A(new_n671), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n990), .B1(new_n991), .B2(new_n776), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n395), .A2(KEYINPUT50), .A3(G50), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT50), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(new_n247), .B2(new_n201), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n671), .B(new_n267), .C1(new_n203), .C2(new_n350), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n992), .A2(new_n997), .B1(G107), .B2(new_n208), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n716), .B1(new_n998), .B2(new_n774), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n727), .A2(new_n321), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT104), .B(G150), .Z(new_n1001));
  AOI22_X1  g0801(.A1(new_n739), .A2(G50), .B1(new_n723), .B2(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n751), .A2(new_n350), .B1(new_n747), .B2(new_n203), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n306), .B(new_n1003), .C1(G97), .C2(new_n817), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n247), .A2(new_n742), .B1(G159), .B2(new_n744), .ZN(new_n1005));
  AND4_X1   g0805(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n744), .A2(G322), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n585), .B2(new_n747), .C1(new_n743), .C2(new_n764), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n739), .B2(G317), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT48), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n727), .A2(G283), .B1(G294), .B2(new_n755), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT105), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1013), .A2(KEYINPUT49), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n723), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n306), .B1(new_n590), .B2(new_n749), .C1(new_n1015), .C2(new_n762), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n1013), .B2(KEYINPUT49), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1006), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n999), .B1(new_n1018), .B2(new_n718), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n961), .A2(new_n669), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n708), .A2(new_n960), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n988), .B1(new_n989), .B2(new_n1019), .C1(new_n1020), .C2(new_n1021), .ZN(G393));
  OAI221_X1 g0822(.A(new_n774), .B1(new_n485), .B2(new_n208), .C1(new_n239), .C2(new_n780), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n713), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n738), .A2(new_n969), .B1(new_n808), .B2(new_n745), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT51), .Z(new_n1026));
  OAI22_X1  g0826(.A1(new_n395), .A2(new_n747), .B1(new_n203), .B2(new_n751), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n306), .B(new_n1027), .C1(G87), .C2(new_n817), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n201), .B2(new_n743), .C1(new_n809), .C2(new_n1015), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n728), .A2(new_n350), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT106), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(KEYINPUT106), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n739), .A2(G311), .B1(G317), .B2(new_n744), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT52), .Z(new_n1035));
  OAI221_X1 g0835(.A(new_n306), .B1(new_n749), .B2(new_n490), .C1(new_n765), .C2(new_n751), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G322), .B2(new_n723), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT107), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n743), .A2(new_n585), .B1(new_n747), .B2(new_n820), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n727), .B2(G116), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1035), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1032), .A2(new_n1033), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1024), .B1(new_n1042), .B2(new_n717), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n788), .B2(new_n937), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n958), .B2(new_n711), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n962), .A2(new_n669), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n958), .A2(new_n961), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1046), .B1(new_n1047), .B2(new_n1049), .ZN(G390));
  OAI21_X1  g0850(.A(new_n713), .B1(new_n247), .B2(new_n805), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n739), .A2(G116), .B1(new_n723), .B2(G294), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n747), .A2(new_n485), .B1(new_n749), .B2(new_n203), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n276), .B(new_n1053), .C1(G87), .C2(new_n755), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n742), .A2(G107), .B1(new_n744), .B2(G283), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n755), .A2(new_n1001), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT53), .Z(new_n1058));
  NAND2_X1  g0858(.A1(new_n739), .A2(G132), .ZN(new_n1059));
  INV_X1    g0859(.A(G125), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1059), .C1(new_n1060), .C2(new_n1015), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n727), .A2(G159), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n817), .A2(G50), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(KEYINPUT54), .B(G143), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n306), .B1(new_n806), .B2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n742), .A2(G137), .B1(new_n744), .B2(G128), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1062), .A2(new_n1063), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1030), .A2(new_n1056), .B1(new_n1061), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1051), .B1(new_n1069), .B2(new_n717), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT100), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n920), .A2(new_n921), .ZN(new_n1072));
  AOI21_X1  g0872(.A(KEYINPUT38), .B1(new_n1072), .B2(new_n863), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT39), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n917), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1071), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n883), .A3(new_n878), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1070), .B1(new_n1077), .B2(new_n772), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT111), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n895), .A2(new_n850), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1080), .A2(new_n1076), .A3(new_n883), .A4(new_n878), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT108), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n894), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n891), .A2(new_n893), .A3(KEYINPUT108), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n658), .B(new_n794), .C1(new_n706), .C2(new_n631), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n795), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(new_n850), .A3(new_n923), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1081), .A2(new_n1089), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n914), .A2(G330), .A3(new_n913), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT109), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1091), .A2(KEYINPUT109), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n699), .A2(new_n799), .A3(new_n894), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1081), .B(new_n1089), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1079), .B1(new_n1099), .B2(new_n712), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n463), .A2(G330), .A3(new_n913), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n904), .B(new_n1101), .C1(new_n622), .C2(new_n623), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n913), .A2(G330), .A3(new_n799), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n1084), .A3(new_n1083), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT110), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1087), .A2(new_n795), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1103), .A2(new_n1083), .A3(KEYINPUT110), .A4(new_n1084), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1106), .A2(new_n1096), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n894), .B1(new_n699), .B2(new_n799), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n889), .B1(new_n1110), .B2(new_n1091), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1102), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1098), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1094), .A2(new_n1112), .A3(new_n1097), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n669), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1100), .A2(new_n1116), .ZN(G378));
  NAND2_X1  g0917(.A1(new_n296), .A2(new_n853), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT55), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n298), .B(new_n1119), .ZN(new_n1120));
  XOR2_X1   g0920(.A(KEYINPUT112), .B(KEYINPUT56), .Z(new_n1121));
  XNOR2_X1  g0921(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n924), .B2(G330), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n915), .A2(new_n907), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n916), .A2(new_n923), .ZN(new_n1125));
  AND4_X1   g0925(.A1(G330), .A2(new_n1124), .A3(new_n1125), .A4(new_n1122), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT101), .B1(new_n886), .B2(new_n898), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n900), .B(new_n897), .C1(new_n1077), .C2(new_n851), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1124), .A2(new_n1125), .A3(G330), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1122), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n924), .A2(G330), .A3(new_n1122), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n901), .A2(new_n902), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1130), .A2(new_n1136), .A3(KEYINPUT113), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT113), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n903), .A2(new_n1138), .A3(new_n1127), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1139), .A3(new_n712), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n713), .B1(G50), .B2(new_n805), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(G33), .A2(G41), .ZN(new_n1142));
  AOI211_X1 g0942(.A(G50), .B(new_n1142), .C1(new_n306), .C2(new_n266), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n739), .A2(G107), .B1(new_n723), .B2(G283), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n743), .A2(new_n485), .B1(new_n745), .B2(new_n590), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n320), .A2(new_n747), .B1(new_n749), .B2(new_n202), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n266), .B(new_n306), .C1(new_n751), .C2(new_n350), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1144), .A2(new_n968), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT58), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1143), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n745), .A2(new_n1060), .ZN(new_n1152));
  INV_X1    g0952(.A(G137), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n751), .A2(new_n1064), .B1(new_n747), .B2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(G132), .C2(new_n742), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n739), .A2(G128), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(new_n808), .C2(new_n728), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1142), .B1(new_n749), .B2(new_n969), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n723), .B2(G124), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1151), .B1(new_n1150), .B2(new_n1149), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1141), .B1(new_n1163), .B2(new_n717), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1122), .B2(new_n772), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1140), .A2(KEYINPUT114), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(KEYINPUT114), .B1(new_n1140), .B2(new_n1165), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1102), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1115), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT115), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT115), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1115), .A2(new_n1173), .A3(new_n1170), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT57), .B1(new_n1169), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n669), .B1(new_n1176), .B2(KEYINPUT117), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1115), .A2(new_n1173), .A3(new_n1170), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1173), .B1(new_n1115), .B2(new_n1170), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1182));
  OAI211_X1 g0982(.A(KEYINPUT117), .B(new_n1178), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT116), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1178), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n1175), .B2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1184), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1183), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1168), .B1(new_n1177), .B2(new_n1189), .ZN(G375));
  NAND2_X1  g0990(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(new_n1170), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1192), .A2(new_n952), .A3(new_n1112), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT118), .Z(new_n1194));
  OAI21_X1  g0994(.A(new_n713), .B1(G68), .B2(new_n805), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n739), .A2(G283), .B1(new_n723), .B2(G303), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n751), .A2(new_n485), .B1(new_n747), .B2(new_n490), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n276), .B(new_n1197), .C1(G77), .C2(new_n817), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n742), .A2(G116), .B1(new_n744), .B2(G294), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1196), .A2(new_n1000), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT120), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n739), .A2(G137), .B1(new_n723), .B2(G128), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n744), .A2(G132), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT121), .Z(new_n1204));
  NAND2_X1  g1004(.A1(new_n727), .A2(G50), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n276), .B1(new_n749), .B2(new_n202), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n751), .A2(new_n969), .B1(new_n747), .B2(new_n808), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n742), .C2(new_n1065), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1200), .A2(KEYINPUT120), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1201), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1195), .B1(new_n1211), .B2(new_n717), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1085), .B2(new_n772), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n711), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT119), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1213), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1215), .B2(new_n1214), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1194), .A2(new_n1217), .ZN(G381));
  INV_X1    g1018(.A(G390), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n830), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(G387), .A2(new_n1220), .A3(G396), .A4(G393), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n1217), .A3(new_n1194), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT122), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G375), .A2(G378), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(G407));
  NAND2_X1  g1025(.A1(new_n650), .A2(G213), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1224), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(G407), .A2(G213), .A3(new_n1228), .ZN(G409));
  XNOR2_X1  g1029(.A(G393), .B(new_n790), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n964), .A2(new_n986), .A3(G390), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G390), .B1(new_n964), .B2(new_n986), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1231), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1234), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT126), .Z(new_n1239));
  OAI211_X1 g1039(.A(G378), .B(new_n1168), .C1(new_n1177), .C2(new_n1189), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1130), .A2(new_n1136), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1169), .A2(new_n1175), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1165), .B1(new_n711), .B2(new_n1241), .C1(new_n1242), .C2(new_n952), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n1116), .A3(new_n1100), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1240), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1113), .A2(KEYINPUT60), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1191), .B2(new_n1170), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1113), .A2(new_n1192), .A3(KEYINPUT60), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n669), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1217), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n830), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1249), .A2(G384), .A3(new_n1217), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1245), .A2(new_n1226), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT62), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1245), .A2(new_n1226), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT123), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1251), .A2(new_n1259), .A3(new_n1253), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1227), .A2(G2897), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT123), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1260), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1263), .B1(new_n1265), .B2(new_n1261), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1258), .A2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1257), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1256), .A2(KEYINPUT62), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1239), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1235), .A2(new_n1237), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1258), .B2(new_n1266), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1227), .B1(new_n1240), .B2(new_n1244), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n1255), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1276), .B1(new_n1275), .B2(new_n1255), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1274), .B(KEYINPUT124), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1256), .A2(KEYINPUT63), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1275), .A2(new_n1276), .A3(new_n1255), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT124), .B1(new_n1283), .B2(new_n1274), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1271), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT127), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT127), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1287), .B(new_n1271), .C1(new_n1280), .C2(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(G405));
  XNOR2_X1  g1089(.A(G375), .B(G378), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(new_n1255), .ZN(new_n1291));
  XOR2_X1   g1091(.A(new_n1291), .B(new_n1239), .Z(G402));
endmodule


