//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1332, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G50), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AND2_X1   g0013(.A1(KEYINPUT64), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(KEYINPUT64), .A2(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n202), .A2(G50), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT66), .Z(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  OAI21_X1  g0027(.A(new_n210), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n213), .B1(new_n219), .B2(new_n220), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT67), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n217), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n216), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G77), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G68), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n253), .A2(G50), .B1(G20), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n249), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g0056(.A1(new_n256), .A2(KEYINPUT11), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT72), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT72), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n261), .A2(new_n258), .A3(G13), .A4(G20), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n248), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n258), .A2(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G68), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n256), .A2(KEYINPUT11), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n262), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n254), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT12), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n257), .A2(new_n265), .A3(new_n266), .A4(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT13), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT68), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(KEYINPUT68), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n276), .A2(new_n281), .A3(G226), .A4(new_n282), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n276), .A2(new_n281), .A3(G232), .A4(G1698), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n283), .B(new_n284), .C1(new_n278), .C2(new_n206), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G1), .A3(G13), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  INV_X1    g0090(.A(G45), .ZN(new_n291));
  AOI21_X1  g0091(.A(G1), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(new_n287), .A3(G274), .ZN(new_n293));
  INV_X1    g0093(.A(G238), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n293), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n272), .B1(new_n289), .B2(new_n298), .ZN(new_n299));
  AOI211_X1 g0099(.A(KEYINPUT13), .B(new_n297), .C1(new_n285), .C2(new_n288), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G179), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT14), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n303), .B(G169), .C1(new_n299), .C2(new_n300), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n289), .A2(new_n298), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT13), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n289), .A2(new_n272), .A3(new_n298), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n303), .B1(new_n309), .B2(G169), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n271), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(G200), .B1(new_n299), .B2(new_n300), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(KEYINPUT74), .B1(new_n301), .B2(G190), .ZN(new_n314));
  INV_X1    g0114(.A(new_n271), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n307), .A2(KEYINPUT74), .A3(G190), .A4(new_n308), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n276), .A2(new_n281), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(G1698), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G222), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT69), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(KEYINPUT69), .A3(G222), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n320), .A2(new_n282), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT70), .B(G223), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n327), .A2(new_n328), .B1(G77), .B2(new_n320), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n287), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n293), .ZN(new_n331));
  INV_X1    g0131(.A(new_n296), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n331), .B1(G226), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n264), .A2(G50), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n267), .A2(new_n249), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT73), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT73), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n263), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n338), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G50), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n343), .B1(new_n344), .B2(new_n268), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT8), .B(G58), .ZN(new_n346));
  INV_X1    g0146(.A(G150), .ZN(new_n347));
  INV_X1    g0147(.A(new_n253), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n250), .A2(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G20), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n349), .A2(KEYINPUT71), .B1(new_n350), .B2(new_n203), .ZN(new_n351));
  INV_X1    g0151(.A(new_n349), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT71), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n248), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n345), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n337), .B(new_n356), .C1(G169), .C2(new_n335), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n335), .A2(G190), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT9), .B1(new_n345), .B2(new_n355), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(G200), .B1(new_n330), .B2(new_n334), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n345), .A2(new_n355), .A3(KEYINPUT9), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n359), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT10), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n361), .A2(new_n363), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT10), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(new_n359), .A4(new_n362), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n358), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT15), .B(G87), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n250), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G77), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n216), .A2(new_n372), .B1(new_n346), .B2(new_n348), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n248), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n263), .A2(G77), .A3(new_n264), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n268), .A2(new_n372), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n327), .A2(G238), .B1(G107), .B2(new_n320), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n321), .A2(G232), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n287), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G244), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n293), .B1(new_n382), .B2(new_n296), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G169), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n378), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n381), .A2(new_n383), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n336), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n384), .A2(G200), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n377), .B1(new_n387), .B2(G190), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT75), .ZN(new_n394));
  INV_X1    g0194(.A(new_n346), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n264), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n340), .B2(new_n342), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n267), .A2(new_n395), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n396), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n341), .B1(new_n267), .B2(new_n249), .ZN(new_n401));
  AOI211_X1 g0201(.A(KEYINPUT73), .B(new_n248), .C1(new_n260), .C2(new_n262), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n398), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(KEYINPUT75), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n350), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n276), .B2(new_n281), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n274), .A2(new_n275), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n407), .B1(new_n216), .B2(new_n410), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n409), .A2(new_n411), .A3(new_n254), .ZN(new_n412));
  AND2_X1   g0212(.A1(G58), .A2(G68), .ZN(new_n413));
  OAI21_X1  g0213(.A(G20), .B1(new_n413), .B2(new_n201), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n253), .A2(G159), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n406), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n279), .A2(new_n350), .A3(new_n280), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n254), .B1(new_n418), .B2(KEYINPUT7), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n216), .A2(new_n410), .A3(new_n407), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n249), .B1(new_n421), .B2(KEYINPUT16), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n399), .A2(new_n405), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n282), .A2(G223), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT76), .B1(new_n410), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G87), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n278), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT3), .B(G33), .ZN(new_n428));
  AND2_X1   g0228(.A1(G226), .A2(G1698), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT76), .ZN(new_n431));
  INV_X1    g0231(.A(new_n424), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n425), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n288), .ZN(new_n435));
  INV_X1    g0235(.A(G232), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n293), .B1(new_n436), .B2(new_n296), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT77), .B1(new_n439), .B2(G179), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n385), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n437), .B1(new_n434), .B2(new_n288), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT77), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(new_n336), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT18), .B1(new_n423), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G190), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n435), .A2(new_n447), .A3(new_n438), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(G200), .B2(new_n442), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n417), .A2(new_n422), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n403), .A2(KEYINPUT75), .A3(new_n404), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT75), .B1(new_n403), .B2(new_n404), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n449), .B(new_n450), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT17), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  AOI211_X1 g0257(.A(G179), .B(new_n437), .C1(new_n434), .C2(new_n288), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n458), .A2(new_n443), .B1(new_n439), .B2(new_n385), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n456), .A2(new_n457), .A3(new_n440), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n399), .A2(new_n405), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n461), .A2(KEYINPUT17), .A3(new_n450), .A4(new_n449), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n446), .A2(new_n455), .A3(new_n460), .A4(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n393), .B1(KEYINPUT78), .B2(new_n463), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n463), .A2(KEYINPUT78), .ZN(new_n465));
  AND4_X1   g0265(.A1(new_n319), .A2(new_n369), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT81), .ZN(new_n468));
  OAI211_X1 g0268(.A(G244), .B(new_n282), .C1(new_n274), .C2(new_n275), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT4), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n469), .A2(new_n470), .B1(G33), .B2(G283), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n276), .A2(new_n281), .A3(G250), .A4(G1698), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n470), .A2(new_n382), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n276), .A2(new_n281), .A3(new_n282), .A4(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n288), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n291), .A2(G1), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n477), .A2(G274), .A3(new_n287), .A4(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  NOR2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n258), .A2(G45), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n287), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G257), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n479), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n476), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n385), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(KEYINPUT80), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT80), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n491), .B(new_n479), .C1(new_n484), .C2(new_n485), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n476), .A2(new_n336), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n258), .A2(G33), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n206), .B1(new_n263), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT79), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n267), .A2(new_n206), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n499), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT79), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n207), .A2(KEYINPUT6), .A3(G97), .ZN(new_n503));
  XOR2_X1   g0303(.A(G97), .B(G107), .Z(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n505));
  OR2_X1    g0305(.A1(KEYINPUT64), .A2(G20), .ZN(new_n506));
  NAND2_X1  g0306(.A1(KEYINPUT64), .A2(G20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n505), .A2(new_n508), .B1(G77), .B2(new_n253), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT7), .B1(new_n508), .B2(new_n428), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n276), .A2(new_n281), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(new_n408), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n509), .B1(new_n512), .B2(new_n207), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n500), .A2(new_n502), .B1(new_n513), .B2(new_n248), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n468), .B1(new_n494), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n500), .A2(new_n502), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(new_n248), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(KEYINPUT81), .A3(new_n493), .A4(new_n489), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n476), .A2(new_n490), .A3(new_n492), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n514), .B(new_n521), .C1(new_n447), .C2(new_n488), .ZN(new_n522));
  NAND3_X1  g0322(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n506), .A2(new_n507), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(G87), .B2(new_n208), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n506), .A2(G33), .A3(G97), .A4(new_n507), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT19), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n216), .A2(new_n428), .A3(G68), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n525), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(new_n248), .B1(new_n268), .B2(new_n370), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n263), .A2(G87), .A3(new_n495), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n287), .A2(G250), .A3(new_n483), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n287), .A2(G274), .A3(new_n478), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G116), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(G238), .A2(G1698), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n382), .B2(G1698), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n538), .B1(new_n540), .B2(new_n428), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n536), .B(G190), .C1(new_n287), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n294), .A2(new_n282), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n382), .A2(G1698), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(new_n274), .C2(new_n275), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n287), .B1(new_n545), .B2(new_n537), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n534), .A2(new_n535), .ZN(new_n547));
  OAI21_X1  g0347(.A(G200), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n542), .A2(new_n548), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n546), .A2(new_n547), .A3(G179), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n536), .B1(new_n287), .B2(new_n541), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n550), .B1(new_n385), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n370), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n263), .A2(new_n553), .A3(new_n495), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n531), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n533), .A2(new_n549), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n515), .A2(new_n519), .A3(new_n522), .A4(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(G116), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n268), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n263), .A2(G116), .A3(new_n495), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n278), .A2(G97), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G283), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n506), .A2(new_n561), .A3(new_n507), .A4(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n247), .A2(new_n217), .B1(G20), .B2(new_n558), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT20), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n563), .A2(KEYINPUT20), .A3(new_n564), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n559), .B(new_n560), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G303), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n276), .B2(new_n281), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n485), .A2(new_n282), .ZN(new_n570));
  INV_X1    g0370(.A(G264), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G1698), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(new_n572), .C1(new_n274), .C2(new_n275), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n288), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G270), .B(new_n287), .C1(new_n482), .C2(new_n483), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n576), .A2(new_n479), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n567), .A2(new_n578), .A3(G169), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(G200), .ZN(new_n582));
  INV_X1    g0382(.A(new_n567), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n575), .A2(new_n577), .A3(G190), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n575), .A2(new_n577), .A3(G179), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n567), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n567), .A2(new_n578), .A3(KEYINPUT21), .A4(G169), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n581), .A2(new_n585), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n263), .A2(G107), .A3(new_n495), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n260), .A2(new_n207), .A3(new_n262), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT25), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT22), .B1(new_n511), .B2(G87), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n216), .A2(new_n428), .A3(KEYINPUT22), .A4(G87), .ZN(new_n596));
  AND2_X1   g0396(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n597));
  NOR2_X1   g0397(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n597), .A2(new_n598), .B1(new_n350), .B2(G107), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n508), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n538), .A2(new_n350), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n596), .A2(new_n599), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT24), .B1(new_n595), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT22), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n320), .B2(new_n426), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n601), .A2(new_n599), .A3(new_n602), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT24), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .A4(new_n596), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n594), .B1(new_n610), .B2(new_n248), .ZN(new_n611));
  OAI211_X1 g0411(.A(G264), .B(new_n287), .C1(new_n482), .C2(new_n483), .ZN(new_n612));
  INV_X1    g0412(.A(G294), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n278), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(G250), .A2(G1698), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n485), .B2(G1698), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n616), .B2(new_n428), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n479), .B(new_n612), .C1(new_n617), .C2(new_n287), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT83), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n619), .A3(G169), .ZN(new_n620));
  INV_X1    g0420(.A(new_n615), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n485), .A2(G1698), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n621), .B(new_n622), .C1(new_n274), .C2(new_n275), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n288), .B1(new_n624), .B2(new_n614), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n625), .A2(G179), .A3(new_n479), .A4(new_n612), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n619), .B1(new_n618), .B2(G169), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT84), .B1(new_n611), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT84), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n249), .B1(new_n604), .B2(new_n609), .ZN(new_n632));
  OAI221_X1 g0432(.A(new_n631), .B1(new_n627), .B2(new_n628), .C1(new_n632), .C2(new_n594), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n618), .A2(KEYINPUT85), .A3(G190), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n618), .A2(G190), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT85), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(G200), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n618), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n634), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n611), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n630), .A2(new_n633), .A3(new_n641), .ZN(new_n642));
  NOR4_X1   g0442(.A1(new_n467), .A2(new_n557), .A3(new_n589), .A4(new_n642), .ZN(G372));
  NAND2_X1  g0443(.A1(new_n365), .A2(new_n368), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n455), .A2(new_n462), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n313), .A2(KEYINPUT74), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n447), .B2(new_n309), .ZN(new_n647));
  INV_X1    g0447(.A(new_n317), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n388), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n377), .B1(new_n387), .B2(G169), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n645), .B1(new_n653), .B2(new_n311), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n446), .A2(new_n460), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n644), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(new_n357), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n530), .A2(new_n248), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n268), .A2(new_n370), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n658), .A2(new_n659), .A3(new_n554), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n385), .B1(new_n546), .B2(new_n547), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n551), .B2(G179), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n531), .A2(new_n532), .A3(new_n542), .A4(new_n548), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n660), .B2(new_n662), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n494), .A2(new_n665), .A3(new_n514), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n663), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n665), .B1(new_n515), .B2(new_n519), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n611), .A2(new_n629), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n581), .A2(new_n587), .A3(new_n588), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n665), .B1(new_n640), .B2(new_n611), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n515), .A3(new_n519), .A4(new_n522), .ZN(new_n674));
  OAI221_X1 g0474(.A(new_n668), .B1(new_n669), .B2(new_n667), .C1(new_n672), .C2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n657), .B1(new_n467), .B2(new_n676), .ZN(G369));
  OR2_X1    g0477(.A1(new_n589), .A2(KEYINPUT86), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n258), .A2(G13), .ZN(new_n679));
  OR3_X1    g0479(.A1(new_n508), .A2(KEYINPUT27), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT27), .B1(new_n508), .B2(new_n679), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n583), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n589), .B2(KEYINPUT86), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n581), .A2(new_n587), .A3(new_n588), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n678), .A2(new_n687), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n642), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n611), .B2(new_n685), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n670), .A2(new_n684), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n671), .A2(new_n685), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n642), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n684), .B(KEYINPUT87), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n698), .B1(new_n670), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n696), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n211), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G1), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n426), .A2(new_n206), .A3(new_n207), .A4(new_n558), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n706), .A2(new_n707), .B1(new_n220), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n486), .B1(new_n475), .B2(new_n288), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n612), .B1(new_n617), .B2(new_n287), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n551), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n586), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n551), .A2(new_n618), .A3(new_n336), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n520), .A2(new_n716), .A3(new_n578), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n586), .A2(new_n712), .A3(new_n710), .A4(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(KEYINPUT31), .B(new_n699), .C1(new_n715), .C2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT88), .B1(new_n713), .B2(new_n714), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n719), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n713), .A2(KEYINPUT88), .A3(new_n714), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n685), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n720), .B1(new_n725), .B2(KEYINPUT31), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n688), .A2(new_n585), .A3(new_n700), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n557), .A2(new_n642), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(G330), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT89), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n723), .A2(new_n721), .A3(new_n719), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n732), .B1(new_n733), .B2(new_n685), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n589), .A2(new_n699), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n630), .A3(new_n633), .A4(new_n641), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n734), .B(new_n720), .C1(new_n557), .C2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(KEYINPUT89), .A3(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n731), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT29), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n668), .B1(new_n667), .B2(new_n669), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n674), .A2(new_n672), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n740), .B(new_n700), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  AND4_X1   g0543(.A1(new_n515), .A2(new_n673), .A3(new_n519), .A4(new_n522), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n630), .A2(new_n633), .A3(new_n688), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n663), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n489), .A2(new_n493), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n747), .A2(new_n556), .A3(KEYINPUT26), .A4(new_n518), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT90), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n494), .A2(new_n514), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT90), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT26), .A4(new_n556), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n749), .B(new_n752), .C1(new_n669), .C2(KEYINPUT26), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n684), .B1(new_n746), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n743), .B1(new_n754), .B2(new_n740), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n739), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT91), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(KEYINPUT91), .B1(new_n739), .B2(new_n755), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n709), .B1(new_n760), .B2(G1), .ZN(G364));
  INV_X1    g0561(.A(G13), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n508), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G45), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(new_n705), .A3(G1), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT92), .Z(new_n766));
  NOR2_X1   g0566(.A1(new_n691), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n689), .A2(G330), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT93), .Z(new_n771));
  OR3_X1    g0571(.A1(new_n689), .A2(G20), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n217), .B1(G20), .B2(new_n385), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n703), .A2(new_n428), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G45), .B2(new_n220), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n245), .B2(G45), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n511), .A2(G355), .A3(new_n211), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G116), .B2(new_n211), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n775), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n766), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT32), .ZN(new_n783));
  NOR3_X1   g0583(.A1(G179), .A2(G190), .A3(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n508), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G159), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n216), .A2(new_n336), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n447), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G58), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n783), .A2(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n783), .B2(new_n787), .ZN(new_n793));
  NOR4_X1   g0593(.A1(new_n350), .A2(new_n447), .A3(new_n638), .A4(G179), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G87), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n511), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n508), .A2(new_n336), .A3(new_n447), .A4(G200), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(G107), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G190), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n788), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n216), .B1(new_n336), .B2(new_n789), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n802), .A2(G77), .B1(new_n804), .B2(G97), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n788), .A2(G200), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n447), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(G190), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G50), .A2(new_n807), .B1(new_n808), .B2(G68), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n793), .A2(new_n799), .A3(new_n805), .A4(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G311), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n801), .A2(new_n811), .B1(new_n803), .B2(new_n613), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G326), .B2(new_n807), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT94), .Z(new_n814));
  INV_X1    g0614(.A(new_n785), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n798), .A2(G283), .B1(new_n815), .B2(G329), .ZN(new_n816));
  INV_X1    g0616(.A(new_n794), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n320), .C1(new_n568), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n790), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(G322), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n808), .ZN(new_n821));
  XOR2_X1   g0621(.A(KEYINPUT33), .B(G317), .Z(new_n822));
  OAI21_X1  g0622(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n810), .B1(new_n814), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n782), .B1(new_n824), .B2(new_n774), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n767), .A2(new_n769), .B1(new_n772), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  OR2_X1    g0627(.A1(new_n774), .A2(new_n770), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n766), .B1(G77), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n320), .B1(new_n817), .B2(new_n207), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n797), .A2(new_n426), .B1(new_n785), .B2(new_n811), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n830), .B(new_n831), .C1(G283), .C2(new_n808), .ZN(new_n832));
  INV_X1    g0632(.A(new_n807), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n568), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n802), .A2(G116), .B1(new_n804), .B2(G97), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n613), .B2(new_n790), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT95), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n802), .A2(G159), .B1(new_n819), .B2(G143), .ZN(new_n839));
  INV_X1    g0639(.A(G137), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(new_n833), .B2(new_n840), .C1(new_n347), .C2(new_n821), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT34), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n797), .A2(new_n254), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n428), .B1(new_n785), .B2(new_n846), .C1(new_n817), .C2(new_n344), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n845), .B(new_n847), .C1(G58), .C2(new_n804), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n843), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n838), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n829), .B1(new_n850), .B2(new_n774), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT96), .Z(new_n852));
  NAND3_X1  g0652(.A1(new_n386), .A2(new_n388), .A3(new_n685), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n390), .A2(new_n391), .B1(new_n377), .B2(new_n684), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n854), .B1(new_n389), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n771), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT97), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n700), .B(new_n853), .C1(new_n855), .C2(new_n652), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n741), .B2(new_n742), .ZN(new_n863));
  INV_X1    g0663(.A(new_n857), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n676), .B2(new_n699), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n739), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(new_n766), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n739), .A2(new_n863), .A3(new_n865), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n860), .A2(new_n869), .ZN(G384));
  NOR2_X1   g0670(.A1(new_n763), .A2(new_n258), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n755), .A2(new_n466), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n657), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT105), .Z(new_n874));
  NAND2_X1  g0674(.A1(new_n312), .A2(new_n685), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n419), .A2(new_n420), .ZN(new_n876));
  INV_X1    g0676(.A(new_n416), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(KEYINPUT16), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n248), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n421), .A2(KEYINPUT16), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n403), .B(new_n404), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n682), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n655), .B2(new_n645), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT100), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n463), .A2(KEYINPUT100), .A3(new_n884), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n459), .A2(new_n881), .A3(new_n440), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(new_n453), .A3(new_n883), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT101), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT37), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n442), .A2(new_n443), .A3(new_n336), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n443), .B1(new_n442), .B2(new_n336), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n442), .A2(G169), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n456), .B1(new_n896), .B2(new_n882), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(new_n898), .A3(new_n453), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n892), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT101), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n887), .A2(new_n888), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT39), .B1(new_n903), .B2(KEYINPUT38), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT103), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n445), .A2(new_n682), .B1(new_n461), .B2(new_n450), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n906), .B2(KEYINPUT102), .ZN(new_n907));
  INV_X1    g0707(.A(new_n453), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT102), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n897), .B(new_n453), .C1(new_n911), .C2(new_n898), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n905), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT104), .ZN(new_n915));
  INV_X1    g0715(.A(new_n462), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT17), .B1(new_n423), .B2(new_n449), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n446), .A2(new_n460), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n455), .A2(KEYINPUT104), .A3(new_n462), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n456), .A2(new_n882), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n897), .A2(new_n453), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n896), .A2(new_n456), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n911), .A3(new_n922), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(KEYINPUT37), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(KEYINPUT103), .A3(new_n912), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n914), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT38), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n904), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n887), .A2(new_n888), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n902), .A2(new_n899), .A3(new_n892), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n463), .A2(KEYINPUT100), .A3(new_n884), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT100), .B1(new_n463), .B2(new_n884), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n935), .B(KEYINPUT38), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT39), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n875), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT99), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n854), .B1(new_n675), .B2(new_n862), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT98), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n315), .A2(new_n685), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT14), .B1(new_n301), .B2(new_n385), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(new_n302), .A3(new_n304), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n945), .B(new_n946), .C1(new_n318), .C2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n946), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n649), .A2(new_n311), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n305), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n953), .B(new_n947), .C1(new_n314), .C2(new_n317), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n945), .B1(new_n954), .B2(new_n946), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n943), .B1(new_n944), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n863), .A2(new_n853), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n946), .B1(new_n318), .B2(new_n948), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT98), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(new_n951), .A3(new_n949), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n961), .A3(KEYINPUT99), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n931), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n939), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n957), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n919), .A2(new_n882), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n942), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n874), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n928), .A2(new_n912), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n970), .A2(new_n905), .B1(new_n921), .B2(new_n923), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT38), .B1(new_n971), .B2(new_n929), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n940), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n722), .A2(new_n724), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n974), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n975), .B(new_n734), .C1(new_n557), .C2(new_n736), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n857), .B(new_n976), .C1(new_n952), .C2(new_n955), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(KEYINPUT40), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n977), .B1(new_n964), .B2(new_n939), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n973), .A2(new_n979), .B1(new_n980), .B2(KEYINPUT40), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n975), .A2(new_n734), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(new_n728), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n981), .B1(new_n467), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n965), .A2(new_n978), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT40), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n932), .A2(new_n939), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n988), .A2(KEYINPUT40), .A3(new_n978), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n987), .A2(new_n989), .A3(new_n466), .A4(new_n976), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n984), .A2(G330), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n871), .B1(new_n969), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n969), .B2(new_n991), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n994), .A2(G116), .A3(new_n218), .A4(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT36), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n220), .A2(new_n372), .A3(new_n413), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n254), .A2(G50), .ZN(new_n999));
  OAI211_X1 g0799(.A(G1), .B(new_n762), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n993), .A2(new_n997), .A3(new_n1000), .ZN(G367));
  NAND2_X1  g0801(.A1(new_n764), .A2(G1), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT111), .Z(new_n1003));
  INV_X1    g0803(.A(KEYINPUT44), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n699), .A2(new_n518), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n515), .A2(new_n519), .A3(new_n522), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n750), .A2(new_n699), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1004), .B1(new_n701), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n698), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n670), .A2(new_n700), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1008), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(KEYINPUT44), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT45), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n701), .A2(KEYINPUT45), .A3(new_n1008), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1020), .A2(new_n691), .A3(new_n695), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1015), .A2(new_n1019), .A3(new_n696), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1010), .A2(KEYINPUT110), .ZN(new_n1024));
  AND3_X1   g0824(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1010), .A2(KEYINPUT110), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(new_n691), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n760), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n704), .B(KEYINPUT41), .Z(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1003), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1008), .A2(new_n698), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT107), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT107), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT42), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1034), .A2(KEYINPUT42), .A3(new_n1035), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n630), .A2(new_n633), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1008), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n515), .A2(new_n519), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n699), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1040), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n533), .A2(new_n685), .ZN(new_n1048));
  MUX2_X1   g0848(.A(new_n556), .B(new_n663), .S(new_n1048), .Z(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT106), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT43), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1047), .A2(KEYINPUT108), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT108), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1045), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1051), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT43), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1054), .A2(new_n1057), .A3(new_n1050), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1052), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT109), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT109), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1052), .A2(new_n1056), .A3(new_n1061), .A4(new_n1058), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n696), .A2(new_n1013), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1032), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1060), .A2(new_n1064), .A3(new_n1062), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n234), .A2(new_n703), .A3(new_n428), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n775), .B1(new_n211), .B2(new_n370), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n766), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(G283), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n801), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n794), .A2(G116), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT46), .Z(new_n1075));
  AOI211_X1 g0875(.A(new_n1073), .B(new_n1075), .C1(G107), .C2(new_n804), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n428), .B1(new_n815), .B2(G317), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n798), .A2(G97), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT113), .Z(new_n1080));
  OAI211_X1 g0880(.A(new_n1076), .B(new_n1080), .C1(new_n613), .C2(new_n821), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n807), .A2(G311), .B1(new_n819), .B2(G303), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT112), .Z(new_n1083));
  NAND2_X1  g0883(.A1(new_n804), .A2(G68), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n790), .B2(new_n347), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT114), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n797), .A2(new_n372), .B1(new_n785), .B2(new_n840), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n320), .B(new_n1087), .C1(G58), .C2(new_n794), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G143), .A2(new_n807), .B1(new_n808), .B2(G159), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(new_n344), .C2(new_n801), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1081), .A2(new_n1083), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g0891(.A(KEYINPUT115), .B(KEYINPUT47), .Z(new_n1092));
  XNOR2_X1  g0892(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1071), .B1(new_n1093), .B2(new_n774), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1050), .A2(new_n773), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1068), .A2(new_n1096), .ZN(G387));
  AOI21_X1  g0897(.A(new_n1028), .B1(new_n758), .B2(new_n759), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n758), .A2(new_n1028), .A3(new_n759), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n704), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1028), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n693), .A2(new_n694), .A3(new_n773), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n238), .A2(new_n291), .ZN(new_n1104));
  AOI211_X1 g0904(.A(G45), .B(new_n707), .C1(G68), .C2(G77), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n395), .A2(KEYINPUT50), .A3(new_n344), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT50), .B1(new_n395), .B2(new_n344), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1108), .A2(new_n776), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT116), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n511), .A2(new_n211), .A3(new_n707), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(G107), .B2(new_n211), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1104), .A2(new_n1109), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n775), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n766), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n428), .B1(new_n815), .B2(G326), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n803), .A2(new_n1072), .B1(new_n817), .B2(new_n613), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n802), .A2(G303), .B1(new_n819), .B2(G317), .ZN(new_n1119));
  INV_X1    g0919(.A(G322), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1119), .B1(new_n833), .B2(new_n1120), .C1(new_n811), .C2(new_n821), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT48), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1118), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n1122), .B2(new_n1121), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT49), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1117), .B1(new_n558), .B2(new_n797), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n803), .A2(new_n370), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n801), .B2(new_n254), .C1(new_n344), .C2(new_n790), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n794), .A2(G77), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1078), .A2(new_n428), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G150), .B2(new_n815), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n786), .B2(new_n833), .C1(new_n346), .C2(new_n821), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n1126), .A2(new_n1127), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1116), .B1(new_n1135), .B2(new_n774), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1102), .A2(new_n1003), .B1(new_n1103), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1101), .A2(new_n1137), .ZN(G393));
  NAND2_X1  g0938(.A1(new_n1013), .A2(new_n773), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n775), .B1(new_n206), .B2(new_n211), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n242), .A2(new_n776), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n766), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n428), .B1(new_n797), .B2(new_n426), .C1(new_n254), .C2(new_n817), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G143), .B2(new_n815), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n802), .A2(new_n395), .B1(new_n804), .B2(G77), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n344), .C2(new_n821), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n807), .A2(G150), .B1(new_n819), .B2(G159), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT51), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n807), .A2(G317), .B1(new_n819), .B2(G311), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT52), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n801), .A2(new_n613), .B1(new_n803), .B2(new_n558), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n320), .B1(new_n817), .B2(new_n1072), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n797), .A2(new_n207), .B1(new_n785), .B2(new_n1120), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n568), .B2(new_n821), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1146), .A2(new_n1148), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1142), .B1(new_n1156), .B2(new_n774), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1139), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1003), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1023), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1099), .A2(new_n1023), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1023), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n705), .B1(new_n1098), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1160), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(G390));
  OAI21_X1  g0965(.A(new_n875), .B1(new_n944), .B2(new_n956), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n933), .A2(new_n941), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n856), .A2(new_n389), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n753), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n745), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n1170), .A2(new_n674), .B1(new_n660), .B2(new_n662), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n685), .B(new_n1168), .C1(new_n1169), .C2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n853), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n961), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n988), .A2(new_n1174), .A3(new_n875), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n729), .A2(new_n730), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT89), .B1(new_n737), .B2(G330), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n857), .B(new_n961), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1167), .A2(new_n1175), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n976), .A2(G330), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n857), .A3(new_n961), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1167), .B2(new_n1175), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n1003), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(KEYINPUT39), .A2(new_n965), .B1(new_n904), .B2(new_n932), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n771), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n766), .B1(new_n395), .B2(new_n828), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT118), .Z(new_n1190));
  INV_X1    g0990(.A(new_n774), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n845), .B1(G294), .B2(new_n815), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n320), .A3(new_n795), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n207), .A2(new_n821), .B1(new_n833), .B2(new_n1072), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(G97), .C2(new_n802), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n790), .A2(new_n558), .B1(new_n803), .B2(new_n372), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT120), .ZN(new_n1197));
  INV_X1    g0997(.A(G125), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n511), .B1(new_n1198), .B2(new_n785), .C1(new_n344), .C2(new_n797), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT119), .Z(new_n1200));
  INV_X1    g1000(.A(G128), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1201), .A2(new_n833), .B1(new_n821), .B2(new_n840), .ZN(new_n1202));
  OR3_X1    g1002(.A1(new_n817), .A2(KEYINPUT53), .A3(new_n347), .ZN(new_n1203));
  OAI21_X1  g1003(.A(KEYINPUT53), .B1(new_n817), .B2(new_n347), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT54), .B(G143), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1204), .C1(new_n801), .C2(new_n1205), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n790), .A2(new_n846), .B1(new_n803), .B2(new_n786), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1202), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1195), .A2(new_n1197), .B1(new_n1200), .B2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1188), .B(new_n1190), .C1(new_n1191), .C2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1185), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT117), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1167), .A2(new_n1175), .A3(new_n1178), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n875), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n932), .B2(new_n939), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1186), .A2(new_n1166), .B1(new_n1174), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1213), .B1(new_n1216), .B2(new_n1182), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n854), .B1(new_n754), .B2(new_n1168), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n976), .A2(G330), .A3(new_n857), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n956), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1178), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n956), .A2(new_n1180), .A3(new_n864), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n857), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1222), .B1(new_n1223), .B2(new_n956), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1221), .B1(new_n1224), .B2(new_n944), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n466), .A2(new_n1181), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n872), .A2(new_n1226), .A3(new_n657), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1212), .B1(new_n1217), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n864), .B1(new_n731), .B2(new_n738), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1182), .B1(new_n1231), .B2(new_n961), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n958), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1227), .B1(new_n1233), .B2(new_n1221), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT39), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n939), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n972), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n964), .B2(new_n939), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1214), .B1(new_n958), .B2(new_n961), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n875), .B1(new_n972), .B2(new_n940), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1218), .A2(new_n956), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1222), .B1(new_n1240), .B2(new_n1243), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1234), .A2(new_n1244), .A3(KEYINPUT117), .A4(new_n1213), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1230), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n705), .B1(new_n1217), .B2(new_n1229), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1211), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(G378));
  AOI21_X1  g1049(.A(new_n682), .B1(new_n345), .B2(new_n355), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n369), .B(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1251), .B(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1187), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n766), .B1(G50), .B2(new_n828), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n819), .A2(G128), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n802), .A2(G137), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1259), .B1(new_n347), .B2(new_n803), .C1(new_n817), .C2(new_n1205), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1198), .A2(new_n833), .B1(new_n821), .B2(new_n846), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1263), .A2(KEYINPUT59), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(KEYINPUT59), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n278), .B(new_n290), .C1(new_n797), .C2(new_n786), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(G124), .B2(new_n815), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1264), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1084), .B1(new_n801), .B2(new_n370), .C1(new_n207), .C2(new_n790), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n798), .A2(G58), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n428), .A2(G41), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n1131), .A3(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G283), .B2(new_n815), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n206), .B2(new_n821), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1269), .B(new_n1274), .C1(G116), .C2(new_n807), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT58), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1275), .A2(KEYINPUT58), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1271), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1278), .B(new_n344), .C1(G33), .C2(G41), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1268), .A2(new_n1276), .A3(new_n1277), .A4(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1256), .B1(new_n1280), .B2(new_n774), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1255), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(G330), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1254), .B1(new_n981), .B2(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1251), .B(new_n1252), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1285), .A2(new_n987), .A3(new_n989), .A4(G330), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1284), .A2(new_n968), .A3(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n968), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1282), .B1(new_n1289), .B2(new_n1159), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT117), .B1(new_n1184), .B2(new_n1234), .ZN(new_n1292));
  AND4_X1   g1092(.A1(KEYINPUT117), .A2(new_n1234), .A3(new_n1244), .A4(new_n1213), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1228), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT57), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1227), .B1(new_n1230), .B2(new_n1245), .ZN(new_n1297));
  OAI21_X1  g1097(.A(KEYINPUT57), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n704), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1291), .B1(new_n1296), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT121), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1300), .A2(KEYINPUT121), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(G375));
  OAI211_X1 g1104(.A(new_n1227), .B(new_n1221), .C1(new_n1224), .C2(new_n944), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1229), .A2(new_n1031), .A3(new_n1305), .ZN(new_n1306));
  OAI221_X1 g1106(.A(new_n1129), .B1(new_n801), .B2(new_n207), .C1(new_n1072), .C2(new_n790), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n511), .B1(G97), .B2(new_n794), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n798), .A2(G77), .B1(new_n815), .B2(G303), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1308), .B(new_n1309), .C1(new_n821), .C2(new_n558), .ZN(new_n1310));
  AOI211_X1 g1110(.A(new_n1307), .B(new_n1310), .C1(G294), .C2(new_n807), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1270), .B(new_n428), .C1(new_n347), .C2(new_n801), .ZN(new_n1312));
  OAI22_X1  g1112(.A1(new_n817), .A2(new_n786), .B1(new_n1201), .B2(new_n785), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1313), .B(KEYINPUT123), .ZN(new_n1314));
  AOI211_X1 g1114(.A(new_n1312), .B(new_n1314), .C1(G50), .C2(new_n804), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1315), .B(KEYINPUT124), .ZN(new_n1316));
  OAI22_X1  g1116(.A1(new_n821), .A2(new_n1205), .B1(new_n840), .B2(new_n790), .ZN(new_n1317));
  OR3_X1    g1117(.A1(new_n833), .A2(KEYINPUT122), .A3(new_n846), .ZN(new_n1318));
  OAI21_X1  g1118(.A(KEYINPUT122), .B1(new_n833), .B2(new_n846), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1317), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1311), .B1(new_n1316), .B2(new_n1320), .ZN(new_n1321));
  OAI221_X1 g1121(.A(new_n766), .B1(G68), .B2(new_n828), .C1(new_n1321), .C2(new_n1191), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(new_n956), .B2(new_n770), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1323), .B1(new_n1225), .B2(new_n1003), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1306), .A2(new_n1324), .ZN(G381));
  NAND3_X1  g1125(.A1(new_n1101), .A2(new_n826), .A3(new_n1137), .ZN(new_n1326));
  NOR4_X1   g1126(.A1(G390), .A2(new_n1326), .A3(G381), .A4(G384), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1096), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1328), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1327), .A2(new_n1329), .A3(new_n1248), .ZN(new_n1330));
  OR2_X1    g1130(.A1(G375), .A2(new_n1330), .ZN(G407));
  OAI21_X1  g1131(.A(new_n1248), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1332));
  OAI211_X1 g1132(.A(G407), .B(G213), .C1(G343), .C2(new_n1332), .ZN(G409));
  INV_X1    g1133(.A(KEYINPUT63), .ZN(new_n1334));
  OAI211_X1 g1134(.A(G378), .B(new_n1291), .C1(new_n1296), .C2(new_n1299), .ZN(new_n1335));
  NOR3_X1   g1135(.A1(new_n1297), .A2(new_n1030), .A3(new_n1289), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1248), .B1(new_n1336), .B2(new_n1290), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n683), .A2(G213), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT125), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT60), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1341), .B1(new_n1305), .B2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n705), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1344));
  AND2_X1   g1144(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1345));
  AOI22_X1  g1145(.A1(new_n1232), .A2(new_n958), .B1(new_n1345), .B2(new_n1178), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1346), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n1227), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1305), .A2(new_n1342), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1343), .A2(new_n1344), .A3(new_n1347), .A4(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1324), .ZN(new_n1350));
  INV_X1    g1150(.A(G384), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1349), .A2(G384), .A3(new_n1324), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1334), .B1(new_n1340), .B2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1339), .ZN(new_n1356));
  AND3_X1   g1156(.A1(new_n1349), .A2(G384), .A3(new_n1324), .ZN(new_n1357));
  AOI21_X1  g1157(.A(G384), .B1(new_n1349), .B2(new_n1324), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  OAI211_X1 g1159(.A(G2897), .B(new_n1356), .C1(new_n1359), .C2(KEYINPUT126), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT126), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1356), .A2(G2897), .ZN(new_n1362));
  OAI211_X1 g1162(.A(new_n1361), .B(new_n1362), .C1(new_n1357), .C2(new_n1358), .ZN(new_n1363));
  AOI22_X1  g1163(.A1(new_n1360), .A2(new_n1363), .B1(KEYINPUT126), .B2(new_n1359), .ZN(new_n1364));
  AOI21_X1  g1164(.A(KEYINPUT61), .B1(new_n1340), .B2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1326), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n826), .B1(new_n1101), .B2(new_n1137), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1164), .B1(new_n1366), .B2(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1367), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1369), .A2(G390), .A3(new_n1326), .ZN(new_n1370));
  AND3_X1   g1170(.A1(new_n1329), .A2(new_n1368), .A3(new_n1370), .ZN(new_n1371));
  AOI22_X1  g1171(.A1(new_n1368), .A2(new_n1370), .B1(new_n1068), .B2(new_n1096), .ZN(new_n1372));
  NOR2_X1   g1172(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1356), .B1(new_n1335), .B2(new_n1337), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1374), .A2(KEYINPUT63), .A3(new_n1359), .ZN(new_n1375));
  NAND4_X1  g1175(.A1(new_n1355), .A2(new_n1365), .A3(new_n1373), .A4(new_n1375), .ZN(new_n1376));
  INV_X1    g1176(.A(KEYINPUT62), .ZN(new_n1377));
  AND3_X1   g1177(.A1(new_n1374), .A2(new_n1377), .A3(new_n1359), .ZN(new_n1378));
  INV_X1    g1178(.A(KEYINPUT61), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1359), .A2(KEYINPUT126), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1362), .B1(new_n1354), .B2(new_n1361), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1363), .ZN(new_n1382));
  OAI21_X1  g1182(.A(new_n1380), .B1(new_n1381), .B2(new_n1382), .ZN(new_n1383));
  OAI21_X1  g1183(.A(new_n1379), .B1(new_n1374), .B2(new_n1383), .ZN(new_n1384));
  AOI21_X1  g1184(.A(new_n1377), .B1(new_n1374), .B2(new_n1359), .ZN(new_n1385));
  NOR3_X1   g1185(.A1(new_n1378), .A2(new_n1384), .A3(new_n1385), .ZN(new_n1386));
  OAI21_X1  g1186(.A(new_n1376), .B1(new_n1386), .B2(new_n1373), .ZN(G405));
  OAI21_X1  g1187(.A(new_n1354), .B1(new_n1371), .B2(new_n1372), .ZN(new_n1388));
  INV_X1    g1188(.A(KEYINPUT127), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1368), .A2(new_n1370), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1390), .A2(G387), .ZN(new_n1391));
  NAND3_X1  g1191(.A1(new_n1329), .A2(new_n1368), .A3(new_n1370), .ZN(new_n1392));
  NAND3_X1  g1192(.A1(new_n1391), .A2(new_n1359), .A3(new_n1392), .ZN(new_n1393));
  NAND3_X1  g1193(.A1(new_n1388), .A2(new_n1389), .A3(new_n1393), .ZN(new_n1394));
  INV_X1    g1194(.A(new_n1394), .ZN(new_n1395));
  AOI21_X1  g1195(.A(new_n1389), .B1(new_n1388), .B2(new_n1393), .ZN(new_n1396));
  OR2_X1    g1196(.A1(new_n1300), .A2(KEYINPUT121), .ZN(new_n1397));
  AOI21_X1  g1197(.A(G378), .B1(new_n1397), .B2(new_n1301), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1300), .A2(G378), .ZN(new_n1399));
  INV_X1    g1199(.A(new_n1399), .ZN(new_n1400));
  OAI22_X1  g1200(.A1(new_n1395), .A2(new_n1396), .B1(new_n1398), .B2(new_n1400), .ZN(new_n1401));
  NAND2_X1  g1201(.A1(new_n1388), .A2(new_n1393), .ZN(new_n1402));
  NAND2_X1  g1202(.A1(new_n1402), .A2(KEYINPUT127), .ZN(new_n1403));
  NAND4_X1  g1203(.A1(new_n1403), .A2(new_n1332), .A3(new_n1399), .A4(new_n1394), .ZN(new_n1404));
  AND2_X1   g1204(.A1(new_n1401), .A2(new_n1404), .ZN(G402));
endmodule


