//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  NAND2_X1  g0009(.A1(G68), .A2(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  AOI211_X1 g0015(.A(new_n213), .B(new_n215), .C1(G77), .C2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n204), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT64), .ZN(new_n229));
  INV_X1    g0029(.A(G58), .ZN(new_n230));
  INV_X1    g0030(.A(G68), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n209), .B(new_n226), .C1(new_n229), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n220), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n227), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n203), .A2(G20), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n253), .A2(G50), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(G20), .B1(new_n232), .B2(G50), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n261), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n256), .B1(G50), .B2(new_n254), .C1(new_n266), .C2(new_n253), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT9), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G223), .A2(G1698), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(G1), .B(G13), .C1(new_n262), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n278), .B(new_n281), .C1(G77), .C2(new_n274), .ZN(new_n282));
  INV_X1    g0082(.A(G45), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G274), .ZN(new_n285));
  INV_X1    g0085(.A(new_n284), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n280), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n282), .B(new_n285), .C1(new_n212), .C2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n269), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT10), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n267), .A2(new_n268), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n288), .A2(G200), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n291), .A2(new_n292), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n269), .A2(new_n294), .A3(new_n290), .ZN(new_n296));
  INV_X1    g0096(.A(new_n293), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT10), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n288), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n301), .B(new_n267), .C1(G179), .C2(new_n288), .ZN(new_n302));
  INV_X1    g0102(.A(G244), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n285), .B1(new_n287), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g0104(.A(new_n304), .B(KEYINPUT66), .Z(new_n305));
  NAND2_X1  g0105(.A1(G238), .A2(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(G232), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n274), .B(new_n306), .C1(new_n307), .C2(G1698), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT67), .B(G107), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n308), .B(new_n281), .C1(new_n274), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G200), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n305), .A2(G190), .A3(new_n310), .ZN(new_n313));
  INV_X1    g0113(.A(new_n254), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT68), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT68), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n254), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n315), .A2(new_n317), .A3(new_n253), .A4(new_n255), .ZN(new_n318));
  INV_X1    g0118(.A(G77), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n265), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n321));
  INV_X1    g0121(.A(new_n263), .ZN(new_n322));
  XOR2_X1   g0122(.A(KEYINPUT15), .B(G87), .Z(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n321), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n320), .B1(new_n252), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n315), .A2(new_n317), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n319), .ZN(new_n328));
  XOR2_X1   g0128(.A(new_n328), .B(KEYINPUT69), .Z(new_n329));
  NAND4_X1  g0129(.A1(new_n312), .A2(new_n313), .A3(new_n326), .A4(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n311), .A2(new_n300), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n326), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n305), .A2(new_n333), .A3(new_n310), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AND4_X1   g0135(.A1(new_n299), .A2(new_n302), .A3(new_n330), .A4(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT70), .ZN(new_n338));
  NOR2_X1   g0138(.A1(G226), .A2(G1698), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n307), .B2(G1698), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n274), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n262), .A2(new_n222), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n338), .B(new_n281), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n274), .B2(new_n340), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT70), .B1(new_n344), .B2(new_n280), .ZN(new_n345));
  INV_X1    g0145(.A(new_n285), .ZN(new_n346));
  INV_X1    g0146(.A(new_n287), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(G238), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n343), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT13), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT13), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n343), .A2(new_n345), .A3(new_n351), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n337), .B1(new_n353), .B2(G169), .ZN(new_n354));
  AOI211_X1 g0154(.A(KEYINPUT14), .B(new_n300), .C1(new_n350), .C2(new_n352), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n353), .A2(new_n333), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n322), .A2(new_n319), .B1(new_n204), .B2(G68), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT71), .B1(new_n259), .B2(G50), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n259), .A2(KEYINPUT71), .A3(G50), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT11), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(new_n252), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT11), .B1(new_n361), .B2(new_n253), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n327), .A2(KEYINPUT12), .A3(new_n231), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n231), .B1(new_n318), .B2(KEYINPUT12), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT12), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n254), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n366), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n357), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n350), .A2(new_n352), .ZN(new_n373));
  INV_X1    g0173(.A(G200), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n350), .A2(G190), .A3(new_n352), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT77), .ZN(new_n380));
  AND2_X1   g0180(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n381));
  NOR2_X1   g0181(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n382));
  OAI21_X1  g0182(.A(G33), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n275), .A2(G223), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n270), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT75), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G87), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n383), .A2(G226), .A3(G1698), .A4(new_n270), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n383), .A2(KEYINPUT75), .A3(new_n270), .A4(new_n384), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n387), .A2(new_n388), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n281), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n285), .B1(new_n287), .B2(new_n307), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(G200), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AOI211_X1 g0195(.A(G190), .B(new_n393), .C1(new_n391), .C2(new_n281), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n380), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(new_n289), .A3(new_n394), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n393), .B1(new_n391), .B2(new_n281), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n398), .B(KEYINPUT77), .C1(G200), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n265), .A2(new_n255), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n253), .A2(new_n254), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n402), .A2(new_n403), .B1(new_n254), .B2(new_n265), .ZN(new_n404));
  XNOR2_X1  g0204(.A(G58), .B(G68), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(G20), .B1(G159), .B2(new_n259), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT7), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n383), .A2(new_n270), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n408), .B1(new_n409), .B2(new_n204), .ZN(new_n410));
  OR2_X1    g0210(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n411));
  NAND2_X1  g0211(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n262), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n270), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT73), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT73), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n383), .A2(new_n416), .A3(new_n270), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(KEYINPUT7), .A2(G20), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n410), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n407), .B1(new_n420), .B2(G68), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n253), .B1(new_n421), .B2(KEYINPUT16), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT7), .B1(new_n273), .B2(new_n204), .ZN(new_n423));
  INV_X1    g0223(.A(new_n272), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n381), .A2(new_n382), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n262), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n408), .A2(G20), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT74), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n411), .A2(new_n262), .A3(new_n412), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n272), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT74), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(new_n427), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n423), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n406), .B1(new_n434), .B2(new_n231), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT16), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n404), .B1(new_n422), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n401), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n401), .A2(new_n438), .A3(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n399), .A2(new_n300), .ZN(new_n446));
  AOI211_X1 g0246(.A(new_n333), .B(new_n393), .C1(new_n391), .C2(new_n281), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n399), .A2(G179), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n449), .B(KEYINPUT76), .C1(new_n300), .C2(new_n399), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n404), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n418), .A2(new_n419), .ZN(new_n453));
  INV_X1    g0253(.A(new_n410), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(G68), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(KEYINPUT16), .A3(new_n406), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n252), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n429), .A2(new_n433), .ZN(new_n458));
  INV_X1    g0258(.A(new_n423), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G68), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT16), .B1(new_n461), .B2(new_n406), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n452), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n451), .A2(new_n463), .A3(KEYINPUT18), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT18), .B1(new_n451), .B2(new_n463), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n336), .A2(new_n379), .A3(new_n444), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT81), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n383), .A2(new_n204), .A3(G68), .A4(new_n270), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT19), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n222), .A2(KEYINPUT78), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT78), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G97), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n471), .B1(new_n475), .B2(new_n322), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(G20), .B1(new_n342), .B2(KEYINPUT19), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT78), .B(G97), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(G87), .ZN(new_n480));
  INV_X1    g0280(.A(new_n309), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n252), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n327), .A2(new_n324), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n403), .B1(new_n203), .B2(G33), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G87), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  OR2_X1    g0287(.A1(G238), .A2(G1698), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n303), .A2(G1698), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n383), .A2(new_n270), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G116), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n280), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n283), .A2(G1), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n218), .A2(KEYINPUT80), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(G274), .ZN(new_n495));
  OAI211_X1 g0295(.A(KEYINPUT80), .B(G250), .C1(new_n283), .C2(G1), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n281), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(G200), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n469), .B1(new_n487), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n492), .A2(new_n497), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G190), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n309), .A2(new_n479), .A3(G87), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n476), .B(new_n470), .C1(new_n503), .C2(new_n478), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n504), .A2(new_n252), .B1(new_n327), .B2(new_n324), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(KEYINPUT81), .A3(new_n498), .A4(new_n486), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n500), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n485), .A2(new_n323), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n505), .A2(new_n508), .B1(new_n333), .B2(new_n501), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(G169), .B2(new_n501), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n479), .A2(KEYINPUT6), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n222), .A2(new_n512), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G97), .A2(G107), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n513), .B1(KEYINPUT6), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G20), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n260), .A2(new_n319), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n518), .B(new_n520), .C1(new_n434), .C2(new_n481), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n252), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n314), .A2(new_n222), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n485), .A2(G97), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n383), .A2(G244), .A3(new_n270), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n270), .A2(new_n272), .A3(G250), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT4), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G1698), .ZN(new_n531));
  AND2_X1   g0331(.A1(KEYINPUT4), .A2(G244), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n270), .A2(new_n272), .A3(new_n532), .A4(new_n275), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G283), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n528), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT79), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT79), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n528), .A2(new_n531), .A3(new_n538), .A4(new_n535), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n281), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(KEYINPUT5), .A2(G41), .ZN(new_n541));
  AND2_X1   g0341(.A1(KEYINPUT5), .A2(G41), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n493), .B(G274), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n493), .B1(new_n542), .B2(new_n541), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n545), .A2(new_n280), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n544), .B1(new_n546), .B2(G257), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n540), .A2(new_n333), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n540), .A2(new_n547), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n300), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n525), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n521), .A2(new_n252), .B1(G97), .B2(new_n485), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n540), .A2(new_n289), .A3(new_n547), .ZN(new_n553));
  AOI21_X1  g0353(.A(G200), .B1(new_n540), .B2(new_n547), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n552), .B(new_n523), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n511), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n219), .A2(G20), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n252), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n475), .A2(G33), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n534), .A2(new_n204), .ZN(new_n561));
  OAI211_X1 g0361(.A(KEYINPUT20), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT20), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n561), .B1(new_n479), .B2(new_n262), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n563), .B1(new_n564), .B2(new_n558), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n327), .A2(new_n219), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n219), .B1(new_n203), .B2(G33), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n315), .A2(new_n317), .A3(new_n253), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n223), .A2(new_n275), .ZN(new_n571));
  OR2_X1    g0371(.A1(new_n275), .A2(G264), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n383), .A2(new_n270), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n273), .A2(G303), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n281), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n545), .A2(G270), .A3(new_n280), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n577), .A2(KEYINPUT82), .A3(new_n543), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT82), .B1(new_n577), .B2(new_n543), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n570), .A2(new_n580), .A3(G169), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n580), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(G179), .A3(new_n570), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n570), .A2(new_n580), .A3(KEYINPUT21), .A4(G169), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n204), .A2(KEYINPUT23), .A3(G107), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n217), .A2(G20), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(new_n270), .A3(new_n272), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT22), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n383), .A2(KEYINPUT22), .A3(new_n270), .A4(new_n590), .ZN(new_n594));
  OAI21_X1  g0394(.A(KEYINPUT23), .B1(new_n309), .B2(new_n204), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n491), .A2(G20), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n593), .A2(new_n594), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT24), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n596), .B(new_n589), .C1(new_n591), .C2(new_n592), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n601), .A2(KEYINPUT24), .A3(new_n595), .A4(new_n594), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n252), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n485), .A2(G107), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n254), .A2(G107), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT84), .ZN(new_n606));
  XNOR2_X1  g0406(.A(KEYINPUT83), .B(KEYINPUT25), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n606), .ZN(new_n609));
  MUX2_X1   g0409(.A(new_n605), .B(new_n608), .S(new_n609), .Z(new_n610));
  NAND3_X1  g0410(.A1(new_n603), .A2(new_n604), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n218), .A2(new_n275), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n223), .A2(G1698), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n383), .A2(new_n270), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(G33), .A2(G294), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n280), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n545), .A2(G264), .A3(new_n280), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n616), .A2(new_n544), .A3(new_n617), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n618), .A2(KEYINPUT85), .A3(G200), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n289), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n621), .B(KEYINPUT85), .C1(G200), .C2(new_n618), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n614), .A2(new_n615), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n617), .B1(new_n624), .B2(new_n281), .ZN(new_n625));
  AOI21_X1  g0425(.A(G169), .B1(new_n625), .B2(new_n543), .ZN(new_n626));
  NOR4_X1   g0426(.A1(new_n616), .A2(G179), .A3(new_n544), .A4(new_n617), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n611), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n580), .A2(G200), .ZN(new_n630));
  INV_X1    g0430(.A(new_n570), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n630), .B(new_n631), .C1(new_n289), .C2(new_n580), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n588), .A2(new_n623), .A3(new_n629), .A4(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n468), .A2(new_n556), .A3(new_n633), .ZN(G372));
  OAI21_X1  g0434(.A(new_n449), .B1(new_n300), .B2(new_n399), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n463), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT18), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n463), .A2(KEYINPUT18), .A3(new_n635), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n375), .A2(new_n377), .ZN(new_n641));
  INV_X1    g0441(.A(new_n335), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n641), .B1(new_n372), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n640), .B1(new_n643), .B2(new_n443), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n299), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(new_n302), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n507), .A2(new_n510), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT26), .B1(new_n551), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n550), .A2(new_n548), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n505), .A2(new_n508), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT86), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n501), .B2(G169), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n490), .A2(new_n491), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n281), .ZN(new_n654));
  INV_X1    g0454(.A(new_n497), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(KEYINPUT86), .A3(new_n300), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n501), .A2(new_n333), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n650), .A2(new_n652), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n487), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n502), .A3(new_n498), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n649), .A2(new_n663), .A3(new_n664), .A4(new_n525), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n648), .A2(new_n665), .A3(new_n659), .ZN(new_n666));
  AOI21_X1  g0466(.A(G200), .B1(new_n625), .B2(new_n543), .ZN(new_n667));
  NOR4_X1   g0467(.A1(new_n616), .A2(G190), .A3(new_n544), .A4(new_n617), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT85), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n670), .A2(new_n611), .A3(new_n619), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(new_n662), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n629), .A2(new_n585), .A3(new_n586), .A4(new_n583), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n672), .A2(new_n555), .A3(new_n551), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT87), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n551), .A2(new_n555), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT87), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n676), .A2(new_n677), .A3(new_n673), .A4(new_n672), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n666), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n646), .B1(new_n468), .B2(new_n679), .ZN(G369));
  NAND3_X1  g0480(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n570), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n632), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n687), .B1(new_n587), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n587), .B2(new_n687), .ZN(new_n690));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n611), .A2(new_n686), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n623), .A2(new_n694), .B1(new_n611), .B2(new_n628), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n629), .A2(new_n686), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n686), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n587), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n696), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(G399));
  NAND2_X1  g0504(.A1(new_n503), .A2(new_n219), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n207), .A2(new_n279), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G1), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n233), .B2(new_n707), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n679), .A2(KEYINPUT29), .A3(new_n686), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  INV_X1    g0512(.A(new_n551), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n664), .A3(new_n511), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT26), .B1(new_n551), .B2(new_n662), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n674), .A2(new_n714), .A3(new_n659), .A4(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n712), .B1(new_n716), .B2(new_n700), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n501), .A2(KEYINPUT88), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n501), .A2(KEYINPUT88), .ZN(new_n720));
  NOR4_X1   g0520(.A1(new_n719), .A2(new_n584), .A3(new_n720), .A4(G179), .ZN(new_n721));
  INV_X1    g0521(.A(new_n618), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT89), .B1(new_n549), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT89), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n724), .B(new_n618), .C1(new_n540), .C2(new_n547), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n721), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT90), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n584), .A2(G179), .ZN(new_n728));
  INV_X1    g0528(.A(new_n625), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n540), .A2(new_n547), .A3(new_n501), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT30), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NOR4_X1   g0534(.A1(new_n731), .A2(new_n728), .A3(new_n734), .A4(new_n729), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT90), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n737), .B(new_n721), .C1(new_n723), .C2(new_n725), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n727), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n686), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n556), .A2(new_n633), .A3(new_n686), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n736), .ZN(new_n744));
  INV_X1    g0544(.A(new_n726), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT31), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n743), .B1(new_n700), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n718), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n710), .B1(new_n749), .B2(G1), .ZN(G364));
  NOR3_X1   g0550(.A1(new_n289), .A2(G179), .A3(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n204), .ZN(new_n752));
  INV_X1    g0552(.A(G294), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n289), .A2(new_n374), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n204), .A2(G179), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G190), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G303), .A2(new_n758), .B1(new_n761), .B2(G329), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n204), .A2(new_n333), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n759), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n755), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT93), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n767), .A2(new_n768), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n754), .B(new_n766), .C1(G326), .C2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n764), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n374), .A2(G190), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(KEYINPUT33), .B(G317), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n274), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  INV_X1    g0582(.A(new_n756), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G322), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n775), .A2(new_n289), .A3(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n781), .B1(new_n782), .B2(new_n785), .C1(new_n786), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n752), .A2(new_n222), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G68), .B2(new_n778), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n757), .A2(new_n217), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n765), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G77), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n788), .A2(new_n230), .B1(new_n785), .B2(new_n512), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G50), .B2(new_n773), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n792), .A2(new_n794), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G159), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n760), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT32), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n274), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n789), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n204), .B1(KEYINPUT92), .B2(new_n300), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n300), .A2(KEYINPUT92), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n227), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G13), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(G20), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G45), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n707), .A2(G1), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n418), .A2(new_n207), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT91), .Z(new_n815));
  NAND2_X1  g0615(.A1(new_n249), .A2(G45), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(G45), .C2(new_n233), .ZN(new_n817));
  INV_X1    g0617(.A(G355), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n207), .A2(new_n274), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(G116), .B2(new_n207), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G13), .A2(G33), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n204), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n807), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n808), .A2(new_n813), .A3(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT95), .Z(new_n827));
  NAND2_X1  g0627(.A1(new_n690), .A2(new_n823), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n690), .A2(new_n691), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n693), .A2(new_n812), .A3(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  NAND2_X1  g0633(.A1(new_n332), .A2(new_n686), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n330), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n335), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n642), .A2(new_n700), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n679), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(new_n840), .B2(new_n700), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n679), .A2(new_n686), .A3(new_n838), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(new_n748), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n812), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n773), .A2(G303), .B1(G283), .B2(new_n778), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n219), .B2(new_n765), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT97), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n784), .A2(G87), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n787), .A2(G294), .B1(G311), .B2(new_n761), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n757), .A2(new_n512), .ZN(new_n852));
  NOR4_X1   g0652(.A1(new_n851), .A2(new_n274), .A3(new_n790), .A4(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n773), .A2(G137), .B1(G150), .B2(new_n778), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n800), .B2(new_n765), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G143), .B2(new_n787), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT34), .ZN(new_n857));
  INV_X1    g0657(.A(new_n752), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n418), .B1(G58), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n784), .A2(G68), .B1(new_n758), .B2(G50), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n760), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n807), .B1(new_n853), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n807), .A2(new_n821), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT96), .Z(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n319), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n838), .A2(new_n821), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n864), .A2(new_n813), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n845), .A2(new_n870), .ZN(G384));
  XNOR2_X1  g0671(.A(new_n684), .B(KEYINPUT99), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n640), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n371), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n686), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n641), .B(new_n875), .C1(new_n357), .C2(new_n371), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT14), .B1(new_n373), .B2(new_n300), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n373), .A2(G179), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n353), .A2(new_n337), .A3(G169), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n874), .B(new_n686), .C1(new_n880), .C2(new_n378), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n840), .A2(new_n700), .A3(new_n839), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n883), .B1(new_n884), .B2(new_n837), .ZN(new_n885));
  INV_X1    g0685(.A(new_n684), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n422), .B1(KEYINPUT16), .B2(new_n421), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n452), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n886), .B(new_n888), .C1(new_n466), .C2(new_n443), .ZN(new_n889));
  INV_X1    g0689(.A(new_n439), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n635), .A2(new_n886), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n452), .B2(new_n887), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT37), .B1(new_n451), .B2(new_n463), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n463), .A2(new_n872), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n439), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n889), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n889), .A2(KEYINPUT38), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n873), .B1(new_n885), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n895), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n401), .A2(new_n438), .A3(KEYINPUT17), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT17), .B1(new_n401), .B2(new_n438), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT101), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT101), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n441), .A2(new_n908), .A3(new_n442), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n909), .A3(new_n640), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n439), .A2(KEYINPUT100), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT100), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n401), .A2(new_n438), .A3(new_n912), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n911), .A2(new_n636), .A3(new_n895), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT37), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n904), .A2(new_n910), .B1(new_n915), .B2(new_n896), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n901), .B1(new_n916), .B2(KEYINPUT38), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n372), .A2(new_n700), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n900), .A2(KEYINPUT39), .A3(new_n901), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n903), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n468), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n711), .B2(new_n717), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n646), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n924), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n882), .A2(new_n839), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n929), .B1(new_n743), .B2(new_n930), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n889), .A2(KEYINPUT38), .A3(new_n897), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT38), .B1(new_n889), .B2(new_n897), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n838), .B1(new_n876), .B2(new_n881), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n673), .A2(new_n671), .A3(new_n688), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n676), .A2(new_n937), .A3(new_n511), .A4(new_n700), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n938), .A2(KEYINPUT31), .B1(new_n739), .B2(new_n686), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n940));
  OAI211_X1 g0740(.A(KEYINPUT40), .B(new_n936), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n934), .A2(new_n935), .B1(new_n917), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n939), .A2(new_n940), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n468), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n943), .B(new_n945), .Z(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(G330), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n928), .B(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n203), .B2(new_n810), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n517), .B(KEYINPUT98), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n219), .B1(new_n950), .B2(KEYINPUT35), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n951), .B(new_n229), .C1(KEYINPUT35), .C2(new_n950), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT36), .ZN(new_n953));
  OAI21_X1  g0753(.A(G77), .B1(new_n230), .B2(new_n231), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n233), .A2(new_n954), .B1(G50), .B2(new_n231), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(G1), .A3(new_n809), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n949), .A2(new_n953), .A3(new_n956), .ZN(G367));
  NAND2_X1  g0757(.A1(new_n525), .A2(new_n686), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n676), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n551), .B2(new_n700), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n702), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT42), .Z(new_n962));
  OAI21_X1  g0762(.A(new_n551), .B1(new_n959), .B2(new_n629), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n700), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n660), .A2(new_n700), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n966), .A2(new_n509), .A3(new_n652), .A4(new_n657), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n662), .B2(new_n966), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n965), .A2(KEYINPUT43), .A3(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n968), .B(KEYINPUT43), .Z(new_n970));
  NAND2_X1  g0770(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(KEYINPUT102), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT102), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n965), .A2(new_n973), .A3(new_n970), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n969), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n698), .A2(new_n960), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n975), .B(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n707), .B(KEYINPUT41), .Z(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n697), .B(new_n701), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(new_n692), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n749), .A2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT104), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n703), .A2(new_n960), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(KEYINPUT103), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT103), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n703), .A2(new_n987), .A3(new_n960), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n703), .A2(new_n960), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT44), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n986), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n698), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n983), .A2(KEYINPUT104), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n991), .A2(new_n993), .A3(new_n699), .A4(new_n994), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n984), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n980), .B1(new_n999), .B2(new_n749), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n811), .A2(G1), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n978), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(G317), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n418), .B1(new_n1003), .B2(new_n760), .C1(new_n475), .C2(new_n785), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT106), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n782), .B2(new_n765), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1004), .A2(KEYINPUT106), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT105), .B1(new_n757), .B2(new_n219), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT46), .ZN(new_n1009));
  INV_X1    g0809(.A(G303), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n772), .A2(new_n763), .B1(new_n1010), .B2(new_n788), .ZN(new_n1011));
  NOR4_X1   g0811(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n778), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1012), .B1(new_n753), .B2(new_n1013), .C1(new_n481), .C2(new_n752), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n273), .B1(new_n795), .B2(G50), .ZN(new_n1015));
  INV_X1    g0815(.A(G137), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1015), .B1(new_n1016), .B2(new_n760), .C1(new_n800), .C2(new_n1013), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G150), .B2(new_n787), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n230), .B2(new_n757), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G143), .B2(new_n773), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n231), .B2(new_n752), .C1(new_n319), .C2(new_n785), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1014), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT47), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n807), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n968), .A2(new_n822), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n815), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n824), .B1(new_n207), .B2(new_n324), .C1(new_n1026), .C2(new_n242), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1024), .A2(new_n813), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1002), .A2(new_n1028), .ZN(G387));
  NAND2_X1  g0829(.A1(new_n984), .A2(new_n997), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n707), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n749), .A2(new_n982), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n265), .A2(new_n778), .B1(new_n795), .B2(G68), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n258), .B2(new_n760), .C1(new_n324), .C2(new_n752), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G77), .B2(new_n758), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n787), .A2(G50), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n773), .A2(G159), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n418), .B1(G97), .B2(new_n784), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n773), .A2(G322), .B1(G311), .B2(new_n778), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n1010), .B2(new_n765), .C1(new_n1003), .C2(new_n788), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT48), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n782), .B2(new_n752), .C1(new_n753), .C2(new_n757), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT49), .Z(new_n1045));
  NAND2_X1  g0845(.A1(new_n761), .A2(G326), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n418), .B(new_n1046), .C1(new_n219), .C2(new_n785), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1040), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n812), .B1(new_n1048), .B2(new_n807), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n697), .A2(new_n823), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n231), .A2(new_n319), .ZN(new_n1052));
  OAI21_X1  g0852(.A(KEYINPUT50), .B1(new_n264), .B2(G50), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT50), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n265), .A2(new_n1054), .A3(new_n211), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n706), .A2(new_n283), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n815), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT107), .Z(new_n1058));
  INV_X1    g0858(.A(new_n239), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1058), .B1(new_n283), .B2(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(G107), .B2(new_n207), .C1(new_n706), .C2(new_n819), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n824), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1051), .A2(new_n1062), .B1(new_n1001), .B2(new_n982), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1033), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(KEYINPUT108), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT108), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1033), .A2(new_n1066), .A3(new_n1063), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1067), .ZN(G393));
  OAI21_X1  g0868(.A(new_n824), .B1(new_n207), .B2(new_n475), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n815), .B2(new_n246), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n785), .A2(new_n217), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n418), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n772), .A2(new_n258), .B1(new_n800), .B2(new_n788), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT51), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1071), .B(new_n1075), .C1(new_n1074), .C2(new_n1073), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n795), .A2(new_n265), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n761), .A2(G143), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n757), .A2(new_n231), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n752), .A2(new_n319), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(G50), .C2(new_n778), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n772), .A2(new_n1003), .B1(new_n763), .B2(new_n788), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT52), .Z(new_n1084));
  AOI211_X1 g0884(.A(new_n274), .B(new_n1084), .C1(G116), .C2(new_n858), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n795), .A2(G294), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n778), .A2(G303), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n784), .A2(G107), .B1(new_n758), .B2(G283), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n760), .A2(new_n786), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1082), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1070), .B1(new_n1091), .B2(new_n807), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1092), .B(new_n813), .C1(new_n822), .C2(new_n960), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n996), .A2(new_n998), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1001), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n707), .B1(new_n1030), .B2(new_n1094), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n999), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(G390));
  NAND2_X1  g0899(.A1(new_n919), .A2(new_n922), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n837), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n882), .B1(new_n842), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n920), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n716), .A2(new_n700), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1101), .B1(new_n1105), .B2(new_n836), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n917), .B(new_n920), .C1(new_n1106), .C2(new_n883), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n747), .A2(G330), .A3(new_n839), .A4(new_n882), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1104), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n944), .A2(new_n691), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n936), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n919), .A2(new_n922), .B1(new_n1102), .B2(new_n920), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1107), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(G330), .B1(new_n939), .B2(new_n940), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n883), .B1(new_n1117), .B2(new_n838), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1108), .A2(new_n1118), .A3(new_n1106), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n746), .A2(new_n700), .ZN(new_n1120));
  OAI211_X1 g0920(.A(G330), .B(new_n839), .C1(new_n939), .C2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1111), .A2(new_n936), .B1(new_n1121), .B2(new_n883), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n842), .A2(new_n1101), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1119), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n925), .B(G330), .C1(new_n939), .C2(new_n940), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1125), .A2(new_n926), .A3(new_n646), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT109), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1125), .A2(new_n926), .A3(new_n646), .A4(KEYINPUT109), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1124), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1116), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1110), .A3(new_n1115), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n1031), .A3(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n785), .A2(new_n231), .B1(new_n760), .B2(new_n753), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n793), .B(new_n1135), .C1(new_n309), .C2(new_n778), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n274), .B(new_n1080), .C1(new_n479), .C2(new_n795), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n787), .A2(G116), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n773), .A2(G283), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(G128), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n772), .A2(new_n1141), .B1(new_n861), .B2(new_n788), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT110), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n758), .A2(G150), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n273), .B1(new_n1144), .B2(KEYINPUT53), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n784), .A2(G50), .B1(new_n761), .B2(G125), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n800), .C2(new_n752), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT54), .B(G143), .Z(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1148), .B1(new_n1016), .B2(new_n1013), .C1(new_n765), .C2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1144), .A2(KEYINPUT53), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1140), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1153), .A2(new_n807), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n812), .B(new_n1154), .C1(new_n1100), .C2(new_n821), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n867), .A2(new_n264), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1116), .A2(new_n1001), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1134), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT111), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1134), .A2(KEYINPUT111), .A3(new_n1157), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(G378));
  NAND2_X1  g0962(.A1(new_n934), .A2(new_n935), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n299), .A2(new_n302), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  XOR2_X1   g0965(.A(new_n1164), .B(new_n1165), .Z(new_n1166));
  AND2_X1   g0966(.A1(new_n267), .A2(new_n886), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1166), .B(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n910), .A2(new_n904), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n915), .A2(new_n896), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT38), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g0971(.A(KEYINPUT40), .B(new_n931), .C1(new_n1171), .C2(new_n932), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1163), .A2(new_n1168), .A3(G330), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1168), .B1(new_n943), .B2(G330), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n924), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n901), .B2(new_n900), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1172), .B(G330), .C1(new_n1178), .C2(KEYINPUT40), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1168), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n903), .A2(new_n923), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n1182), .A3(new_n1173), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT114), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1183), .A2(KEYINPUT113), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n1183), .B2(KEYINPUT113), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1176), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1183), .A2(KEYINPUT113), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT114), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1176), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1183), .A2(KEYINPUT113), .A3(new_n1184), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1187), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1116), .B2(new_n1124), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n707), .A2(KEYINPUT57), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1095), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1168), .A2(new_n821), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n867), .A2(new_n211), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1013), .A2(new_n861), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n752), .A2(new_n258), .B1(new_n765), .B2(new_n1016), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n773), .C2(G125), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n1141), .B2(new_n788), .C1(new_n757), .C2(new_n1150), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT59), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n800), .B2(new_n785), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G41), .B1(new_n1072), .B2(G33), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n1205), .A2(new_n1207), .B1(G50), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n784), .A2(G58), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT112), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G107), .A2(new_n787), .B1(new_n858), .B2(G68), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n782), .C2(new_n760), .ZN(new_n1213));
  AOI21_X1  g1013(.A(G41), .B1(new_n795), .B2(new_n323), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n319), .B2(new_n757), .C1(new_n222), .C2(new_n1013), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n772), .A2(new_n219), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1213), .A2(new_n1072), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT58), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n807), .B1(new_n1209), .B2(new_n1218), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1199), .A2(new_n813), .A3(new_n1200), .A4(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1176), .A2(KEYINPUT115), .A3(new_n1183), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT115), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n924), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(KEYINPUT57), .B(new_n1031), .C1(new_n1224), .C2(new_n1195), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1198), .A2(new_n1220), .A3(new_n1225), .ZN(G375));
  XOR2_X1   g1026(.A(new_n1001), .B(KEYINPUT116), .Z(new_n1227));
  NAND2_X1  g1027(.A1(new_n883), .A2(new_n821), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1013), .A2(new_n219), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n274), .B1(new_n761), .B2(G303), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n222), .B2(new_n757), .C1(new_n785), .C2(new_n319), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1229), .B(new_n1231), .C1(G294), .C2(new_n773), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n788), .A2(new_n782), .B1(new_n324), .B2(new_n752), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT117), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1232), .B(new_n1234), .C1(new_n481), .C2(new_n765), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1211), .B1(new_n258), .B2(new_n765), .C1(new_n1013), .C2(new_n1150), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G132), .B2(new_n773), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n787), .A2(G137), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n757), .A2(new_n800), .B1(new_n760), .B2(new_n1141), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT118), .Z(new_n1240));
  NAND4_X1  g1040(.A1(new_n1237), .A2(new_n1072), .A3(new_n1238), .A4(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n752), .A2(new_n211), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1235), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n812), .B1(new_n1243), .B2(new_n807), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(G68), .B2(new_n866), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT119), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1124), .A2(new_n1227), .B1(new_n1228), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1124), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1248), .A2(new_n980), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1249), .B2(new_n1131), .ZN(G381));
  AND3_X1   g1050(.A1(new_n1002), .A2(new_n1098), .A3(new_n1028), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1065), .A2(new_n832), .A3(new_n1067), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(new_n1252), .A2(G384), .A3(G381), .A4(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(G375), .A2(new_n1158), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(G407));
  OAI21_X1  g1056(.A(new_n1255), .B1(new_n1254), .B2(new_n685), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(G213), .ZN(G409));
  INV_X1    g1058(.A(new_n1158), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1221), .A2(new_n1223), .A3(new_n1227), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1220), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT120), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT120), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1260), .A2(new_n1263), .A3(new_n1220), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n980), .B(new_n1195), .C1(new_n1187), .C2(new_n1192), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1259), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(G378), .A2(new_n1198), .A3(new_n1220), .A4(new_n1225), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(G213), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(G343), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT122), .ZN(new_n1273));
  INV_X1    g1073(.A(G384), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT121), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1124), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT60), .B1(new_n1276), .B2(new_n1194), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1275), .B1(new_n1277), .B2(new_n1131), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n707), .B1(new_n1248), .B2(KEYINPUT60), .ZN(new_n1279));
  OAI211_X1 g1079(.A(KEYINPUT121), .B(new_n1130), .C1(new_n1248), .C2(KEYINPUT60), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1273), .B(new_n1274), .C1(new_n1281), .C2(new_n1247), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1274), .A2(new_n1273), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1281), .A2(new_n1247), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1282), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1269), .A2(KEYINPUT63), .A3(new_n1272), .A4(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT124), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1065), .A2(new_n832), .A3(new_n1067), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n832), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G393), .A2(G396), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(KEYINPUT124), .A3(new_n1253), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G387), .A2(G390), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1294), .A2(new_n1296), .A3(new_n1252), .A4(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G387), .A2(KEYINPUT125), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(G390), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1295), .A2(new_n1253), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(G387), .A2(KEYINPUT125), .A3(new_n1098), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1298), .A2(new_n1303), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1289), .A2(new_n1290), .A3(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1269), .A2(new_n1272), .A3(new_n1288), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1271), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1281), .A2(new_n1247), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(KEYINPUT122), .A3(G384), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1271), .A2(G2897), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1311), .A2(new_n1285), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1312), .B1(new_n1311), .B2(new_n1285), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(KEYINPUT123), .B1(new_n1309), .B2(new_n1315), .ZN(new_n1316));
  OR3_X1    g1116(.A1(new_n1309), .A2(new_n1315), .A3(KEYINPUT123), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1305), .A2(new_n1308), .A3(new_n1316), .A4(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1304), .ZN(new_n1319));
  AOI211_X1 g1119(.A(new_n1271), .B(new_n1287), .C1(new_n1267), .C2(new_n1268), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1290), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1323));
  OAI22_X1  g1123(.A1(new_n1306), .A2(new_n1323), .B1(new_n1309), .B2(new_n1315), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1319), .B1(new_n1322), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1318), .A2(new_n1325), .ZN(G405));
  NAND2_X1  g1126(.A1(G375), .A2(new_n1259), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1268), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1327), .A2(KEYINPUT127), .A3(new_n1268), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1287), .A3(new_n1331), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1288), .A2(new_n1327), .A3(KEYINPUT127), .A4(new_n1268), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1304), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1332), .A2(new_n1333), .A3(new_n1319), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(G402));
endmodule


