//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n203));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G169gat), .B2(G176gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n209), .B(KEYINPUT24), .Z(new_n210));
  NOR2_X1   g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n208), .B(KEYINPUT25), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n209), .B(KEYINPUT24), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n207), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n212), .B1(new_n215), .B2(KEYINPUT25), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT27), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n217), .A2(KEYINPUT27), .ZN(new_n220));
  NOR3_X1   g019(.A1(new_n220), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n219), .A2(new_n221), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT26), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n202), .A2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(KEYINPUT67), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(KEYINPUT67), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n204), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT28), .ZN(new_n230));
  INV_X1    g029(.A(new_n220), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(new_n218), .A3(KEYINPUT66), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n217), .A2(KEYINPUT27), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(new_n220), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G190gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n230), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n216), .B1(new_n229), .B2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(G127gat), .B(G134gat), .Z(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241));
  OR3_X1    g040(.A1(new_n240), .A2(KEYINPUT1), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n240), .B1(KEYINPUT1), .B2(new_n241), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n238), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(new_n228), .A3(new_n222), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n241), .A2(KEYINPUT1), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(new_n240), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n249), .A3(new_n216), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G227gat), .A2(G233gat), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n253));
  XNOR2_X1  g052(.A(G15gat), .B(G43gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(G71gat), .B(G99gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n245), .A2(new_n250), .A3(new_n252), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n252), .B1(new_n245), .B2(new_n250), .ZN(new_n260));
  INV_X1    g059(.A(new_n253), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n259), .B(new_n256), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT34), .ZN(new_n263));
  OAI211_X1 g062(.A(KEYINPUT32), .B(new_n263), .C1(new_n251), .C2(new_n252), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT32), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT34), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n258), .A2(new_n262), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT36), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n264), .A2(new_n262), .A3(new_n258), .A4(new_n266), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n268), .A2(new_n269), .A3(new_n270), .A4(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n270), .ZN(new_n273));
  NAND2_X1  g072(.A1(KEYINPUT69), .A2(KEYINPUT36), .ZN(new_n274));
  INV_X1    g073(.A(new_n271), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n273), .B(new_n274), .C1(new_n275), .C2(new_n267), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT82), .ZN(new_n279));
  NAND2_X1  g078(.A1(G228gat), .A2(G233gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT80), .ZN(new_n281));
  XNOR2_X1  g080(.A(G197gat), .B(G204gat), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n283), .A2(KEYINPUT70), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(KEYINPUT70), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G211gat), .B(G218gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G155gat), .B(G162gat), .ZN(new_n290));
  XOR2_X1   g089(.A(G141gat), .B(G148gat), .Z(new_n291));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT2), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT3), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n291), .B(new_n296), .C1(new_n292), .C2(new_n290), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n289), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n299), .B1(new_n288), .B2(KEYINPUT29), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n298), .A2(new_n300), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n281), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n280), .B1(new_n306), .B2(new_n307), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT81), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n305), .B2(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n301), .A2(new_n302), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n301), .A2(new_n302), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT29), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n315), .A2(KEYINPUT81), .A3(new_n289), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n309), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n279), .B1(new_n317), .B2(G22gat), .ZN(new_n318));
  XOR2_X1   g117(.A(G78gat), .B(G106gat), .Z(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT31), .B(G50gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n317), .A2(G22gat), .ZN(new_n323));
  INV_X1    g122(.A(G22gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n311), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT81), .B1(new_n315), .B2(new_n289), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n310), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n324), .B1(new_n327), .B2(new_n309), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n318), .A2(new_n322), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n328), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(new_n324), .A3(new_n309), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n330), .A2(new_n279), .A3(new_n331), .A4(new_n321), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G57gat), .B(G85gat), .Z(new_n334));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n249), .A2(new_n300), .A3(new_n298), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n307), .A2(new_n244), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342));
  OAI211_X1 g141(.A(KEYINPUT77), .B(KEYINPUT5), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n342), .B1(new_n339), .B2(new_n340), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT5), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n249), .B1(new_n307), .B2(KEYINPUT3), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n303), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n303), .A2(KEYINPUT75), .A3(new_n349), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n342), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(new_n339), .B2(KEYINPUT4), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n339), .A2(KEYINPUT4), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n339), .A2(new_n356), .A3(KEYINPUT4), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n355), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n348), .B1(new_n354), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n339), .B(KEYINPUT4), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n355), .A2(KEYINPUT5), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n303), .A2(KEYINPUT75), .A3(new_n349), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT75), .B1(new_n303), .B2(new_n349), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n363), .B(new_n364), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n338), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n361), .B1(new_n366), .B2(new_n365), .ZN(new_n370));
  INV_X1    g169(.A(new_n348), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n338), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n367), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n369), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n338), .B(new_n375), .C1(new_n362), .C2(new_n368), .ZN(new_n378));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(new_n239), .B2(new_n304), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n379), .B1(new_n247), .B2(new_n216), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n288), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT71), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n381), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n239), .A2(new_n380), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(KEYINPUT72), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT72), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n389), .B1(new_n239), .B2(new_n380), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n386), .B(new_n289), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(KEYINPUT71), .B(new_n288), .C1(new_n381), .C2(new_n382), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n385), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n396), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n385), .A2(new_n391), .A3(new_n392), .A4(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(KEYINPUT30), .A3(new_n399), .ZN(new_n400));
  OR3_X1    g199(.A1(new_n393), .A2(KEYINPUT30), .A3(new_n396), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n377), .A2(new_n378), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n278), .B1(new_n333), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT84), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT39), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n341), .B2(new_n342), .ZN(new_n406));
  INV_X1    g205(.A(new_n363), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n407), .B1(new_n352), .B2(new_n353), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n408), .B2(new_n342), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(new_n405), .A3(new_n355), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n409), .A2(KEYINPUT40), .A3(new_n373), .A4(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n412), .A2(new_n369), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(new_n373), .A3(new_n411), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT40), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n413), .A2(new_n401), .A3(new_n400), .A4(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n399), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT37), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n385), .A2(new_n391), .A3(new_n419), .A4(new_n392), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n420), .A2(new_n396), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n247), .B2(new_n216), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n289), .B(new_n387), .C1(new_n422), .C2(new_n380), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n386), .A2(KEYINPUT83), .A3(new_n289), .A4(new_n387), .ZN(new_n426));
  INV_X1    g225(.A(new_n390), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n382), .A2(new_n389), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n381), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n425), .B(new_n426), .C1(new_n429), .C2(new_n289), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT38), .B1(new_n430), .B2(KEYINPUT37), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n418), .B1(new_n421), .B2(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n393), .A2(KEYINPUT37), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n420), .A2(new_n396), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT38), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n432), .A2(new_n435), .A3(new_n377), .A4(new_n378), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n436), .A3(new_n333), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n403), .B1(new_n404), .B2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n417), .A2(new_n436), .A3(KEYINPUT84), .A4(new_n333), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n275), .A2(new_n267), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n329), .A2(new_n332), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT86), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT86), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n329), .A2(new_n332), .A3(new_n443), .A4(new_n440), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n402), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT35), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n377), .A2(new_n378), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT35), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n400), .A2(new_n401), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n447), .B1(new_n451), .B2(new_n441), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n329), .A2(new_n332), .A3(new_n440), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n453), .A2(KEYINPUT85), .A3(new_n449), .A4(new_n402), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n438), .A2(new_n439), .B1(new_n446), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G43gat), .B(G50gat), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT15), .ZN(new_n458));
  INV_X1    g257(.A(G29gat), .ZN(new_n459));
  INV_X1    g258(.A(G36gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT14), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(new_n459), .A3(new_n460), .ZN(new_n464));
  AOI211_X1 g263(.A(new_n458), .B(new_n461), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n464), .A2(new_n462), .B1(G29gat), .B2(G36gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(KEYINPUT15), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n457), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(KEYINPUT15), .ZN(new_n469));
  INV_X1    g268(.A(new_n457), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT17), .ZN(new_n473));
  XNOR2_X1  g272(.A(G15gat), .B(G22gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(G1gat), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n476));
  OAI21_X1  g275(.A(G8gat), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT16), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n474), .B1(new_n478), .B2(G1gat), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(G1gat), .B2(new_n474), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n477), .B(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT17), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n468), .A2(new_n482), .A3(new_n471), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n473), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT88), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n477), .B(new_n480), .Z(new_n488));
  INV_X1    g287(.A(new_n472), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT18), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n484), .A2(KEYINPUT18), .A3(new_n490), .A4(new_n487), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n481), .A2(new_n472), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n486), .B(new_n497), .Z(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G113gat), .B(G141gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(G197gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT11), .B(G169gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n504), .B(KEYINPUT12), .Z(new_n505));
  NAND4_X1  g304(.A1(new_n493), .A2(new_n494), .A3(new_n500), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT90), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n491), .A2(new_n492), .B1(new_n496), .B2(new_n499), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT90), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(new_n494), .A4(new_n505), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n494), .ZN(new_n512));
  INV_X1    g311(.A(new_n505), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G57gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(G64gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(G64gat), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(KEYINPUT94), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(KEYINPUT94), .B2(new_n519), .ZN(new_n521));
  INV_X1    g320(.A(G71gat), .ZN(new_n522));
  INV_X1    g321(.A(G78gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT9), .ZN(new_n524));
  NAND2_X1  g323(.A1(G71gat), .A2(G78gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G64gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(G57gat), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT92), .B1(new_n529), .B2(new_n518), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(G57gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n519), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT9), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n525), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n530), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n537));
  OR3_X1    g336(.A1(KEYINPUT91), .A2(G71gat), .A3(G78gat), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT91), .B1(G71gat), .B2(G78gat), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n538), .A2(new_n539), .B1(G71gat), .B2(G78gat), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n537), .B1(new_n536), .B2(new_n540), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n527), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n488), .B1(new_n544), .B2(KEYINPUT21), .ZN(new_n545));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n545), .B(new_n546), .Z(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G127gat), .B(G155gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(G183gat), .ZN(new_n554));
  INV_X1    g353(.A(G211gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n551), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT101), .B(G85gat), .ZN(new_n560));
  INV_X1    g359(.A(G92gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n560), .A2(new_n561), .B1(KEYINPUT8), .B2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G99gat), .B(G106gat), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AND3_X1   g364(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n566));
  OR2_X1    g365(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n567));
  NAND2_X1  g366(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n570));
  AND2_X1   g369(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n571));
  NOR2_X1   g370(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n563), .A2(new_n565), .A3(new_n569), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n573), .ZN(new_n575));
  AND2_X1   g374(.A1(KEYINPUT101), .A2(G85gat), .ZN(new_n576));
  NOR2_X1   g375(.A1(KEYINPUT101), .A2(G85gat), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n561), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n562), .A2(KEYINPUT8), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n564), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n489), .A2(new_n582), .B1(KEYINPUT41), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n574), .A2(new_n581), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n473), .A2(new_n483), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G190gat), .B(G218gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT102), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n587), .B(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n583), .A2(KEYINPUT41), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT98), .ZN(new_n593));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n591), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n543), .A2(new_n585), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT10), .ZN(new_n598));
  XNOR2_X1  g397(.A(G57gat), .B(G64gat), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n535), .B1(new_n599), .B2(new_n532), .ZN(new_n600));
  INV_X1    g399(.A(new_n533), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n540), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT93), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(new_n527), .A3(new_n582), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n597), .A2(new_n598), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n544), .A2(KEYINPUT10), .A3(new_n582), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT103), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n612));
  INV_X1    g411(.A(new_n610), .ZN(new_n613));
  AOI211_X1 g412(.A(new_n612), .B(new_n613), .C1(new_n607), .C2(new_n608), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n606), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n613), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n609), .A2(new_n610), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n617), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n559), .A2(new_n596), .A3(new_n627), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n456), .A2(new_n516), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n448), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G1gat), .ZN(G1324gat));
  INV_X1    g431(.A(new_n450), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G8gat), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT42), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n478), .A2(new_n635), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  MUX2_X1   g438(.A(KEYINPUT42), .B(new_n636), .S(new_n639), .Z(G1325gat));
  AOI21_X1  g439(.A(G15gat), .B1(new_n629), .B2(new_n440), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n277), .A2(G15gat), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n629), .B2(new_n642), .ZN(G1326gat));
  NAND2_X1  g442(.A1(new_n329), .A2(new_n332), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT43), .B(G22gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1327gat));
  XOR2_X1   g446(.A(new_n551), .B(new_n558), .Z(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n627), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n515), .A2(KEYINPUT105), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT105), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n511), .A2(new_n652), .A3(new_n514), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n446), .A2(new_n455), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n437), .A2(new_n404), .ZN(new_n657));
  INV_X1    g456(.A(new_n402), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n277), .B1(new_n658), .B2(new_n644), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n439), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662));
  INV_X1    g461(.A(new_n596), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT107), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n596), .B1(new_n656), .B2(new_n660), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n667), .A3(new_n662), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT106), .B1(new_n666), .B2(new_n662), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n671), .B(KEYINPUT44), .C1(new_n456), .C2(new_n596), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n655), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G29gat), .B1(new_n675), .B2(new_n448), .ZN(new_n676));
  NOR4_X1   g475(.A1(new_n456), .A2(new_n516), .A3(new_n596), .A4(new_n649), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n459), .A3(new_n630), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n676), .A2(new_n680), .ZN(G1328gat));
  OAI21_X1  g480(.A(G36gat), .B1(new_n675), .B2(new_n450), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n677), .A2(new_n460), .A3(new_n633), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(KEYINPUT46), .Z(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(G1329gat));
  INV_X1    g484(.A(G43gat), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n677), .A2(new_n686), .A3(new_n440), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI211_X1 g488(.A(new_n278), .B(new_n655), .C1(new_n669), .C2(new_n673), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691));
  OAI21_X1  g490(.A(G43gat), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n674), .A2(new_n691), .A3(new_n277), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n690), .A2(new_n686), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n688), .B1(new_n695), .B2(new_n687), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(G1330gat));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n674), .A2(new_n644), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G50gat), .ZN(new_n700));
  INV_X1    g499(.A(G50gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n677), .A2(new_n701), .A3(new_n644), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n698), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n702), .ZN(new_n704));
  AOI211_X1 g503(.A(KEYINPUT48), .B(new_n704), .C1(new_n699), .C2(G50gat), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(G1331gat));
  NOR4_X1   g505(.A1(new_n648), .A2(new_n663), .A3(new_n627), .A4(new_n654), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n448), .B(KEYINPUT109), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n661), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n661), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT110), .Z(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n450), .ZN(new_n713));
  NOR2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  AND2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n713), .B2(new_n714), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n712), .B2(new_n278), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n707), .A2(new_n661), .A3(new_n522), .A4(new_n440), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1334gat));
  NOR2_X1   g521(.A1(new_n712), .A2(new_n333), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(new_n523), .ZN(G1335gat));
  NOR2_X1   g523(.A1(new_n559), .A2(new_n654), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n666), .A2(KEYINPUT51), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT51), .B1(new_n666), .B2(new_n725), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(new_n626), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n630), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n725), .A2(new_n626), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n669), .B2(new_n673), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n448), .A2(new_n560), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n730), .A2(new_n560), .B1(new_n732), .B2(new_n733), .ZN(G1336gat));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n450), .B(new_n731), .C1(new_n669), .C2(new_n673), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(new_n561), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n728), .A2(new_n561), .A3(new_n633), .A4(new_n626), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n736), .B2(new_n561), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n739), .A3(KEYINPUT52), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741));
  OAI221_X1 g540(.A(new_n738), .B1(new_n735), .B2(new_n741), .C1(new_n736), .C2(new_n561), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1337gat));
  AOI21_X1  g542(.A(G99gat), .B1(new_n729), .B2(new_n440), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n277), .A2(G99gat), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n732), .B2(new_n745), .ZN(G1338gat));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(KEYINPUT53), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n644), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G106gat), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n333), .A2(G106gat), .A3(new_n627), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(KEYINPUT112), .Z(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n726), .B2(new_n727), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(KEYINPUT113), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n749), .B1(new_n751), .B2(new_n757), .ZN(new_n758));
  AOI211_X1 g557(.A(new_n748), .B(new_n756), .C1(new_n750), .C2(G106gat), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(G1339gat));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n611), .B2(new_n614), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n607), .A2(new_n613), .A3(new_n608), .ZN(new_n764));
  AND4_X1   g563(.A1(new_n763), .A2(new_n623), .A3(KEYINPUT54), .A4(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n761), .B1(new_n609), .B2(new_n610), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n763), .B1(new_n766), .B2(new_n764), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n621), .B(new_n762), .C1(new_n765), .C2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n625), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT115), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n772), .B(new_n625), .C1(new_n768), .C2(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n768), .A2(new_n769), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n771), .A2(new_n654), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n484), .A2(new_n490), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n486), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n490), .A2(new_n495), .A3(new_n498), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n504), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n507), .B2(new_n510), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n626), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n663), .B1(new_n775), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n780), .A2(KEYINPUT116), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784));
  AOI211_X1 g583(.A(new_n784), .B(new_n779), .C1(new_n507), .C2(new_n510), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n783), .A2(new_n785), .A3(new_n596), .ZN(new_n786));
  AND4_X1   g585(.A1(new_n773), .A2(new_n786), .A3(new_n771), .A4(new_n774), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n648), .B1(new_n782), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n654), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n559), .A2(new_n596), .A3(new_n627), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(new_n708), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n442), .A2(new_n444), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(new_n450), .ZN(new_n795));
  INV_X1    g594(.A(G113gat), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n796), .A3(new_n654), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n441), .B1(new_n788), .B2(new_n790), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n633), .A2(new_n448), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G113gat), .B1(new_n800), .B2(new_n516), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n801), .ZN(G1340gat));
  INV_X1    g601(.A(G120gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n795), .A2(new_n803), .A3(new_n626), .ZN(new_n804));
  OAI21_X1  g603(.A(G120gat), .B1(new_n800), .B2(new_n627), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1341gat));
  INV_X1    g605(.A(G127gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n800), .A2(new_n807), .A3(new_n648), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n795), .A2(new_n559), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n807), .ZN(G1342gat));
  INV_X1    g609(.A(G134gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n450), .A2(new_n663), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT117), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n794), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n815), .A2(KEYINPUT56), .ZN(new_n816));
  OAI21_X1  g615(.A(G134gat), .B1(new_n800), .B2(new_n596), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(KEYINPUT56), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(G1343gat));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n799), .A2(new_n278), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n333), .B1(new_n788), .B2(new_n790), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(KEYINPUT57), .ZN(new_n825));
  INV_X1    g624(.A(new_n768), .ZN(new_n826));
  XOR2_X1   g625(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n827));
  OAI21_X1  g626(.A(new_n515), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n828), .A2(new_n770), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n663), .B1(new_n829), .B2(new_n781), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n648), .B1(new_n830), .B2(new_n787), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n790), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(KEYINPUT57), .A3(new_n644), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n825), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n824), .A2(new_n823), .A3(KEYINPUT57), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n515), .B(new_n822), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G141gat), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n333), .A2(new_n277), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n516), .A2(G141gat), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n792), .A2(new_n450), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n820), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  AOI211_X1 g643(.A(KEYINPUT120), .B(new_n842), .C1(new_n836), .C2(G141gat), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n654), .B(new_n822), .C1(new_n834), .C2(new_n835), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n792), .A2(new_n838), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n633), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n846), .A2(G141gat), .B1(new_n848), .B2(new_n839), .ZN(new_n849));
  OAI22_X1  g648(.A1(new_n844), .A2(new_n845), .B1(new_n841), .B2(new_n849), .ZN(G1344gat));
  INV_X1    g649(.A(G148gat), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(new_n851), .A3(new_n626), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n822), .B1(new_n834), .B2(new_n835), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n627), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(KEYINPUT59), .A3(new_n851), .ZN(new_n855));
  INV_X1    g654(.A(new_n824), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n559), .A2(new_n516), .A3(new_n596), .A4(new_n627), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n831), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n333), .A2(KEYINPUT57), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n856), .A2(KEYINPUT57), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n626), .ZN(new_n861));
  OAI21_X1  g660(.A(G148gat), .B1(new_n861), .B2(new_n821), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n862), .A2(KEYINPUT59), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n852), .B1(new_n855), .B2(new_n863), .ZN(G1345gat));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n559), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n294), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n648), .A2(new_n294), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n822), .B(new_n867), .C1(new_n834), .C2(new_n835), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n866), .A2(new_n871), .A3(new_n868), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(G1346gat));
  OAI21_X1  g672(.A(G162gat), .B1(new_n853), .B2(new_n596), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n814), .A2(new_n295), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n847), .B2(new_n875), .ZN(G1347gat));
  AOI21_X1  g675(.A(new_n630), .B1(new_n788), .B2(new_n790), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n877), .A2(new_n633), .A3(new_n793), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT122), .ZN(new_n879));
  INV_X1    g678(.A(G169gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n880), .A3(new_n654), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n708), .A2(new_n450), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n798), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G169gat), .B1(new_n883), .B2(new_n516), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(G1348gat));
  INV_X1    g684(.A(G176gat), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n883), .A2(new_n886), .A3(new_n627), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n879), .A2(new_n626), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(new_n886), .ZN(G1349gat));
  NAND3_X1  g688(.A1(new_n878), .A2(new_n236), .A3(new_n559), .ZN(new_n890));
  OAI21_X1  g689(.A(G183gat), .B1(new_n883), .B2(new_n648), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g692(.A1(new_n879), .A2(new_n237), .A3(new_n663), .ZN(new_n894));
  OAI21_X1  g693(.A(G190gat), .B1(new_n883), .B2(new_n596), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT61), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1351gat));
  NOR3_X1   g696(.A1(new_n333), .A2(new_n277), .A3(new_n450), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n877), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(G197gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n654), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n901), .B(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n882), .A2(new_n278), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n860), .A2(new_n904), .A3(new_n515), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n858), .A2(new_n859), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n908), .B(new_n906), .C1(new_n909), .C2(new_n824), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT124), .B1(new_n910), .B2(new_n516), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n907), .A2(new_n911), .A3(G197gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n903), .A2(KEYINPUT125), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1352gat));
  INV_X1    g716(.A(G204gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n899), .A2(new_n918), .A3(new_n626), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT62), .Z(new_n920));
  OAI21_X1  g719(.A(G204gat), .B1(new_n861), .B2(new_n905), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1353gat));
  OAI211_X1 g721(.A(KEYINPUT63), .B(G211gat), .C1(new_n910), .C2(new_n648), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n923), .A2(KEYINPUT126), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(KEYINPUT126), .ZN(new_n925));
  INV_X1    g724(.A(new_n910), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n555), .B1(new_n926), .B2(new_n559), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n924), .B(new_n925), .C1(KEYINPUT63), .C2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n899), .A2(new_n555), .A3(new_n559), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1354gat));
  AND2_X1   g729(.A1(new_n899), .A2(new_n663), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n931), .A2(G218gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n663), .A2(G218gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n910), .B2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n932), .B(KEYINPUT127), .C1(new_n910), .C2(new_n933), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1355gat));
endmodule


