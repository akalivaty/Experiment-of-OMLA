//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n544,
    new_n546, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n561, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  AND3_X1   g038(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT68), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT68), .B1(new_n461), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n461), .A2(new_n463), .A3(new_n459), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  INV_X1    g045(.A(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n459), .A2(G2104), .ZN(new_n472));
  OAI22_X1  g047(.A1(new_n469), .A2(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  INV_X1    g049(.A(new_n469), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n461), .A2(new_n463), .A3(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(new_n459), .B2(G112), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n476), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  NOR3_X1   g058(.A1(new_n483), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n464), .B2(new_n465), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT71), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT4), .B1(new_n469), .B2(new_n483), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(new_n484), .C1(new_n464), .C2(new_n465), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n460), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI221_X1 g069(.A(new_n494), .B1(new_n493), .B2(new_n492), .C1(G102), .C2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n477), .A2(G126), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .A3(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n508), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n517));
  INV_X1    g092(.A(G51), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT74), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n517), .B(KEYINPUT73), .C1(new_n512), .C2(new_n518), .ZN(new_n525));
  INV_X1    g100(.A(new_n510), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT75), .B(G89), .Z(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n521), .A2(new_n524), .A3(new_n525), .A4(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n507), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n510), .A2(new_n533), .B1(new_n512), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  AOI22_X1  g111(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n507), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT76), .B(G43), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n510), .A2(new_n539), .B1(new_n512), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT77), .ZN(G188));
  INV_X1    g124(.A(G53), .ZN(new_n550));
  OR3_X1    g125(.A1(new_n512), .A2(KEYINPUT9), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT9), .B1(new_n512), .B2(new_n550), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n526), .A2(G91), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT78), .Z(new_n556));
  XNOR2_X1  g131(.A(KEYINPUT79), .B(G65), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n556), .B1(new_n505), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n553), .B(new_n554), .C1(new_n507), .C2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  NAND2_X1  g135(.A1(new_n526), .A2(G87), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n562));
  INV_X1    g137(.A(new_n512), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G49), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(G288));
  NAND2_X1  g140(.A1(new_n505), .A2(G61), .ZN(new_n566));
  NAND2_X1  g141(.A1(G73), .A2(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT80), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n507), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(KEYINPUT81), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n526), .A2(G86), .B1(new_n563), .B2(G48), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(KEYINPUT81), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G305));
  AOI22_X1  g148(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n574), .A2(new_n507), .ZN(new_n575));
  INV_X1    g150(.A(G47), .ZN(new_n576));
  INV_X1    g151(.A(G85), .ZN(new_n577));
  OAI221_X1 g152(.A(new_n575), .B1(new_n576), .B2(new_n512), .C1(new_n577), .C2(new_n510), .ZN(G290));
  NAND2_X1  g153(.A1(G301), .A2(G868), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G54), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n580), .A2(new_n507), .B1(new_n512), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT83), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT83), .ZN(new_n584));
  OAI221_X1 g159(.A(new_n584), .B1(new_n512), .B2(new_n581), .C1(new_n580), .C2(new_n507), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n505), .A2(G92), .A3(new_n509), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT82), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT82), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n505), .A2(new_n590), .A3(G92), .A4(new_n509), .ZN(new_n591));
  AOI21_X1  g166(.A(KEYINPUT10), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n589), .A2(KEYINPUT10), .A3(new_n591), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n579), .B1(new_n596), .B2(G868), .ZN(G321));
  XNOR2_X1  g172(.A(G321), .B(KEYINPUT84), .ZN(G284));
  NAND2_X1  g173(.A1(G286), .A2(G868), .ZN(new_n599));
  INV_X1    g174(.A(G299), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(G297));
  OAI21_X1  g176(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n596), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g183(.A1(new_n464), .A2(new_n465), .ZN(new_n609));
  INV_X1    g184(.A(new_n472), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT12), .Z(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  INV_X1    g188(.A(G2100), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n475), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n477), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(new_n459), .B2(G111), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT85), .ZN(new_n621));
  INV_X1    g196(.A(G2096), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n615), .A2(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT86), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  XOR2_X1   g205(.A(G2443), .B(G2446), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT87), .B(KEYINPUT16), .Z(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(G14), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2072), .B(G2078), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT88), .ZN(new_n643));
  XOR2_X1   g218(.A(G2067), .B(G2678), .Z(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(KEYINPUT17), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n645), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT89), .ZN(new_n649));
  INV_X1    g224(.A(new_n644), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n650), .A2(new_n641), .A3(new_n642), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT18), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n641), .A3(new_n644), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(new_n614), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT90), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(new_n622), .ZN(G227));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n659), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  AOI22_X1  g240(.A1(new_n663), .A2(KEYINPUT20), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n659), .A3(new_n662), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n666), .B(new_n668), .C1(KEYINPUT20), .C2(new_n663), .ZN(new_n669));
  XOR2_X1   g244(.A(G1991), .B(G1996), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G229));
  XNOR2_X1  g250(.A(KEYINPUT92), .B(G16), .ZN(new_n676));
  INV_X1    g251(.A(G24), .ZN(new_n677));
  OAI21_X1  g252(.A(KEYINPUT93), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OR3_X1    g253(.A1(new_n676), .A2(KEYINPUT93), .A3(new_n677), .ZN(new_n679));
  INV_X1    g254(.A(G290), .ZN(new_n680));
  INV_X1    g255(.A(new_n676), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n678), .B(new_n679), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n682), .A2(G1986), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(G1986), .ZN(new_n684));
  AND2_X1   g259(.A1(KEYINPUT91), .A2(G29), .ZN(new_n685));
  NOR2_X1   g260(.A1(KEYINPUT91), .A2(G29), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G25), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n475), .A2(G131), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n477), .A2(G119), .ZN(new_n691));
  OR2_X1    g266(.A1(G95), .A2(G2105), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n692), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n689), .B1(new_n695), .B2(new_n688), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT35), .B(G1991), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n683), .A2(new_n684), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G23), .ZN(new_n701));
  INV_X1    g276(.A(G288), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT33), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1976), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n700), .A2(G6), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G305), .B2(G16), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT32), .B(G1981), .Z(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n681), .A2(G22), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G166), .B2(new_n681), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(G1971), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n707), .A2(new_n708), .B1(new_n711), .B2(G1971), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n705), .A2(new_n709), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n699), .B1(new_n714), .B2(KEYINPUT34), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n715), .B1(KEYINPUT34), .B2(new_n714), .C1(new_n697), .C2(new_n696), .ZN(new_n716));
  NAND2_X1  g291(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n688), .A2(G35), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n688), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT104), .B(KEYINPUT29), .ZN(new_n721));
  INV_X1    g296(.A(G2090), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n720), .B(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n716), .A2(new_n717), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n688), .B1(new_n727), .B2(G34), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT99), .Z(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n727), .B2(G34), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G160), .B2(G29), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(G2084), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT102), .Z(new_n733));
  NOR2_X1   g308(.A1(new_n542), .A2(new_n681), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G19), .B2(new_n681), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G1341), .ZN(new_n737));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G32), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n475), .A2(G141), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n477), .A2(G129), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT26), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n610), .A2(G105), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n740), .A2(new_n741), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n739), .B1(new_n746), .B2(new_n738), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT100), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  NOR2_X1   g325(.A1(G16), .A2(G21), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G168), .B2(G16), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n749), .A2(new_n750), .B1(G1966), .B2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n752), .ZN(new_n754));
  INV_X1    g329(.A(G1966), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n754), .A2(new_n755), .B1(new_n736), .B2(G1341), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n733), .A2(new_n737), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(KEYINPUT28), .B1(new_n688), .B2(G26), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n688), .A2(KEYINPUT28), .A3(G26), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n475), .A2(G140), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n477), .A2(G128), .ZN(new_n762));
  OR3_X1    g337(.A1(KEYINPUT95), .A2(G104), .A3(G2105), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n459), .A2(G116), .ZN(new_n764));
  OAI21_X1  g339(.A(KEYINPUT95), .B1(G104), .B2(G2105), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n763), .A2(new_n764), .A3(G2104), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n761), .A2(new_n762), .A3(new_n766), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n758), .B(new_n760), .C1(new_n767), .C2(G29), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G28), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n771), .B2(KEYINPUT30), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(KEYINPUT30), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g348(.A1(G5), .A2(G16), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G171), .B2(G16), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n773), .B1(new_n775), .B2(G1961), .C1(new_n621), .C2(new_n688), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n770), .B(new_n776), .C1(G1961), .C2(new_n775), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT101), .B(KEYINPUT31), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G11), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n681), .A2(KEYINPUT23), .A3(G20), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT23), .ZN(new_n781));
  INV_X1    g356(.A(G20), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n676), .B2(new_n782), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n780), .B(new_n783), .C1(new_n600), .C2(new_n700), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G1956), .Z(new_n785));
  INV_X1    g360(.A(new_n750), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n731), .A2(G2084), .B1(new_n748), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n777), .A2(new_n779), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n609), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(new_n459), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n475), .A2(G139), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n610), .A2(G103), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n790), .A2(new_n791), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n792), .B(new_n795), .C1(new_n789), .C2(new_n459), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(KEYINPUT97), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n738), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n738), .B2(G33), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT98), .B(G2072), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n596), .A2(new_n700), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G4), .B2(new_n700), .ZN(new_n804));
  INV_X1    g379(.A(G1348), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT103), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n688), .A2(G27), .ZN(new_n808));
  AOI211_X1 g383(.A(new_n807), .B(new_n808), .C1(new_n498), .C2(new_n687), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n807), .B2(new_n808), .ZN(new_n810));
  INV_X1    g385(.A(G2078), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n804), .A2(new_n805), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n806), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NOR4_X1   g389(.A1(new_n757), .A2(new_n788), .A3(new_n802), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n718), .A2(new_n724), .A3(new_n726), .A4(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  AOI22_X1  g392(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n507), .ZN(new_n819));
  INV_X1    g394(.A(G93), .ZN(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n510), .A2(new_n820), .B1(new_n512), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G860), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  INV_X1    g401(.A(new_n542), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(new_n823), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n824), .A2(new_n542), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n596), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n833), .A2(KEYINPUT105), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(KEYINPUT105), .B1(new_n833), .B2(new_n834), .ZN(new_n836));
  OR3_X1    g411(.A1(new_n835), .A2(new_n836), .A3(G860), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n833), .A2(new_n834), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n826), .B1(new_n837), .B2(new_n838), .ZN(G145));
  NAND2_X1  g414(.A1(new_n475), .A2(G142), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n477), .A2(G130), .ZN(new_n841));
  NOR2_X1   g416(.A1(G106), .A2(G2105), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(new_n459), .B2(G118), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n498), .B(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(new_n746), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n746), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n695), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n694), .A3(new_n847), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n796), .A2(new_n798), .A3(KEYINPUT106), .ZN(new_n852));
  INV_X1    g427(.A(new_n767), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n796), .A2(new_n798), .A3(KEYINPUT106), .A4(new_n767), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n612), .ZN(new_n857));
  INV_X1    g432(.A(new_n612), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n858), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n849), .A2(new_n857), .A3(new_n859), .A4(new_n850), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n621), .B(G160), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(G162), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G37), .ZN(new_n867));
  INV_X1    g442(.A(new_n865), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n861), .A2(new_n862), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n866), .A2(KEYINPUT107), .A3(new_n867), .A4(new_n869), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT40), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(G395));
  XNOR2_X1  g453(.A(new_n830), .B(KEYINPUT108), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n605), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n600), .B1(new_n587), .B2(new_n595), .ZN(new_n881));
  INV_X1    g456(.A(new_n594), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(new_n592), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(G299), .A3(new_n586), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(KEYINPUT109), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n884), .ZN(new_n888));
  AOI21_X1  g463(.A(G299), .B1(new_n883), .B2(new_n586), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n881), .A2(KEYINPUT41), .A3(new_n884), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT109), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n880), .A2(new_n887), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n885), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n894), .B1(new_n895), .B2(new_n880), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT112), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G305), .B(G166), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT110), .ZN(new_n900));
  XNOR2_X1  g475(.A(G290), .B(new_n702), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n900), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(new_n899), .ZN(new_n904));
  XNOR2_X1  g479(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n894), .B(KEYINPUT112), .C1(new_n895), .C2(new_n880), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n898), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n896), .A2(new_n897), .A3(new_n906), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(G868), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT113), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n823), .A2(G868), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT113), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n909), .A2(new_n914), .A3(G868), .A4(new_n910), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(G295));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(G331));
  NAND2_X1  g492(.A1(new_n890), .A2(KEYINPUT117), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT117), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n885), .A2(new_n919), .A3(new_n886), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n918), .A2(new_n920), .B1(new_n895), .B2(KEYINPUT41), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT118), .ZN(new_n923));
  NOR2_X1   g498(.A1(G286), .A2(G171), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G286), .A2(G171), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n925), .A2(new_n829), .A3(new_n828), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n828), .A2(new_n829), .ZN(new_n928));
  INV_X1    g503(.A(new_n926), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(new_n929), .B2(new_n924), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n922), .A2(new_n923), .A3(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n927), .A2(new_n930), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT118), .B1(new_n921), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n927), .A2(new_n930), .A3(KEYINPUT114), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT114), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n830), .A2(new_n936), .A3(new_n925), .A4(new_n926), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n885), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n932), .A2(new_n934), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n904), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n933), .A2(KEYINPUT115), .A3(new_n885), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT115), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(new_n931), .B2(new_n895), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n893), .A2(new_n887), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n943), .B(new_n945), .C1(new_n946), .C2(new_n938), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(new_n904), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n941), .A2(new_n942), .A3(new_n867), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n904), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT116), .B1(new_n951), .B2(new_n867), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT116), .ZN(new_n953));
  AOI211_X1 g528(.A(new_n953), .B(G37), .C1(new_n947), .C2(new_n904), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n952), .A2(new_n954), .A3(new_n948), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n950), .B1(new_n955), .B2(new_n942), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n952), .A2(new_n954), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT43), .B1(new_n959), .B2(new_n949), .ZN(new_n960));
  AND4_X1   g535(.A1(KEYINPUT43), .A2(new_n941), .A3(new_n867), .A4(new_n949), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT44), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n498), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT119), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  AOI21_X1  g542(.A(G1384), .B1(new_n490), .B2(new_n497), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT119), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(G160), .A2(G40), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OR3_X1    g550(.A1(new_n975), .A2(KEYINPUT120), .A3(new_n745), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n767), .B(new_n769), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n974), .B2(new_n746), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT120), .B1(new_n975), .B2(new_n745), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n694), .B(new_n697), .Z(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n982), .A2(KEYINPUT121), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(KEYINPUT121), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n973), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n976), .A2(new_n979), .A3(new_n980), .A4(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n973), .ZN(new_n987));
  OR2_X1    g562(.A1(G290), .A2(G1986), .ZN(new_n988));
  NAND2_X1  g563(.A1(G290), .A2(G1986), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1981), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n570), .A2(new_n992), .A3(new_n571), .A4(new_n572), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G40), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n468), .A2(new_n995), .A3(new_n473), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n968), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G8), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n571), .ZN(new_n1000));
  OAI21_X1  g575(.A(G1981), .B1(new_n1000), .B2(new_n569), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n993), .A2(new_n1001), .A3(KEYINPUT49), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n993), .A2(new_n1001), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n999), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n994), .B1(new_n1008), .B2(new_n702), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n702), .A2(G1976), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(G288), .B2(new_n1007), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n999), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n998), .B1(G1976), .B2(new_n702), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1006), .B(new_n1012), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT45), .B1(new_n498), .B2(new_n964), .ZN(new_n1016));
  AOI211_X1 g591(.A(new_n967), .B(G1384), .C1(new_n490), .C2(new_n497), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n972), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT50), .B1(new_n498), .B2(new_n964), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  AOI211_X1 g595(.A(new_n1020), .B(G1384), .C1(new_n490), .C2(new_n497), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n996), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  OAI22_X1  g597(.A1(new_n1018), .A2(G1971), .B1(new_n1022), .B2(G2090), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G303), .A2(G8), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT55), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(G8), .A3(new_n1026), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1009), .A2(new_n998), .B1(new_n1015), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1023), .A2(G8), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n1025), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1015), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n1027), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n972), .B1(KEYINPUT45), .B2(new_n968), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n965), .A2(new_n967), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n755), .ZN(new_n1037));
  INV_X1    g612(.A(G2084), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(new_n996), .C1(new_n1019), .C2(new_n1021), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1033), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1032), .A2(KEYINPUT63), .A3(G168), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT63), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1030), .A2(new_n1031), .A3(new_n1040), .A4(new_n1027), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1042), .B1(new_n1043), .B2(G286), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1028), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n1046));
  XNOR2_X1  g621(.A(G299), .B(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT56), .B(G2072), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1034), .A2(new_n1035), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1022), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1047), .B(new_n1049), .C1(new_n1050), .C2(G1956), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1051), .B(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n596), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1022), .A2(new_n805), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n968), .A2(new_n769), .A3(new_n996), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1054), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1049), .B1(new_n1050), .B2(G1956), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1047), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1053), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT58), .B(G1341), .Z(new_n1063));
  AND2_X1   g638(.A1(new_n997), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n1018), .B2(new_n974), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT59), .B1(new_n1065), .B2(new_n827), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1036), .A2(G1996), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1067), .B(new_n542), .C1(new_n1068), .C2(new_n1064), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1056), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n596), .B(new_n1071), .C1(new_n1022), .C2(new_n805), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT60), .B1(new_n1057), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT60), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1055), .A2(new_n1074), .A3(new_n596), .A4(new_n1056), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1061), .A2(KEYINPUT61), .A3(new_n1051), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1061), .A2(KEYINPUT123), .A3(KEYINPUT61), .A4(new_n1051), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1076), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT61), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1061), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1082), .B1(new_n1053), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1062), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1034), .A2(new_n1035), .A3(new_n811), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n1087));
  INV_X1    g662(.A(G1961), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1086), .A2(new_n1087), .B1(new_n1022), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G171), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT124), .B(G2078), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n971), .A2(KEYINPUT53), .A3(new_n1034), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1091), .B(new_n1092), .C1(G171), .C2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(KEYINPUT125), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1097), .A2(G301), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1090), .A2(G301), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT54), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1096), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(G168), .A2(new_n1033), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT51), .B1(new_n1040), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1039), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1966), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1107));
  OAI21_X1  g682(.A(G8), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1104), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1105), .A2(new_n1111), .B1(new_n1104), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1030), .A2(new_n1031), .A3(new_n1027), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1103), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1045), .B1(new_n1085), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1112), .A2(new_n1104), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1111), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1109), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1032), .B1(new_n1122), .B2(KEYINPUT62), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1091), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1113), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1118), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1091), .B1(new_n1122), .B2(KEYINPUT62), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1114), .B1(new_n1113), .B2(new_n1125), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(KEYINPUT126), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n991), .B1(new_n1117), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n987), .B1(new_n746), .B2(new_n977), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT46), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n975), .B1(KEYINPUT127), .B2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT127), .B(KEYINPUT46), .Z(new_n1136));
  AOI211_X1 g711(.A(new_n1133), .B(new_n1135), .C1(new_n975), .C2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT47), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n694), .A2(new_n697), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n976), .A2(new_n979), .A3(new_n980), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n853), .A2(new_n769), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n987), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n987), .A2(new_n988), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT48), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n986), .A2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1138), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1132), .A2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g722(.A(G401), .B1(new_n872), .B2(new_n873), .ZN(new_n1149));
  INV_X1    g723(.A(G319), .ZN(new_n1150));
  NOR3_X1   g724(.A1(G227), .A2(new_n1150), .A3(G229), .ZN(new_n1151));
  AND3_X1   g725(.A1(new_n1149), .A2(new_n956), .A3(new_n1151), .ZN(G308));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n956), .A3(new_n1151), .ZN(G225));
endmodule


