

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737;

  NOR2_X2 U369 ( .A1(G953), .A2(G237), .ZN(n494) );
  XNOR2_X1 U370 ( .A(n452), .B(n451), .ZN(n454) );
  NOR2_X1 U371 ( .A1(n513), .A2(n526), .ZN(n349) );
  AND2_X4 U372 ( .A1(n403), .A2(n401), .ZN(n699) );
  NOR2_X2 U373 ( .A1(n529), .A2(n528), .ZN(n531) );
  INV_X2 U374 ( .A(n533), .ZN(n516) );
  NOR2_X1 U375 ( .A1(n615), .A2(n707), .ZN(n362) );
  NOR2_X1 U376 ( .A1(n622), .A2(n707), .ZN(n624) );
  NAND2_X1 U377 ( .A1(n735), .A2(n737), .ZN(n593) );
  XNOR2_X1 U378 ( .A(n412), .B(KEYINPUT95), .ZN(n481) );
  XNOR2_X1 U379 ( .A(n454), .B(n453), .ZN(n504) );
  OR2_X1 U380 ( .A1(n390), .A2(n389), .ZN(n401) );
  AND2_X1 U381 ( .A1(n609), .A2(n608), .ZN(n726) );
  XNOR2_X1 U382 ( .A(n364), .B(n363), .ZN(n609) );
  NAND2_X1 U383 ( .A1(n594), .A2(n595), .ZN(n364) );
  AND2_X1 U384 ( .A1(n543), .A2(n617), .ZN(n387) );
  XNOR2_X1 U385 ( .A(n487), .B(KEYINPUT101), .ZN(n628) );
  NOR2_X1 U386 ( .A1(n473), .A2(n549), .ZN(n474) );
  XOR2_X1 U387 ( .A(KEYINPUT108), .B(n512), .Z(n643) );
  AND2_X1 U388 ( .A1(n588), .A2(n561), .ZN(n544) );
  XNOR2_X1 U389 ( .A(n365), .B(n348), .ZN(n559) );
  NAND2_X1 U390 ( .A1(n552), .A2(n588), .ZN(n388) );
  XNOR2_X1 U391 ( .A(n450), .B(n449), .ZN(n563) );
  XNOR2_X1 U392 ( .A(n425), .B(n424), .ZN(n552) );
  XNOR2_X1 U393 ( .A(n499), .B(n498), .ZN(n525) );
  XNOR2_X1 U394 ( .A(n708), .B(n419), .ZN(n612) );
  XNOR2_X1 U395 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U396 ( .A(n413), .B(n481), .ZN(n708) );
  XNOR2_X1 U397 ( .A(n379), .B(G104), .ZN(n493) );
  XNOR2_X1 U398 ( .A(G113), .B(G122), .ZN(n379) );
  OR2_X1 U399 ( .A1(n606), .A2(n394), .ZN(n393) );
  NOR2_X1 U400 ( .A1(n710), .A2(n356), .ZN(n368) );
  XNOR2_X1 U401 ( .A(n387), .B(KEYINPUT44), .ZN(n386) );
  INV_X1 U402 ( .A(KEYINPUT75), .ZN(n378) );
  NAND2_X1 U403 ( .A1(n351), .A2(n371), .ZN(n370) );
  NOR2_X1 U404 ( .A1(n580), .A2(n645), .ZN(n369) );
  XOR2_X1 U405 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n453) );
  INV_X1 U406 ( .A(KEYINPUT70), .ZN(n451) );
  XNOR2_X1 U407 ( .A(KEYINPUT4), .B(G131), .ZN(n438) );
  NAND2_X1 U408 ( .A1(n386), .A2(n350), .ZN(n384) );
  INV_X1 U409 ( .A(n505), .ZN(n506) );
  XNOR2_X1 U410 ( .A(n381), .B(n495), .ZN(n380) );
  XNOR2_X1 U411 ( .A(n383), .B(n382), .ZN(n381) );
  XNOR2_X1 U412 ( .A(KEYINPUT104), .B(KEYINPUT103), .ZN(n383) );
  XNOR2_X1 U413 ( .A(G101), .B(G107), .ZN(n439) );
  XOR2_X1 U414 ( .A(G110), .B(G104), .Z(n440) );
  NOR2_X1 U415 ( .A1(n726), .A2(n402), .ZN(n389) );
  NAND2_X1 U416 ( .A1(n368), .A2(n367), .ZN(n390) );
  NAND2_X1 U417 ( .A1(n726), .A2(n392), .ZN(n367) );
  XNOR2_X1 U418 ( .A(n533), .B(n532), .ZN(n561) );
  INV_X1 U419 ( .A(KEYINPUT110), .ZN(n532) );
  XNOR2_X1 U420 ( .A(n511), .B(n510), .ZN(n526) );
  INV_X1 U421 ( .A(KEYINPUT47), .ZN(n373) );
  NAND2_X1 U422 ( .A1(n375), .A2(n374), .ZN(n371) );
  NOR2_X1 U423 ( .A1(n633), .A2(n378), .ZN(n374) );
  NOR2_X1 U424 ( .A1(n643), .A2(n349), .ZN(n655) );
  INV_X1 U425 ( .A(G237), .ZN(n420) );
  XNOR2_X1 U426 ( .A(G137), .B(G113), .ZN(n478) );
  XNOR2_X1 U427 ( .A(KEYINPUT3), .B(KEYINPUT73), .ZN(n409) );
  NAND2_X1 U428 ( .A1(n358), .A2(n375), .ZN(n385) );
  INV_X1 U429 ( .A(n642), .ZN(n359) );
  INV_X1 U430 ( .A(n628), .ZN(n360) );
  XNOR2_X1 U431 ( .A(G131), .B(KEYINPUT11), .ZN(n382) );
  INV_X1 U432 ( .A(KEYINPUT48), .ZN(n363) );
  NAND2_X1 U433 ( .A1(G234), .A2(G237), .ZN(n430) );
  XNOR2_X1 U434 ( .A(n573), .B(n429), .ZN(n566) );
  XNOR2_X1 U435 ( .A(n719), .B(n462), .ZN(n463) );
  INV_X1 U436 ( .A(G119), .ZN(n462) );
  AND2_X1 U437 ( .A1(n606), .A2(n355), .ZN(n399) );
  NAND2_X1 U438 ( .A1(n607), .A2(n400), .ZN(n398) );
  NAND2_X1 U439 ( .A1(n404), .A2(n397), .ZN(n396) );
  NAND2_X1 U440 ( .A1(n400), .A2(KEYINPUT2), .ZN(n397) );
  NAND2_X1 U441 ( .A1(n391), .A2(KEYINPUT65), .ZN(n394) );
  XNOR2_X1 U442 ( .A(n521), .B(n405), .ZN(n682) );
  XNOR2_X1 U443 ( .A(KEYINPUT90), .B(KEYINPUT39), .ZN(n584) );
  BUF_X1 U444 ( .A(n552), .Z(n601) );
  XNOR2_X1 U445 ( .A(n525), .B(KEYINPUT105), .ZN(n513) );
  XNOR2_X1 U446 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U447 ( .A(n380), .B(n493), .ZN(n496) );
  XNOR2_X1 U448 ( .A(n444), .B(n443), .ZN(n445) );
  NOR2_X1 U449 ( .A1(n728), .A2(G952), .ZN(n707) );
  INV_X1 U450 ( .A(n401), .ZN(n648) );
  NOR2_X1 U451 ( .A1(n372), .A2(n665), .ZN(n645) );
  XNOR2_X1 U452 ( .A(n575), .B(n353), .ZN(n372) );
  OR2_X1 U453 ( .A1(n540), .A2(n535), .ZN(n632) );
  BUF_X1 U454 ( .A(n628), .Z(n366) );
  AND2_X1 U455 ( .A1(n376), .A2(n373), .ZN(n347) );
  XOR2_X1 U456 ( .A(n469), .B(n468), .Z(n348) );
  AND2_X1 U457 ( .A1(n385), .A2(n625), .ZN(n350) );
  AND2_X1 U458 ( .A1(n347), .A2(n377), .ZN(n351) );
  XNOR2_X1 U459 ( .A(n655), .B(KEYINPUT86), .ZN(n567) );
  INV_X1 U460 ( .A(n567), .ZN(n375) );
  NOR2_X1 U461 ( .A1(n606), .A2(KEYINPUT2), .ZN(n352) );
  XOR2_X1 U462 ( .A(n568), .B(KEYINPUT36), .Z(n353) );
  XOR2_X1 U463 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n354) );
  INV_X1 U464 ( .A(n607), .ZN(n404) );
  INV_X1 U465 ( .A(KEYINPUT2), .ZN(n391) );
  INV_X1 U466 ( .A(KEYINPUT88), .ZN(n402) );
  AND2_X1 U467 ( .A1(n404), .A2(n400), .ZN(n355) );
  AND2_X1 U468 ( .A1(KEYINPUT88), .A2(n391), .ZN(n356) );
  AND2_X1 U469 ( .A1(n398), .A2(n396), .ZN(n357) );
  XOR2_X2 U470 ( .A(KEYINPUT6), .B(n516), .Z(n569) );
  NAND2_X1 U471 ( .A1(n360), .A2(n359), .ZN(n358) );
  NOR2_X2 U472 ( .A1(n697), .A2(n707), .ZN(n698) );
  NAND2_X1 U473 ( .A1(n504), .A2(G221), .ZN(n458) );
  XNOR2_X1 U474 ( .A(n585), .B(n584), .ZN(n596) );
  NOR2_X1 U475 ( .A1(n361), .A2(n551), .ZN(n583) );
  XNOR2_X1 U476 ( .A(n550), .B(KEYINPUT77), .ZN(n361) );
  XNOR2_X1 U477 ( .A(n362), .B(n616), .ZN(G51) );
  NOR2_X1 U478 ( .A1(n705), .A2(G902), .ZN(n365) );
  NAND2_X1 U479 ( .A1(n395), .A2(n393), .ZN(n403) );
  NAND2_X1 U480 ( .A1(n570), .A2(n349), .ZN(n571) );
  AND2_X1 U481 ( .A1(n370), .A2(n369), .ZN(n581) );
  NAND2_X1 U482 ( .A1(n633), .A2(n378), .ZN(n376) );
  NAND2_X1 U483 ( .A1(n567), .A2(n378), .ZN(n377) );
  INV_X1 U484 ( .A(n522), .ZN(n473) );
  NAND2_X1 U485 ( .A1(n522), .A2(n406), .ZN(n515) );
  XNOR2_X2 U486 ( .A(n436), .B(n435), .ZN(n522) );
  XNOR2_X2 U487 ( .A(n384), .B(n354), .ZN(n710) );
  NOR2_X2 U488 ( .A1(n710), .A2(n605), .ZN(n606) );
  NAND2_X1 U489 ( .A1(n566), .A2(n434), .ZN(n436) );
  XNOR2_X2 U490 ( .A(n388), .B(KEYINPUT92), .ZN(n573) );
  AND2_X1 U491 ( .A1(n402), .A2(KEYINPUT2), .ZN(n392) );
  NOR2_X1 U492 ( .A1(n399), .A2(n357), .ZN(n395) );
  INV_X1 U493 ( .A(KEYINPUT65), .ZN(n400) );
  XNOR2_X2 U494 ( .A(G146), .B(G125), .ZN(n461) );
  XNOR2_X1 U495 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n405) );
  XOR2_X1 U496 ( .A(n514), .B(KEYINPUT109), .Z(n406) );
  INV_X1 U497 ( .A(KEYINPUT5), .ZN(n477) );
  XNOR2_X1 U498 ( .A(n478), .B(n477), .ZN(n479) );
  INV_X1 U499 ( .A(G469), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n480), .B(n479), .ZN(n482) );
  INV_X1 U501 ( .A(KEYINPUT80), .ZN(n441) );
  NAND2_X1 U502 ( .A1(n662), .A2(n661), .ZN(n666) );
  XNOR2_X1 U503 ( .A(n448), .B(KEYINPUT72), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n500), .B(n407), .ZN(n408) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n509), .B(n508), .ZN(n700) );
  INV_X2 U507 ( .A(G953), .ZN(n728) );
  XOR2_X2 U508 ( .A(G116), .B(G107), .Z(n500) );
  XOR2_X1 U509 ( .A(KEYINPUT16), .B(G110), .Z(n407) );
  XNOR2_X1 U510 ( .A(n408), .B(n493), .ZN(n413) );
  INV_X1 U511 ( .A(n409), .ZN(n411) );
  XNOR2_X1 U512 ( .A(G119), .B(G101), .ZN(n410) );
  XNOR2_X1 U513 ( .A(n411), .B(n410), .ZN(n412) );
  NAND2_X1 U514 ( .A1(n728), .A2(G224), .ZN(n414) );
  XNOR2_X1 U515 ( .A(n414), .B(KEYINPUT4), .ZN(n415) );
  XNOR2_X1 U516 ( .A(n415), .B(n461), .ZN(n418) );
  XNOR2_X1 U517 ( .A(G143), .B(G128), .ZN(n437) );
  XNOR2_X1 U518 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n416) );
  XNOR2_X1 U519 ( .A(n437), .B(n416), .ZN(n417) );
  XNOR2_X1 U520 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U521 ( .A(KEYINPUT15), .B(G902), .ZN(n607) );
  NAND2_X1 U522 ( .A1(n612), .A2(n607), .ZN(n425) );
  INV_X1 U523 ( .A(G902), .ZN(n421) );
  NAND2_X1 U524 ( .A1(n421), .A2(n420), .ZN(n426) );
  NAND2_X1 U525 ( .A1(n426), .A2(G210), .ZN(n423) );
  INV_X1 U526 ( .A(KEYINPUT96), .ZN(n422) );
  XNOR2_X1 U527 ( .A(n423), .B(n422), .ZN(n424) );
  NAND2_X1 U528 ( .A1(n426), .A2(G214), .ZN(n428) );
  INV_X1 U529 ( .A(KEYINPUT97), .ZN(n427) );
  XNOR2_X1 U530 ( .A(n428), .B(n427), .ZN(n588) );
  XNOR2_X1 U531 ( .A(KEYINPUT78), .B(KEYINPUT19), .ZN(n429) );
  XNOR2_X1 U532 ( .A(n430), .B(KEYINPUT14), .ZN(n431) );
  NAND2_X1 U533 ( .A1(G952), .A2(n431), .ZN(n680) );
  NOR2_X1 U534 ( .A1(G953), .A2(n680), .ZN(n548) );
  INV_X1 U535 ( .A(G898), .ZN(n713) );
  NAND2_X1 U536 ( .A1(G953), .A2(n713), .ZN(n709) );
  NAND2_X1 U537 ( .A1(G902), .A2(n431), .ZN(n545) );
  NOR2_X1 U538 ( .A1(n709), .A2(n545), .ZN(n432) );
  OR2_X1 U539 ( .A1(n548), .A2(n432), .ZN(n433) );
  XNOR2_X1 U540 ( .A(n433), .B(KEYINPUT98), .ZN(n434) );
  INV_X1 U541 ( .A(KEYINPUT0), .ZN(n435) );
  XNOR2_X1 U542 ( .A(n437), .B(G134), .ZN(n505) );
  XNOR2_X1 U543 ( .A(n505), .B(n438), .ZN(n483) );
  XNOR2_X1 U544 ( .A(G137), .B(G140), .ZN(n459) );
  XNOR2_X1 U545 ( .A(n483), .B(n459), .ZN(n720) );
  XNOR2_X1 U546 ( .A(G146), .B(KEYINPUT79), .ZN(n446) );
  XNOR2_X1 U547 ( .A(n440), .B(n439), .ZN(n444) );
  NAND2_X1 U548 ( .A1(G227), .A2(n728), .ZN(n442) );
  XNOR2_X1 U549 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U550 ( .A(n720), .B(n447), .ZN(n690) );
  NOR2_X1 U551 ( .A1(G902), .A2(n690), .ZN(n450) );
  NAND2_X1 U552 ( .A1(G234), .A2(n728), .ZN(n452) );
  XOR2_X1 U553 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n456) );
  XNOR2_X1 U554 ( .A(G128), .B(KEYINPUT23), .ZN(n455) );
  XNOR2_X1 U555 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U556 ( .A(n458), .B(n457), .ZN(n466) );
  XNOR2_X1 U557 ( .A(G110), .B(n459), .ZN(n464) );
  INV_X1 U558 ( .A(KEYINPUT10), .ZN(n460) );
  XNOR2_X2 U559 ( .A(n461), .B(n460), .ZN(n719) );
  XNOR2_X1 U560 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U561 ( .A(n466), .B(n465), .ZN(n705) );
  XOR2_X1 U562 ( .A(KEYINPUT99), .B(KEYINPUT25), .Z(n469) );
  NAND2_X1 U563 ( .A1(G234), .A2(n607), .ZN(n467) );
  XNOR2_X1 U564 ( .A(KEYINPUT20), .B(n467), .ZN(n470) );
  NAND2_X1 U565 ( .A1(n470), .A2(G217), .ZN(n468) );
  INV_X1 U566 ( .A(n559), .ZN(n662) );
  NAND2_X1 U567 ( .A1(n470), .A2(G221), .ZN(n471) );
  XNOR2_X1 U568 ( .A(KEYINPUT21), .B(n471), .ZN(n557) );
  INV_X1 U569 ( .A(n557), .ZN(n661) );
  INV_X1 U570 ( .A(n666), .ZN(n472) );
  NAND2_X1 U571 ( .A1(n563), .A2(n472), .ZN(n549) );
  XNOR2_X1 U572 ( .A(n474), .B(KEYINPUT100), .ZN(n486) );
  XOR2_X1 U573 ( .A(G116), .B(G146), .Z(n476) );
  NAND2_X1 U574 ( .A1(n494), .A2(G210), .ZN(n475) );
  XNOR2_X1 U575 ( .A(n476), .B(n475), .ZN(n480) );
  XNOR2_X1 U576 ( .A(n482), .B(n481), .ZN(n484) );
  XOR2_X1 U577 ( .A(n484), .B(n483), .Z(n619) );
  NOR2_X1 U578 ( .A1(G902), .A2(n619), .ZN(n485) );
  XNOR2_X2 U579 ( .A(n485), .B(G472), .ZN(n533) );
  NAND2_X1 U580 ( .A1(n486), .A2(n533), .ZN(n487) );
  XNOR2_X1 U581 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n488) );
  XNOR2_X1 U582 ( .A(n563), .B(n488), .ZN(n517) );
  NOR2_X1 U583 ( .A1(n666), .A2(n517), .ZN(n520) );
  AND2_X1 U584 ( .A1(n516), .A2(n520), .ZN(n672) );
  NAND2_X1 U585 ( .A1(n522), .A2(n672), .ZN(n489) );
  XNOR2_X1 U586 ( .A(n489), .B(KEYINPUT31), .ZN(n642) );
  XOR2_X1 U587 ( .A(KEYINPUT102), .B(KEYINPUT12), .Z(n491) );
  XNOR2_X1 U588 ( .A(G143), .B(G140), .ZN(n490) );
  XNOR2_X1 U589 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U590 ( .A(n719), .B(n492), .ZN(n497) );
  NAND2_X1 U591 ( .A1(G214), .A2(n494), .ZN(n495) );
  XNOR2_X1 U592 ( .A(n497), .B(n496), .ZN(n694) );
  NOR2_X1 U593 ( .A1(G902), .A2(n694), .ZN(n499) );
  XNOR2_X1 U594 ( .A(KEYINPUT13), .B(G475), .ZN(n498) );
  XNOR2_X1 U595 ( .A(KEYINPUT107), .B(G478), .ZN(n511) );
  XNOR2_X1 U596 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n503) );
  XNOR2_X1 U597 ( .A(n500), .B(G122), .ZN(n501) );
  XNOR2_X1 U598 ( .A(n501), .B(KEYINPUT106), .ZN(n502) );
  XNOR2_X1 U599 ( .A(n503), .B(n502), .ZN(n509) );
  NAND2_X1 U600 ( .A1(n504), .A2(G217), .ZN(n507) );
  NOR2_X1 U601 ( .A1(G902), .A2(n700), .ZN(n510) );
  NAND2_X1 U602 ( .A1(n513), .A2(n526), .ZN(n512) );
  NOR2_X1 U603 ( .A1(n526), .A2(n525), .ZN(n653) );
  AND2_X1 U604 ( .A1(n653), .A2(n661), .ZN(n514) );
  XNOR2_X1 U605 ( .A(n515), .B(KEYINPUT22), .ZN(n540) );
  NOR2_X1 U606 ( .A1(n569), .A2(n559), .ZN(n518) );
  BUF_X1 U607 ( .A(n517), .Z(n665) );
  NAND2_X1 U608 ( .A1(n518), .A2(n665), .ZN(n519) );
  OR2_X1 U609 ( .A1(n540), .A2(n519), .ZN(n625) );
  NAND2_X1 U610 ( .A1(n520), .A2(n569), .ZN(n521) );
  NAND2_X1 U611 ( .A1(n682), .A2(n522), .ZN(n524) );
  XNOR2_X1 U612 ( .A(KEYINPUT34), .B(KEYINPUT82), .ZN(n523) );
  XNOR2_X1 U613 ( .A(n524), .B(n523), .ZN(n529) );
  NAND2_X1 U614 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U615 ( .A(KEYINPUT111), .B(n527), .ZN(n554) );
  INV_X1 U616 ( .A(n554), .ZN(n528) );
  XNOR2_X1 U617 ( .A(KEYINPUT81), .B(KEYINPUT35), .ZN(n530) );
  XNOR2_X1 U618 ( .A(n531), .B(n530), .ZN(n733) );
  NOR2_X1 U619 ( .A1(n561), .A2(n662), .ZN(n534) );
  NAND2_X1 U620 ( .A1(n534), .A2(n665), .ZN(n535) );
  INV_X1 U621 ( .A(n632), .ZN(n536) );
  NOR2_X1 U622 ( .A1(n733), .A2(n536), .ZN(n543) );
  NOR2_X1 U623 ( .A1(n665), .A2(n662), .ZN(n538) );
  XNOR2_X1 U624 ( .A(n569), .B(KEYINPUT83), .ZN(n537) );
  NAND2_X1 U625 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U626 ( .A1(n540), .A2(n539), .ZN(n542) );
  XOR2_X1 U627 ( .A(KEYINPUT66), .B(KEYINPUT32), .Z(n541) );
  XNOR2_X1 U628 ( .A(n542), .B(n541), .ZN(n617) );
  XOR2_X1 U629 ( .A(n544), .B(KEYINPUT30), .Z(n551) );
  OR2_X1 U630 ( .A1(n728), .A2(n545), .ZN(n546) );
  NOR2_X1 U631 ( .A1(G900), .A2(n546), .ZN(n547) );
  NOR2_X1 U632 ( .A1(n548), .A2(n547), .ZN(n556) );
  NOR2_X1 U633 ( .A1(n556), .A2(n549), .ZN(n550) );
  NAND2_X1 U634 ( .A1(n583), .A2(n601), .ZN(n553) );
  XNOR2_X1 U635 ( .A(n553), .B(KEYINPUT113), .ZN(n555) );
  NAND2_X1 U636 ( .A1(n555), .A2(n554), .ZN(n637) );
  NOR2_X1 U637 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U638 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U639 ( .A(KEYINPUT71), .B(n560), .ZN(n570) );
  AND2_X1 U640 ( .A1(n561), .A2(n570), .ZN(n562) );
  XOR2_X1 U641 ( .A(KEYINPUT28), .B(n562), .Z(n565) );
  INV_X1 U642 ( .A(n563), .ZN(n564) );
  NOR2_X2 U643 ( .A1(n565), .A2(n564), .ZN(n590) );
  NAND2_X1 U644 ( .A1(n590), .A2(n566), .ZN(n633) );
  XNOR2_X1 U645 ( .A(KEYINPUT91), .B(KEYINPUT114), .ZN(n568) );
  INV_X1 U646 ( .A(n569), .ZN(n572) );
  NOR2_X1 U647 ( .A1(n572), .A2(n571), .ZN(n598) );
  INV_X1 U648 ( .A(n573), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n598), .A2(n574), .ZN(n575) );
  NAND2_X1 U650 ( .A1(n655), .A2(KEYINPUT47), .ZN(n576) );
  XOR2_X1 U651 ( .A(n576), .B(KEYINPUT85), .Z(n579) );
  OR2_X1 U652 ( .A1(n633), .A2(KEYINPUT75), .ZN(n577) );
  NAND2_X1 U653 ( .A1(n577), .A2(KEYINPUT47), .ZN(n578) );
  NAND2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n580) );
  AND2_X1 U655 ( .A1(n637), .A2(n581), .ZN(n595) );
  XNOR2_X1 U656 ( .A(KEYINPUT76), .B(KEYINPUT38), .ZN(n582) );
  XOR2_X1 U657 ( .A(n582), .B(n601), .Z(n587) );
  NAND2_X1 U658 ( .A1(n583), .A2(n587), .ZN(n585) );
  NAND2_X1 U659 ( .A1(n349), .A2(n596), .ZN(n586) );
  XNOR2_X2 U660 ( .A(n586), .B(KEYINPUT40), .ZN(n735) );
  INV_X1 U661 ( .A(n587), .ZN(n651) );
  INV_X1 U662 ( .A(n588), .ZN(n650) );
  NOR2_X1 U663 ( .A1(n651), .A2(n650), .ZN(n657) );
  NAND2_X1 U664 ( .A1(n657), .A2(n653), .ZN(n589) );
  XNOR2_X1 U665 ( .A(n589), .B(KEYINPUT41), .ZN(n681) );
  NAND2_X1 U666 ( .A1(n590), .A2(n681), .ZN(n591) );
  XNOR2_X1 U667 ( .A(n591), .B(KEYINPUT42), .ZN(n737) );
  XNOR2_X1 U668 ( .A(KEYINPUT46), .B(KEYINPUT89), .ZN(n592) );
  XNOR2_X1 U669 ( .A(n593), .B(n592), .ZN(n594) );
  AND2_X1 U670 ( .A1(n596), .A2(n643), .ZN(n597) );
  XNOR2_X1 U671 ( .A(n597), .B(KEYINPUT115), .ZN(n732) );
  INV_X1 U672 ( .A(n732), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n598), .A2(n665), .ZN(n599) );
  NOR2_X1 U674 ( .A1(n650), .A2(n599), .ZN(n600) );
  XNOR2_X1 U675 ( .A(n600), .B(KEYINPUT43), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT112), .ZN(n734) );
  NOR2_X1 U678 ( .A1(n604), .A2(n734), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n699), .A2(G210), .ZN(n614) );
  XNOR2_X1 U681 ( .A(KEYINPUT55), .B(KEYINPUT84), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n610), .B(KEYINPUT54), .ZN(n611) );
  XNOR2_X1 U683 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U685 ( .A(KEYINPUT56), .B(KEYINPUT122), .ZN(n616) );
  XNOR2_X1 U686 ( .A(n617), .B(G119), .ZN(G21) );
  NAND2_X1 U687 ( .A1(n699), .A2(G472), .ZN(n621) );
  XNOR2_X1 U688 ( .A(KEYINPUT94), .B(KEYINPUT62), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U690 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U691 ( .A(KEYINPUT93), .B(KEYINPUT63), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n624), .B(n623), .ZN(G57) );
  INV_X1 U693 ( .A(n625), .ZN(n626) );
  XOR2_X1 U694 ( .A(G101), .B(n626), .Z(G3) );
  NAND2_X1 U695 ( .A1(n366), .A2(n349), .ZN(n627) );
  XNOR2_X1 U696 ( .A(n627), .B(G104), .ZN(G6) );
  XOR2_X1 U697 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n630) );
  NAND2_X1 U698 ( .A1(n366), .A2(n643), .ZN(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U700 ( .A(G107), .B(n631), .ZN(G9) );
  XNOR2_X1 U701 ( .A(G110), .B(n632), .ZN(G12) );
  XOR2_X1 U702 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n635) );
  INV_X1 U703 ( .A(n633), .ZN(n638) );
  NAND2_X1 U704 ( .A1(n638), .A2(n643), .ZN(n634) );
  XNOR2_X1 U705 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U706 ( .A(G128), .B(n636), .ZN(G30) );
  XNOR2_X1 U707 ( .A(G143), .B(n637), .ZN(G45) );
  NAND2_X1 U708 ( .A1(n638), .A2(n349), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n639), .B(G146), .ZN(G48) );
  XOR2_X1 U710 ( .A(G113), .B(KEYINPUT117), .Z(n641) );
  NAND2_X1 U711 ( .A1(n642), .A2(n349), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n641), .B(n640), .ZN(G15) );
  NAND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n644), .B(G116), .ZN(G18) );
  XNOR2_X1 U715 ( .A(n645), .B(KEYINPUT37), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n646), .B(KEYINPUT118), .ZN(n647) );
  XNOR2_X1 U717 ( .A(G125), .B(n647), .ZN(G27) );
  NOR2_X1 U718 ( .A1(n352), .A2(n648), .ZN(n649) );
  NOR2_X1 U719 ( .A1(n649), .A2(G953), .ZN(n686) );
  NAND2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n654), .B(KEYINPUT120), .ZN(n659) );
  INV_X1 U723 ( .A(n655), .ZN(n656) );
  NAND2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U726 ( .A1(n682), .A2(n660), .ZN(n676) );
  NOR2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U728 ( .A(n663), .B(KEYINPUT49), .ZN(n664) );
  NAND2_X1 U729 ( .A1(n533), .A2(n664), .ZN(n669) );
  NAND2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U731 ( .A(KEYINPUT50), .B(n667), .Z(n668) );
  NOR2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U733 ( .A(KEYINPUT119), .B(n670), .Z(n671) );
  NOR2_X1 U734 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U735 ( .A(KEYINPUT51), .B(n673), .ZN(n674) );
  NAND2_X1 U736 ( .A1(n674), .A2(n681), .ZN(n675) );
  NAND2_X1 U737 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U738 ( .A(n677), .B(KEYINPUT52), .ZN(n678) );
  XNOR2_X1 U739 ( .A(n678), .B(KEYINPUT121), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n684) );
  AND2_X1 U741 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U742 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U743 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U744 ( .A(KEYINPUT53), .B(n687), .Z(G75) );
  NAND2_X1 U745 ( .A1(n699), .A2(G469), .ZN(n689) );
  XOR2_X1 U746 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n688) );
  XNOR2_X1 U747 ( .A(n689), .B(n688), .ZN(n691) );
  XNOR2_X1 U748 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X1 U749 ( .A1(n707), .A2(n692), .ZN(G54) );
  NAND2_X1 U750 ( .A1(n699), .A2(G475), .ZN(n696) );
  XOR2_X1 U751 ( .A(KEYINPUT59), .B(KEYINPUT68), .Z(n693) );
  XNOR2_X1 U752 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U753 ( .A(KEYINPUT60), .B(n698), .ZN(G60) );
  NAND2_X1 U754 ( .A1(n699), .A2(G478), .ZN(n702) );
  XOR2_X1 U755 ( .A(n700), .B(KEYINPUT123), .Z(n701) );
  XNOR2_X1 U756 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U757 ( .A1(n707), .A2(n703), .ZN(G63) );
  NAND2_X1 U758 ( .A1(n699), .A2(G217), .ZN(n704) );
  XNOR2_X1 U759 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U760 ( .A1(n707), .A2(n706), .ZN(G66) );
  NAND2_X1 U761 ( .A1(n709), .A2(n708), .ZN(n718) );
  NOR2_X1 U762 ( .A1(n710), .A2(G953), .ZN(n716) );
  XOR2_X1 U763 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n712) );
  NAND2_X1 U764 ( .A1(G224), .A2(G953), .ZN(n711) );
  XNOR2_X1 U765 ( .A(n712), .B(n711), .ZN(n714) );
  NOR2_X1 U766 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U767 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U768 ( .A(n718), .B(n717), .ZN(G69) );
  XNOR2_X1 U769 ( .A(n720), .B(n719), .ZN(n727) );
  INV_X1 U770 ( .A(n727), .ZN(n721) );
  XOR2_X1 U771 ( .A(G227), .B(n721), .Z(n722) );
  NAND2_X1 U772 ( .A1(n722), .A2(G900), .ZN(n723) );
  XOR2_X1 U773 ( .A(KEYINPUT125), .B(n723), .Z(n724) );
  NAND2_X1 U774 ( .A1(G953), .A2(n724), .ZN(n725) );
  XNOR2_X1 U775 ( .A(n725), .B(KEYINPUT126), .ZN(n731) );
  XOR2_X1 U776 ( .A(n727), .B(n726), .Z(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n731), .A2(n730), .ZN(G72) );
  XNOR2_X1 U779 ( .A(G134), .B(n732), .ZN(G36) );
  XOR2_X1 U780 ( .A(n733), .B(G122), .Z(G24) );
  XOR2_X1 U781 ( .A(G140), .B(n734), .Z(G42) );
  XOR2_X1 U782 ( .A(n735), .B(G131), .Z(n736) );
  XNOR2_X1 U783 ( .A(KEYINPUT127), .B(n736), .ZN(G33) );
  XNOR2_X1 U784 ( .A(G137), .B(n737), .ZN(G39) );
endmodule

