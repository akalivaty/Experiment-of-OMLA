//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n561, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G234));
  NAND2_X1  g025(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT66), .Z(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  OR2_X1    g051(.A1(new_n465), .A2(new_n466), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n471), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  XNOR2_X1  g061(.A(KEYINPUT68), .B(G114), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n472), .C1(new_n465), .C2(new_n466), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT67), .Z(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT71), .B1(new_n497), .B2(KEYINPUT5), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(new_n497), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT70), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT71), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n507), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT69), .B1(new_n512), .B2(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(new_n509), .A3(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n511), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n510), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n517), .B1(new_n513), .B2(new_n515), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n507), .A2(G89), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(G543), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n524), .B(new_n526), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g108(.A1(G63), .A2(G651), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n533), .B1(new_n507), .B2(new_n535), .ZN(new_n536));
  AOI211_X1 g111(.A(KEYINPUT72), .B(new_n534), .C1(new_n500), .C2(new_n506), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n532), .A2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n509), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n527), .A2(G52), .A3(G543), .A4(new_n529), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n507), .A2(G90), .A3(new_n525), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n543), .B1(new_n542), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n541), .B1(new_n545), .B2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n500), .B2(new_n506), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT75), .B(G43), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n527), .A2(G543), .A3(new_n529), .A4(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n507), .A2(G81), .A3(new_n525), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(new_n563));
  XOR2_X1   g138(.A(new_n563), .B(KEYINPUT76), .Z(G188));
  INV_X1    g139(.A(G78), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT77), .B1(new_n565), .B2(new_n497), .ZN(new_n566));
  OR3_X1    g141(.A1(new_n565), .A2(new_n497), .A3(KEYINPUT77), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT71), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n568), .B1(new_n501), .B2(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n505), .B2(G543), .ZN(new_n570));
  AOI211_X1 g145(.A(new_n568), .B(new_n497), .C1(new_n502), .C2(new_n504), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g147(.A(KEYINPUT78), .B(G65), .Z(new_n573));
  OAI211_X1 g148(.A(new_n566), .B(new_n567), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n519), .B1(new_n500), .B2(new_n506), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n574), .A2(G651), .B1(G91), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT9), .B1(new_n530), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(G543), .B1(new_n525), .B2(new_n528), .ZN(new_n579));
  AOI211_X1 g154(.A(KEYINPUT73), .B(new_n517), .C1(new_n513), .C2(new_n515), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n581), .A2(new_n582), .A3(G53), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n576), .A2(new_n584), .ZN(G299));
  OR2_X1    g160(.A1(new_n532), .A2(new_n538), .ZN(G286));
  XOR2_X1   g161(.A(new_n521), .B(KEYINPUT79), .Z(G303));
  OR2_X1    g162(.A1(new_n507), .A2(G74), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(G87), .B2(new_n575), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n581), .A2(G49), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT80), .ZN(G288));
  NAND2_X1  g167(.A1(new_n575), .A2(G86), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n525), .A2(G48), .A3(G543), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n572), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n596), .B1(new_n599), .B2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n595), .A2(new_n600), .ZN(G305));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n507), .A2(new_n525), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n530), .A2(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(new_n509), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n605), .A2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n603), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n575), .A2(G92), .A3(new_n610), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n613), .A2(new_n614), .B1(G54), .B2(new_n581), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n500), .B2(new_n506), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n618));
  AND2_X1   g193(.A1(G79), .A2(G543), .ZN(new_n619));
  OR3_X1    g194(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n618), .B1(new_n617), .B2(new_n619), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(G651), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n609), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n609), .B1(new_n624), .B2(G868), .ZN(G321));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NOR2_X1   g202(.A1(G286), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G299), .B(KEYINPUT84), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n627), .ZN(G297));
  AOI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(new_n627), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n624), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n557), .A2(new_n627), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n623), .A2(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n627), .ZN(G323));
  XOR2_X1   g211(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n637));
  XNOR2_X1  g212(.A(G323), .B(new_n637), .ZN(G282));
  NAND2_X1  g213(.A1(new_n477), .A2(new_n473), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT13), .Z(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n471), .A2(G135), .ZN(new_n645));
  INV_X1    g220(.A(G123), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n472), .A2(G111), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  OAI221_X1 g223(.A(new_n645), .B1(new_n478), .B2(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(G2096), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n643), .A2(new_n644), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT86), .ZN(G156));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n658), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(G401));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT17), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT87), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n672), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n675), .B(new_n671), .C1(new_n668), .C2(new_n672), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n670), .A2(new_n668), .A3(new_n672), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT18), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT88), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(new_n693), .B(new_n692), .S(new_n685), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G23), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n591), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT33), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1976), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(G6), .ZN(new_n707));
  INV_X1    g282(.A(G305), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n702), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT32), .B(G1981), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G22), .ZN(new_n713));
  OR3_X1    g288(.A1(new_n713), .A2(KEYINPUT92), .A3(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(KEYINPUT92), .B1(new_n713), .B2(G16), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n714), .B(new_n715), .C1(G166), .C2(new_n702), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(G1971), .Z(new_n717));
  NAND4_X1  g292(.A1(new_n706), .A2(new_n711), .A3(new_n712), .A4(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT34), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(KEYINPUT34), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n702), .A2(G24), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n605), .A2(new_n607), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n702), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT91), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1986), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G25), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT89), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n471), .A2(G131), .ZN(new_n729));
  INV_X1    g304(.A(G119), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n472), .A2(G107), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n732));
  OAI221_X1 g307(.A(new_n729), .B1(new_n478), .B2(new_n730), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n728), .B1(new_n737), .B2(G29), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n738), .B(new_n740), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n719), .A2(new_n720), .A3(new_n725), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT36), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT25), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n471), .A2(G139), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n477), .A2(G127), .ZN(new_n750));
  NAND2_X1  g325(.A1(G115), .A2(G2104), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n472), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G29), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G29), .B2(G33), .ZN(new_n755));
  INV_X1    g330(.A(G2072), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(KEYINPUT24), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(KEYINPUT24), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n726), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G160), .B2(new_n726), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n757), .B(new_n758), .C1(G2084), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n726), .A2(G35), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G162), .B2(new_n726), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT29), .B(G2090), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n726), .A2(G26), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT28), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n471), .A2(G140), .ZN(new_n771));
  OR2_X1    g346(.A1(G104), .A2(G2105), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n772), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n773));
  INV_X1    g348(.A(G128), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n771), .B(new_n773), .C1(new_n774), .C2(new_n478), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n770), .B1(new_n775), .B2(G29), .ZN(new_n776));
  INV_X1    g351(.A(G2067), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT31), .B(G11), .Z(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT30), .B(G28), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n779), .B1(new_n726), .B2(new_n780), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n781), .B1(new_n726), .B2(new_n649), .C1(new_n763), .C2(G2084), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n768), .A2(new_n778), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G164), .A2(new_n726), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G27), .B2(new_n726), .ZN(new_n785));
  INV_X1    g360(.A(G2078), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n764), .A2(new_n783), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n702), .A2(G19), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n558), .B2(new_n702), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1341), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n471), .A2(G141), .B1(G105), .B2(new_n473), .ZN(new_n794));
  NAND3_X1  g369(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT26), .Z(new_n796));
  INV_X1    g371(.A(G129), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n794), .B(new_n796), .C1(new_n797), .C2(new_n478), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT94), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(KEYINPUT94), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G29), .ZN(new_n803));
  NOR2_X1   g378(.A1(G29), .A2(G32), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(KEYINPUT95), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(KEYINPUT95), .B2(new_n803), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT27), .B(G1996), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G168), .A2(new_n702), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n702), .B2(G21), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1966), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n793), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G4), .A2(G16), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n624), .B2(G16), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT93), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1348), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n702), .A2(G20), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT23), .Z(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G299), .B2(G16), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(G1956), .Z(new_n820));
  NOR3_X1   g395(.A1(new_n812), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n702), .A2(G5), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G171), .B2(new_n702), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT96), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n821), .B1(G1961), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(G1961), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT97), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n743), .A2(new_n828), .ZN(G150));
  INV_X1    g404(.A(G150), .ZN(G311));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n581), .A2(G55), .B1(new_n575), .B2(G93), .ZN(new_n832));
  INV_X1    g407(.A(G67), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n500), .B2(new_n506), .ZN(new_n834));
  AND2_X1   g409(.A1(G80), .A2(G543), .ZN(new_n835));
  OAI21_X1  g410(.A(G651), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n557), .A2(new_n831), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(G56), .B1(new_n570), .B2(new_n571), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n551), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n839), .A2(G651), .B1(G81), .B2(new_n575), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n840), .A2(KEYINPUT98), .A3(new_n841), .A4(new_n555), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n553), .A2(KEYINPUT98), .A3(new_n555), .A4(new_n556), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT99), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n837), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n832), .A2(new_n836), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n557), .A2(new_n831), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n842), .A2(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT38), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n623), .A2(new_n632), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT100), .ZN(new_n855));
  AOI21_X1  g430(.A(G860), .B1(new_n852), .B2(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n846), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(new_n649), .B(new_n475), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n484), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n801), .A2(new_n775), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n801), .A2(new_n775), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n495), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n495), .B1(new_n863), .B2(new_n864), .ZN(new_n867));
  OAI22_X1  g442(.A1(new_n866), .A2(new_n867), .B1(new_n752), .B2(new_n749), .ZN(new_n868));
  INV_X1    g443(.A(new_n867), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(new_n753), .A3(new_n865), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n479), .A2(G130), .ZN(new_n873));
  INV_X1    g448(.A(new_n471), .ZN(new_n874));
  INV_X1    g449(.A(G142), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n472), .A2(G118), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT101), .B1(G106), .B2(G2105), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  OAI221_X1 g455(.A(new_n873), .B1(new_n874), .B2(new_n875), .C1(new_n878), .C2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n737), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n737), .A2(new_n882), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n884), .A2(new_n885), .A3(new_n640), .ZN(new_n886));
  INV_X1    g461(.A(new_n640), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n735), .A2(new_n736), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT102), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n889), .B2(new_n883), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n881), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n640), .B1(new_n884), .B2(new_n885), .ZN(new_n892));
  INV_X1    g467(.A(new_n881), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n887), .A3(new_n883), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(KEYINPUT103), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT103), .B1(new_n891), .B2(new_n895), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n872), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n896), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n900), .A2(new_n871), .A3(new_n897), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n862), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n891), .A2(new_n895), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n862), .B1(new_n872), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n871), .B1(new_n900), .B2(new_n897), .ZN(new_n905));
  AOI21_X1  g480(.A(G37), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g483(.A1(new_n846), .A2(new_n627), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n591), .A2(new_n722), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n589), .A2(new_n590), .ZN(new_n911));
  NAND2_X1  g486(.A1(G290), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT104), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G305), .A2(G166), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n708), .A2(new_n521), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n910), .A2(new_n912), .A3(KEYINPUT104), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n917), .A2(new_n913), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n915), .A2(new_n914), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT42), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n849), .B(new_n635), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n623), .A2(G299), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n615), .A2(new_n622), .A3(new_n576), .A4(new_n584), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n924), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT41), .B1(new_n923), .B2(new_n924), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n926), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n921), .B(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n909), .B1(new_n931), .B2(new_n627), .ZN(G295));
  OAI21_X1  g507(.A(new_n909), .B1(new_n931), .B2(new_n627), .ZN(G331));
  INV_X1    g508(.A(G37), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n935));
  NAND2_X1  g510(.A1(G301), .A2(G286), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n542), .A2(new_n544), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT74), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(G168), .A3(new_n541), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n845), .B2(new_n848), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n847), .A2(new_n846), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n843), .A2(KEYINPUT99), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n843), .A2(KEYINPUT99), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n837), .A2(new_n842), .A3(new_n844), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n936), .A4(new_n941), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n943), .A2(new_n944), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n942), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n849), .A2(KEYINPUT105), .A3(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n951), .A2(new_n929), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n943), .A2(new_n955), .A3(new_n950), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n942), .B(KEYINPUT106), .C1(new_n845), .C2(new_n848), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n925), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n919), .B1(new_n913), .B2(new_n917), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n919), .B2(new_n913), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n935), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n956), .A2(new_n957), .ZN(new_n963));
  INV_X1    g538(.A(new_n925), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n951), .A2(new_n929), .A3(new_n953), .ZN(new_n966));
  AND4_X1   g541(.A1(new_n935), .A2(new_n965), .A3(new_n961), .A4(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n934), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n956), .A2(new_n929), .A3(new_n957), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n951), .A2(new_n953), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n969), .B1(new_n970), .B2(new_n925), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT108), .B1(new_n971), .B2(new_n920), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n956), .A2(new_n929), .A3(new_n957), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n925), .B1(new_n951), .B2(new_n953), .ZN(new_n974));
  OAI211_X1 g549(.A(KEYINPUT108), .B(new_n920), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n968), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n959), .A2(new_n935), .A3(new_n961), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n965), .A2(new_n961), .A3(new_n966), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT107), .ZN(new_n982));
  AOI21_X1  g557(.A(G37), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n920), .B1(new_n954), .B2(new_n958), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT43), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT44), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n978), .B1(new_n968), .B2(new_n977), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(KEYINPUT43), .A3(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n986), .B1(KEYINPUT44), .B2(new_n989), .ZN(G397));
  XNOR2_X1  g565(.A(new_n775), .B(G2067), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n801), .B2(G1996), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n470), .A2(new_n474), .A3(G40), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n492), .B2(new_n494), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT45), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1996), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n1000), .B(KEYINPUT109), .Z(new_n1001));
  AOI21_X1  g576(.A(new_n998), .B1(new_n1001), .B2(new_n802), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n888), .A2(new_n739), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n737), .A2(new_n740), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n996), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1006), .A2(KEYINPUT126), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(KEYINPUT126), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n997), .A2(G1986), .A3(G290), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT48), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  XOR2_X1   g586(.A(new_n1001), .B(KEYINPUT46), .Z(new_n1012));
  OAI21_X1  g587(.A(new_n996), .B1(new_n801), .B2(new_n991), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n1014), .B(KEYINPUT47), .Z(new_n1015));
  NAND2_X1  g590(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(G2067), .B2(new_n775), .ZN(new_n1017));
  AOI211_X1 g592(.A(new_n1011), .B(new_n1015), .C1(new_n996), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n995), .A2(new_n993), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(G1976), .B2(new_n591), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n1023));
  INV_X1    g598(.A(G288), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(G1976), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1022), .B1(new_n1025), .B2(KEYINPUT111), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(KEYINPUT111), .B2(new_n1025), .ZN(new_n1027));
  OR2_X1    g602(.A1(G305), .A2(G1981), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n600), .A2(new_n593), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G1981), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT49), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n1020), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(KEYINPUT49), .A3(new_n1030), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1032), .A2(new_n1033), .B1(KEYINPUT52), .B2(new_n1022), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G303), .A2(G8), .ZN(new_n1035));
  XOR2_X1   g610(.A(new_n1035), .B(KEYINPUT55), .Z(new_n1036));
  INV_X1    g611(.A(G8), .ZN(new_n1037));
  INV_X1    g612(.A(G1384), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n495), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(KEYINPUT50), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n993), .B1(new_n995), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G2090), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT110), .B(G1971), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n995), .A2(KEYINPUT45), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n993), .B1(new_n995), .B2(KEYINPUT45), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1037), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1027), .B(new_n1034), .C1(new_n1036), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT45), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n994), .B1(new_n1039), .B2(new_n1053), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n1054), .A2(KEYINPUT116), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(KEYINPUT116), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(new_n1047), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  INV_X1    g633(.A(G2084), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1057), .A2(new_n1058), .B1(new_n1059), .B2(new_n1043), .ZN(new_n1060));
  OR3_X1    g635(.A1(new_n1060), .A2(new_n1037), .A3(G286), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT63), .B1(new_n1052), .B2(new_n1061), .ZN(new_n1062));
  AOI211_X1 g637(.A(G1976), .B(G288), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1028), .B(KEYINPUT112), .ZN(new_n1064));
  OAI211_X1 g639(.A(G8), .B(new_n1019), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1027), .A2(new_n1034), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1036), .A2(new_n1051), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1062), .B(new_n1065), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1061), .A2(KEYINPUT63), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G286), .A2(G8), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT121), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1060), .A2(new_n1072), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1071), .A2(KEYINPUT122), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(KEYINPUT122), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1074), .B(new_n1075), .C1(new_n1037), .C2(new_n1060), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1071), .A2(KEYINPUT51), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n1037), .B2(new_n1060), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1076), .A2(KEYINPUT51), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1073), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1054), .A2(new_n786), .A3(new_n1047), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1961), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1084), .A2(G2078), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1085), .B(new_n1087), .C1(new_n1057), .C2(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1090), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1069), .B1(new_n1082), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(G171), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(KEYINPUT62), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1095));
  XNOR2_X1  g670(.A(G299), .B(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT117), .B(G1956), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1039), .B2(KEYINPUT50), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n995), .A2(KEYINPUT113), .A3(new_n1041), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1042), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1098), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1097), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1098), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(new_n1096), .A3(new_n1107), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT61), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(G1348), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n995), .A2(new_n777), .A3(new_n993), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1116), .A2(new_n623), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n623), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT60), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n623), .A2(KEYINPUT60), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1114), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1054), .A2(new_n999), .A3(new_n1047), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1054), .A2(KEYINPUT119), .A3(new_n999), .A4(new_n1047), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(KEYINPUT58), .B(G1341), .Z(new_n1130));
  NAND2_X1  g705(.A1(new_n1019), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT120), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1131), .ZN(new_n1134));
  AOI211_X1 g709(.A(new_n1133), .B(new_n1134), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n558), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(KEYINPUT59), .B(new_n558), .C1(new_n1132), .C2(new_n1135), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1109), .A2(new_n1113), .A3(KEYINPUT61), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1124), .A2(new_n1138), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1142), .A2(new_n1109), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT53), .B1(new_n1105), .B2(new_n786), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(G171), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1054), .A2(new_n1047), .A3(new_n1088), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(new_n1087), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT54), .B1(new_n1093), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1087), .A2(new_n1147), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT124), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1085), .A2(new_n1152), .A3(new_n1087), .A4(new_n1147), .ZN(new_n1153));
  AOI21_X1  g728(.A(G301), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1154), .B(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT54), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1057), .A2(new_n1089), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1158), .A2(new_n1087), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1157), .B1(new_n1159), .B2(new_n1146), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1149), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1094), .B1(new_n1144), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1092), .B1(new_n1162), .B2(new_n1082), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1066), .A2(KEYINPUT115), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1067), .B1(new_n1066), .B2(KEYINPUT115), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1110), .A2(KEYINPUT114), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1044), .B1(new_n1110), .B2(KEYINPUT114), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1050), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1036), .B1(new_n1168), .B2(G8), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1164), .A2(new_n1165), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1068), .B1(new_n1163), .B2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n722), .B(G1986), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1002), .B(new_n1005), .C1(new_n997), .C2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1018), .B1(new_n1171), .B2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g749(.A1(G227), .A2(new_n461), .ZN(new_n1176));
  OR3_X1    g750(.A1(G229), .A2(G401), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g751(.A(new_n1177), .B1(new_n902), .B2(new_n906), .ZN(new_n1178));
  NAND3_X1  g752(.A1(new_n987), .A2(new_n988), .A3(new_n1178), .ZN(G225));
  NAND2_X1  g753(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1180));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n1181));
  NAND4_X1  g755(.A1(new_n987), .A2(new_n1178), .A3(new_n1181), .A4(new_n988), .ZN(new_n1182));
  AND2_X1   g756(.A1(new_n1180), .A2(new_n1182), .ZN(G308));
endmodule


