//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n603, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n463), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n463), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT68), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n477), .A2(G2105), .ZN(new_n481));
  MUX2_X1   g056(.A(G100), .B(G112), .S(G2105), .Z(new_n482));
  AOI22_X1  g057(.A1(new_n481), .A2(G136), .B1(G2104), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .A3(G138), .ZN(new_n487));
  OR2_X1    g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(G102), .A2(G2104), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n463), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n488), .B2(new_n489), .ZN(new_n495));
  NAND2_X1  g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2105), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n463), .C1(new_n475), .C2(new_n476), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n493), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT70), .A2(G651), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n508), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n515), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  AND2_X1   g095(.A1(new_n511), .A2(new_n512), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n511), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n523), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n522), .A2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(new_n509), .A2(G52), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n513), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n517), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G171));
  AOI22_X1  g111(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n517), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n521), .A2(G81), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n509), .A2(G43), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT71), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n538), .A2(new_n543), .A3(new_n539), .A4(new_n540), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OAI211_X1 g129(.A(KEYINPUT72), .B(new_n553), .C1(new_n526), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(KEYINPUT72), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n509), .A2(G53), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n553), .A2(KEYINPUT72), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(new_n512), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(new_n521), .B2(G91), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT73), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  NAND2_X1  g144(.A1(new_n509), .A2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n570), .B(new_n571), .C1(new_n513), .C2(new_n572), .ZN(G288));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  OR3_X1    g149(.A1(new_n563), .A2(KEYINPUT74), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT74), .B1(new_n563), .B2(new_n574), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n521), .A2(G86), .B1(G48), .B2(new_n509), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n517), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT75), .Z(new_n584));
  AOI22_X1  g159(.A1(new_n521), .A2(G85), .B1(G47), .B2(new_n509), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G290));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G301), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n521), .A2(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT10), .Z(new_n590));
  NAND2_X1  g165(.A1(new_n512), .A2(G66), .ZN(new_n591));
  INV_X1    g166(.A(G79), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT76), .B1(new_n592), .B2(new_n504), .ZN(new_n593));
  OR3_X1    g168(.A1(new_n592), .A2(new_n504), .A3(KEYINPUT76), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G54), .B2(new_n509), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n588), .B1(new_n597), .B2(new_n587), .ZN(G284));
  AOI21_X1  g173(.A(new_n588), .B1(new_n597), .B2(new_n587), .ZN(G321));
  NAND2_X1  g174(.A1(G299), .A2(new_n587), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n587), .B2(G168), .ZN(G297));
  OAI21_X1  g176(.A(new_n600), .B1(new_n587), .B2(G168), .ZN(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n597), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND3_X1  g179(.A1(new_n597), .A2(new_n603), .A3(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n546), .A2(new_n587), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT11), .Z(G282));
  INV_X1    g183(.A(new_n607), .ZN(G323));
  NAND2_X1  g184(.A1(new_n481), .A2(G2104), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XOR2_X1   g186(.A(KEYINPUT77), .B(KEYINPUT13), .Z(new_n612));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n611), .A2(new_n612), .B1(new_n613), .B2(G2100), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n611), .B2(new_n612), .ZN(new_n615));
  OR3_X1    g190(.A1(new_n615), .A2(new_n613), .A3(G2100), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n613), .B2(G2100), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n481), .A2(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n478), .A2(G123), .ZN(new_n619));
  MUX2_X1   g194(.A(G99), .B(G111), .S(G2105), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G2104), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2096), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n616), .A2(new_n617), .A3(new_n624), .ZN(G156));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT15), .B(G2435), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2427), .ZN(new_n629));
  INV_X1    g204(.A(G2430), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(new_n629), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XOR2_X1   g209(.A(G2443), .B(G2446), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT79), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n632), .A2(new_n639), .ZN(new_n641));
  AND3_X1   g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT80), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n645), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n644), .A2(new_n647), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(KEYINPUT17), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(KEYINPUT17), .A3(new_n646), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n646), .B1(new_n651), .B2(KEYINPUT17), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n644), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n650), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2100), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT82), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT20), .Z(new_n669));
  NOR2_X1   g244(.A1(new_n662), .A2(new_n664), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n671), .A2(new_n667), .A3(new_n665), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n669), .B(new_n672), .C1(new_n667), .C2(new_n671), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G229));
  MUX2_X1   g254(.A(G6), .B(G305), .S(G16), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT32), .B(G1981), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  MUX2_X1   g257(.A(G23), .B(G288), .S(G16), .Z(new_n683));
  XOR2_X1   g258(.A(KEYINPUT33), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G22), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT85), .Z(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G166), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1971), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n682), .A2(new_n685), .A3(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n481), .A2(G131), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT84), .Z(new_n696));
  MUX2_X1   g271(.A(G95), .B(G107), .S(G2105), .Z(new_n697));
  AOI22_X1  g272(.A1(new_n478), .A2(G119), .B1(G2104), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G29), .ZN(new_n700));
  INV_X1    g275(.A(G25), .ZN(new_n701));
  OAI21_X1  g276(.A(KEYINPUT83), .B1(new_n701), .B2(G29), .ZN(new_n702));
  OR3_X1    g277(.A1(new_n701), .A2(KEYINPUT83), .A3(G29), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT35), .B(G1991), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(G16), .A2(G24), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G290), .B2(new_n686), .ZN(new_n709));
  INV_X1    g284(.A(G1986), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n707), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n693), .A2(new_n694), .A3(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT36), .Z(new_n715));
  NAND2_X1  g290(.A1(G299), .A2(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n686), .A2(G20), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT23), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1956), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n597), .A2(G16), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G4), .B2(G16), .ZN(new_n722));
  INV_X1    g297(.A(G1348), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G26), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  MUX2_X1   g302(.A(G104), .B(G116), .S(G2105), .Z(new_n728));
  AOI22_X1  g303(.A1(new_n478), .A2(G128), .B1(G2104), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G140), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n468), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n727), .B1(new_n734), .B2(new_n725), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT87), .B(G2067), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n722), .A2(new_n723), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n735), .A2(new_n736), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n724), .A2(new_n737), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n465), .A2(KEYINPUT25), .A3(G103), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT25), .ZN(new_n742));
  INV_X1    g317(.A(G103), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n464), .B2(new_n743), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n481), .A2(G139), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n463), .B2(new_n746), .ZN(new_n747));
  MUX2_X1   g322(.A(G33), .B(new_n747), .S(G29), .Z(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G2072), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n686), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G168), .B2(new_n686), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G1966), .ZN(new_n752));
  NAND2_X1  g327(.A1(G164), .A2(G29), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G27), .B2(G29), .ZN(new_n754));
  INV_X1    g329(.A(G2078), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n751), .A2(G1966), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n749), .A2(new_n752), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n622), .A2(new_n725), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT90), .Z(new_n760));
  XOR2_X1   g335(.A(KEYINPUT27), .B(G1996), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT88), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n725), .A2(G32), .ZN(new_n764));
  AOI22_X1  g339(.A1(G129), .A2(new_n478), .B1(new_n481), .B2(G141), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n465), .A2(G105), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT26), .Z(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n764), .B1(new_n769), .B2(G29), .ZN(new_n770));
  NAND2_X1  g345(.A1(G160), .A2(G29), .ZN(new_n771));
  AND2_X1   g346(.A1(KEYINPUT24), .A2(G34), .ZN(new_n772));
  NOR2_X1   g347(.A1(KEYINPUT24), .A2(G34), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n725), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G2084), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n763), .A2(new_n770), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n760), .B(new_n777), .C1(new_n776), .C2(new_n775), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G28), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n725), .B1(new_n779), .B2(G28), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(KEYINPUT91), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(KEYINPUT91), .B2(new_n781), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT31), .B(G11), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT89), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  OAI221_X1 g361(.A(new_n786), .B1(new_n770), .B2(new_n763), .C1(new_n754), .C2(new_n755), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n740), .A2(new_n758), .A3(new_n778), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n686), .A2(G19), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n546), .B2(new_n686), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1341), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G29), .A2(G35), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G162), .B2(G29), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT29), .Z(new_n795));
  INV_X1    g370(.A(G2090), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G5), .A2(G16), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G171), .B2(G16), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT92), .Z(new_n800));
  INV_X1    g375(.A(G1961), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT93), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n795), .A2(new_n796), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n797), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n715), .A2(new_n720), .A3(new_n792), .A4(new_n806), .ZN(G311));
  INV_X1    g382(.A(G311), .ZN(G150));
  NAND2_X1  g383(.A1(new_n509), .A2(G55), .ZN(new_n809));
  INV_X1    g384(.A(G93), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n513), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(new_n517), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G860), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT37), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n597), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n541), .A2(new_n814), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n545), .B2(new_n814), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT39), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n815), .B1(new_n824), .B2(KEYINPUT39), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n817), .B1(new_n825), .B2(new_n826), .ZN(G145));
  XNOR2_X1  g402(.A(new_n733), .B(new_n502), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n769), .B(new_n747), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n831));
  MUX2_X1   g406(.A(G106), .B(G118), .S(G2105), .Z(new_n832));
  AOI22_X1  g407(.A1(new_n478), .A2(G130), .B1(G2104), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G142), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n468), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n611), .B(new_n835), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n699), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n830), .B1(new_n831), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n831), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n484), .B(new_n622), .ZN(new_n841));
  XOR2_X1   g416(.A(G160), .B(KEYINPUT95), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT97), .ZN(new_n846));
  AOI21_X1  g421(.A(G37), .B1(new_n840), .B2(new_n844), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT40), .ZN(G395));
  NOR3_X1   g424(.A1(new_n811), .A2(new_n813), .A3(G868), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n597), .A2(new_n603), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n822), .Z(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n597), .ZN(new_n854));
  XNOR2_X1  g429(.A(G299), .B(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT98), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n855), .B(KEYINPUT41), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n853), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT101), .ZN(new_n861));
  XOR2_X1   g436(.A(G290), .B(G288), .Z(new_n862));
  XNOR2_X1  g437(.A(G303), .B(KEYINPUT99), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G305), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n864), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(KEYINPUT100), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n865), .B2(new_n866), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT42), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(KEYINPUT42), .B2(new_n867), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n861), .B(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n850), .B1(new_n873), .B2(G868), .ZN(G295));
  AOI21_X1  g449(.A(new_n850), .B1(new_n873), .B2(G868), .ZN(G331));
  OR2_X1    g450(.A1(G301), .A2(KEYINPUT102), .ZN(new_n876));
  NAND2_X1  g451(.A1(G301), .A2(KEYINPUT102), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(G286), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(G286), .B2(new_n876), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(new_n822), .Z(new_n880));
  NAND2_X1  g455(.A1(new_n858), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n880), .A2(new_n855), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n868), .A2(new_n870), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT103), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT103), .B1(new_n883), .B2(new_n884), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n883), .A2(new_n884), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT43), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(G37), .B1(new_n883), .B2(new_n884), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n884), .B2(new_n883), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n887), .B2(new_n890), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n893), .A2(KEYINPUT43), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  MUX2_X1   g474(.A(new_n896), .B(new_n899), .S(KEYINPUT44), .Z(G397));
  INV_X1    g475(.A(G1384), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n486), .A2(KEYINPUT4), .A3(G138), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n492), .B1(new_n467), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n501), .B1(new_n903), .B2(G2105), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n467), .A2(G126), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n463), .B1(new_n905), .B2(new_n496), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n901), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n471), .A2(new_n472), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(G2105), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n481), .A2(G137), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n911), .A2(G40), .A3(new_n466), .A4(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT104), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(G1996), .A3(new_n769), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n733), .B(G2067), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n915), .ZN(new_n918));
  INV_X1    g493(.A(G1996), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n920), .A2(new_n769), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n916), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n699), .A2(new_n706), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(G2067), .B2(new_n733), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n915), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n920), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(new_n915), .B2(new_n769), .ZN(new_n931));
  NOR2_X1   g506(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n929), .B1(new_n920), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n931), .A2(new_n918), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT47), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n705), .B1(new_n696), .B2(new_n698), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n915), .B1(new_n936), .B2(new_n923), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n922), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n914), .A2(new_n710), .A3(new_n584), .A4(new_n585), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n939), .B(KEYINPUT126), .Z(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT48), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n928), .B(new_n935), .C1(new_n938), .C2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT127), .ZN(new_n943));
  INV_X1    g518(.A(G1981), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n579), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(G305), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT49), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n491), .B1(new_n477), .B2(new_n487), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n951), .A2(new_n463), .B1(new_n500), .B2(new_n499), .ZN(new_n952));
  AOI21_X1  g527(.A(G1384), .B1(new_n952), .B2(new_n498), .ZN(new_n953));
  INV_X1    g528(.A(G40), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n470), .A2(new_n473), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(G8), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n949), .A2(new_n950), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G1976), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT52), .B1(G288), .B2(new_n959), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n956), .B(G8), .C1(new_n959), .C2(G288), .ZN(new_n961));
  MUX2_X1   g536(.A(new_n960), .B(KEYINPUT52), .S(new_n961), .Z(new_n962));
  NOR2_X1   g537(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n955), .B1(new_n907), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT106), .B1(new_n953), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n907), .A2(new_n969), .A3(KEYINPUT50), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n966), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n796), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n972), .A2(KEYINPUT107), .ZN(new_n973));
  OAI211_X1 g548(.A(KEYINPUT45), .B(new_n901), .C1(new_n904), .C2(new_n906), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n909), .A2(new_n955), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1971), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n972), .B2(KEYINPUT107), .ZN(new_n978));
  OAI21_X1  g553(.A(G8), .B1(new_n973), .B2(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(G303), .B(G8), .C1(KEYINPUT108), .C2(KEYINPUT55), .ZN(new_n980));
  NAND2_X1  g555(.A1(KEYINPUT108), .A2(KEYINPUT55), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n980), .B(new_n981), .Z(new_n982));
  OR2_X1    g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n963), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n977), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n955), .B1(new_n907), .B2(KEYINPUT50), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n964), .B1(new_n502), .B2(new_n901), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n986), .A2(G2090), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(G8), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n982), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n984), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n909), .A2(new_n755), .A3(new_n955), .A4(new_n974), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n974), .B(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT45), .B1(new_n502), .B2(new_n901), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(new_n999), .B2(new_n913), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT111), .B(new_n955), .C1(new_n953), .C2(KEYINPUT45), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n994), .A2(G2078), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n997), .A2(new_n1000), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n913), .B1(new_n953), .B2(new_n964), .ZN(new_n1004));
  AOI211_X1 g579(.A(KEYINPUT106), .B(new_n967), .C1(new_n502), .C2(new_n901), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n969), .B1(new_n907), .B2(KEYINPUT50), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n801), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1003), .A2(new_n1008), .A3(KEYINPUT120), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT120), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1010));
  OAI211_X1 g585(.A(G301), .B(new_n995), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT121), .B1(new_n971), .B2(G1961), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1007), .A2(new_n1014), .A3(new_n801), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n993), .A2(new_n994), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1013), .A2(new_n1015), .A3(new_n995), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1012), .B1(new_n1017), .B2(G171), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1011), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT122), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1011), .A2(new_n1018), .A3(KEYINPUT122), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1024));
  AOI21_X1  g599(.A(G301), .B1(new_n1024), .B2(new_n995), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1017), .A2(G171), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1012), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  INV_X1    g605(.A(G1966), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n974), .A2(KEYINPUT112), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n953), .A2(new_n996), .A3(KEYINPUT45), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1000), .A2(new_n1001), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT113), .B(G2084), .Z(new_n1035));
  OAI211_X1 g610(.A(new_n1004), .B(new_n1035), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1031), .A2(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n971), .A2(KEYINPUT114), .A3(new_n1035), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1030), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G286), .A2(G8), .ZN(new_n1041));
  XOR2_X1   g616(.A(new_n1041), .B(KEYINPUT118), .Z(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1029), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1034), .A2(new_n1031), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(new_n1039), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G8), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(KEYINPUT51), .A3(new_n1042), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1042), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AND4_X1   g626(.A1(new_n1028), .A2(new_n1044), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1043), .B1(new_n1047), .B2(G8), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1050), .B1(new_n1053), .B2(KEYINPUT51), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1028), .B1(new_n1054), .B2(new_n1044), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1023), .B(new_n1027), .C1(new_n1052), .C2(new_n1055), .ZN(new_n1056));
  OAI22_X1  g631(.A1(new_n971), .A2(G1348), .B1(G2067), .B2(new_n956), .ZN(new_n1057));
  INV_X1    g632(.A(G1956), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n986), .B2(new_n987), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n561), .A2(KEYINPUT57), .A3(new_n566), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n565), .A2(G651), .ZN(new_n1062));
  INV_X1    g637(.A(G91), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1062), .B1(new_n1063), .B2(new_n513), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n559), .B1(new_n555), .B2(new_n557), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1061), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1060), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n909), .A2(new_n955), .A3(new_n974), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1059), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1057), .A2(new_n597), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1059), .A2(new_n1069), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1067), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1074), .A2(KEYINPUT61), .A3(new_n1070), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT61), .B1(new_n1074), .B2(new_n1070), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n909), .A2(new_n919), .A3(new_n955), .A4(new_n974), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n956), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n546), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT116), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1082), .A2(new_n1086), .A3(new_n546), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  AOI211_X1 g663(.A(KEYINPUT116), .B(new_n545), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1086), .B1(new_n1082), .B2(new_n546), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT59), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1078), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT117), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1078), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1057), .A2(KEYINPUT60), .A3(new_n854), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1057), .B(new_n597), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(KEYINPUT60), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1075), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1056), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1025), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1053), .A2(KEYINPUT51), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT119), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1054), .A2(new_n1028), .A3(new_n1044), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(KEYINPUT62), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1103), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n992), .B1(new_n1102), .B2(new_n1111), .ZN(new_n1112));
  XOR2_X1   g687(.A(new_n957), .B(KEYINPUT110), .Z(new_n1113));
  NOR3_X1   g688(.A1(new_n958), .A2(G1976), .A3(G288), .ZN(new_n1114));
  NOR2_X1   g689(.A1(G305), .A2(G1981), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n963), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1116), .B1(new_n983), .B2(new_n1117), .ZN(new_n1118));
  XOR2_X1   g693(.A(KEYINPUT115), .B(KEYINPUT63), .Z(new_n1119));
  NOR2_X1   g694(.A1(new_n1048), .A2(G286), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n991), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n979), .A2(new_n982), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n984), .A2(KEYINPUT63), .A3(new_n1120), .A4(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1118), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1112), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(G290), .B(new_n710), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n938), .B1(new_n914), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT123), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1129), .ZN(new_n1132));
  AOI211_X1 g707(.A(new_n1131), .B(new_n1132), .C1(new_n1112), .C2(new_n1125), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n943), .B1(new_n1130), .B2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g709(.A1(G229), .A2(G227), .A3(new_n461), .A4(G401), .ZN(new_n1136));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n848), .A3(new_n1136), .ZN(G225));
  INV_X1    g711(.A(G225), .ZN(G308));
endmodule


