//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n205));
  OAI221_X1 g004(.A(new_n203), .B1(KEYINPUT92), .B2(G8gat), .C1(new_n202), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n206), .B(new_n207), .Z(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT14), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n211), .A2(KEYINPUT91), .ZN(new_n212));
  NAND2_X1  g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(new_n211), .B2(KEYINPUT91), .ZN(new_n214));
  OAI211_X1 g013(.A(KEYINPUT15), .B(new_n209), .C1(new_n212), .C2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(new_n211), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n218), .A3(new_n213), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n208), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G229gat), .A2(G233gat), .ZN(new_n223));
  XOR2_X1   g022(.A(new_n223), .B(KEYINPUT13), .Z(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(new_n225), .B(KEYINPUT94), .Z(new_n226));
  NOR2_X1   g025(.A1(new_n208), .A2(new_n221), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n228), .A2(new_n208), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n227), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n223), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT18), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n226), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT93), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n232), .A2(new_n233), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G113gat), .B(G141gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(G197gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT11), .B(G169gat), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g041(.A(new_n242), .B(KEYINPUT12), .Z(new_n243));
  NAND3_X1  g042(.A1(new_n236), .A2(new_n238), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n243), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n235), .B(new_n237), .C1(KEYINPUT93), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT36), .ZN(new_n249));
  NAND2_X1  g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n251));
  INV_X1    g050(.A(G169gat), .ZN(new_n252));
  INV_X1    g051(.A(G176gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n258));
  AOI22_X1  g057(.A1(KEYINPUT26), .A2(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n254), .A2(KEYINPUT26), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n263));
  INV_X1    g062(.A(G183gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(KEYINPUT27), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT27), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(G183gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n263), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(G183gat), .ZN(new_n269));
  AOI21_X1  g068(.A(G190gat), .B1(new_n269), .B2(KEYINPUT68), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n262), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(KEYINPUT27), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G190gat), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n274), .A2(KEYINPUT28), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n250), .B(new_n261), .C1(new_n271), .C2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278));
  AND2_X1   g077(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(G190gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n250), .A2(KEYINPUT64), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT64), .B1(new_n250), .B2(new_n281), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n280), .B(KEYINPUT65), .C1(new_n282), .C2(new_n283), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n252), .A3(new_n253), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n257), .A2(new_n258), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT25), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n286), .A2(new_n287), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G127gat), .B(G134gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(G113gat), .A2(G120gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(G113gat), .A2(G120gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT1), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n296), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G113gat), .ZN(new_n303));
  INV_X1    g102(.A(G120gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT71), .B1(new_n305), .B2(new_n297), .ZN(new_n306));
  OR2_X1    g105(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n307));
  NAND2_X1  g106(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G134gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G127gat), .ZN(new_n311));
  INV_X1    g110(.A(G127gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G134gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n306), .A2(new_n309), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT71), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n302), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n278), .ZN(new_n318));
  NAND3_X1  g117(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT67), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n318), .B(new_n319), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n320), .A2(new_n321), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n292), .B(new_n291), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT25), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n277), .A2(new_n295), .A3(new_n317), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT73), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n273), .A2(new_n275), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT68), .B1(new_n269), .B2(new_n272), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT68), .B1(new_n264), .B2(KEYINPUT27), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n274), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n328), .B1(new_n332), .B2(new_n262), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n259), .A2(new_n260), .B1(G183gat), .B2(G190gat), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n333), .A2(new_n334), .B1(KEYINPUT25), .B2(new_n324), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n317), .A4(new_n295), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n277), .A2(new_n295), .A3(new_n325), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n309), .A2(new_n314), .ZN(new_n339));
  INV_X1    g138(.A(new_n306), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n340), .A3(new_n316), .ZN(new_n341));
  INV_X1    g140(.A(new_n302), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n337), .A3(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n345), .A2(KEYINPUT74), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT74), .B1(new_n345), .B2(new_n346), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT32), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT33), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(new_n347), .B2(new_n348), .ZN(new_n351));
  XOR2_X1   g150(.A(G15gat), .B(G43gat), .Z(new_n352));
  XNOR2_X1  g151(.A(G71gat), .B(G99gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n349), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n354), .ZN(new_n356));
  OAI221_X1 g155(.A(KEYINPUT32), .B1(new_n350), .B2(new_n356), .C1(new_n347), .C2(new_n348), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n345), .A2(new_n346), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT34), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n359), .B(KEYINPUT34), .Z(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(new_n355), .A3(new_n357), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n249), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(KEYINPUT75), .A3(new_n363), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n358), .A2(new_n366), .A3(new_n360), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n364), .B1(new_n368), .B2(new_n249), .ZN(new_n369));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT82), .ZN(new_n371));
  NAND2_X1  g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372));
  INV_X1    g171(.A(G155gat), .ZN(new_n373));
  INV_X1    g172(.A(G162gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G141gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(G148gat), .ZN(new_n377));
  INV_X1    g176(.A(G148gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G141gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n372), .B(new_n375), .C1(new_n380), .C2(KEYINPUT2), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n372), .B1(new_n375), .B2(KEYINPUT2), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(new_n376), .B2(G148gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(G141gat), .B2(new_n378), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n383), .A2(new_n376), .A3(G148gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(G197gat), .A2(G204gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(G197gat), .A2(G204gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G211gat), .A2(G218gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI22_X1  g193(.A1(new_n390), .A2(new_n392), .B1(new_n394), .B2(KEYINPUT22), .ZN(new_n395));
  NOR2_X1   g194(.A1(G211gat), .A2(G218gat), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n394), .A2(new_n396), .A3(KEYINPUT76), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT76), .ZN(new_n398));
  INV_X1    g197(.A(G211gat), .ZN(new_n399));
  INV_X1    g198(.A(G218gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n398), .B1(new_n401), .B2(new_n393), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n395), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  OR2_X1    g203(.A1(G197gat), .A2(G204gat), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT22), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n405), .A2(new_n391), .B1(new_n406), .B2(new_n393), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT76), .B1(new_n394), .B2(new_n396), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n401), .A2(new_n398), .A3(new_n393), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n403), .A2(new_n404), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT3), .B1(new_n411), .B2(KEYINPUT83), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n403), .A2(new_n413), .A3(new_n410), .A4(new_n404), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n389), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n403), .A2(new_n410), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT77), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n403), .A2(KEYINPUT77), .A3(new_n410), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT3), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n381), .A2(new_n387), .A3(new_n420), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n418), .A2(new_n419), .B1(new_n404), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n371), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n404), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n418), .A2(new_n419), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n421), .A2(KEYINPUT84), .A3(new_n404), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n388), .A2(KEYINPUT3), .ZN(new_n430));
  INV_X1    g229(.A(new_n370), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n389), .A2(new_n411), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(G22gat), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n423), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n423), .B2(new_n435), .ZN(new_n438));
  OAI21_X1  g237(.A(G78gat), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n435), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G22gat), .ZN(new_n441));
  INV_X1    g240(.A(G78gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n435), .A3(new_n436), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT31), .B(G50gat), .ZN(new_n445));
  INV_X1    g244(.A(G106gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n439), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n439), .B2(new_n444), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n343), .B(new_n388), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G225gat), .A2(G233gat), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT79), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n430), .A2(new_n343), .A3(new_n421), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n389), .A2(new_n317), .A3(KEYINPUT4), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n343), .B2(new_n388), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n455), .A2(new_n456), .A3(new_n458), .A4(new_n453), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT79), .ZN(new_n460));
  INV_X1    g259(.A(new_n453), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n451), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n454), .A2(KEYINPUT5), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n455), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(new_n461), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT5), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT81), .B1(new_n456), .B2(new_n458), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n456), .A2(new_n458), .A3(KEYINPUT81), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n465), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(G1gat), .B(G29gat), .Z(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G57gat), .B(G85gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477));
  INV_X1    g276(.A(new_n475), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n478), .A3(new_n469), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n470), .A2(KEYINPUT6), .A3(new_n475), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(G226gat), .A2(G233gat), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(KEYINPUT29), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n338), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(new_n338), .B2(new_n483), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n487), .A2(new_n427), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n427), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G8gat), .B(G36gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(G64gat), .B(G92gat), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n491), .B(new_n492), .Z(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n488), .A2(new_n489), .A3(new_n493), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(KEYINPUT30), .A3(new_n496), .ZN(new_n497));
  OR3_X1    g296(.A1(new_n490), .A2(KEYINPUT30), .A3(new_n494), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n450), .B1(new_n482), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT85), .B1(new_n369), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT36), .B1(new_n365), .B2(new_n367), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n505));
  NOR4_X1   g304(.A1(new_n504), .A2(new_n505), .A3(new_n500), .A4(new_n364), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n482), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n496), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n495), .B1(new_n510), .B2(new_n493), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n487), .A2(KEYINPUT87), .A3(new_n427), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT37), .B(new_n512), .C1(new_n490), .C2(KEYINPUT87), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT38), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT38), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n515), .B1(new_n490), .B2(KEYINPUT37), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n514), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n450), .B1(new_n509), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n499), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT39), .B1(new_n451), .B2(new_n461), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n455), .B1(new_n468), .B2(new_n467), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(new_n461), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT39), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n524), .A3(new_n461), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n523), .A2(new_n478), .A3(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n519), .B(new_n476), .C1(new_n526), .C2(KEYINPUT40), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n523), .A2(KEYINPUT40), .A3(new_n478), .A4(new_n525), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT86), .Z(new_n529));
  NOR2_X1   g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n518), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n503), .A2(new_n507), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n482), .A2(new_n499), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n450), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(KEYINPUT35), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n368), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n361), .A2(new_n450), .A3(new_n363), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT89), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n534), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n361), .A2(new_n450), .A3(KEYINPUT89), .A4(new_n363), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n545), .A2(KEYINPUT90), .A3(KEYINPUT35), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT90), .B1(new_n545), .B2(KEYINPUT35), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n539), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n248), .B1(new_n533), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT7), .ZN(new_n551));
  NAND2_X1  g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552));
  INV_X1    g351(.A(G85gat), .ZN(new_n553));
  INV_X1    g352(.A(G92gat), .ZN(new_n554));
  AOI22_X1  g353(.A1(KEYINPUT8), .A2(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G99gat), .B(G106gat), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT97), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n556), .A2(new_n557), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n228), .A2(new_n230), .A3(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n562), .B(KEYINPUT98), .Z(new_n563));
  INV_X1    g362(.A(KEYINPUT41), .ZN(new_n564));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565));
  OAI221_X1 g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .C1(new_n221), .C2(new_n561), .ZN(new_n566));
  XOR2_X1   g365(.A(G190gat), .B(G218gat), .Z(new_n567));
  OR2_X1    g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n564), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT96), .ZN(new_n572));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT99), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n574), .B(KEYINPUT99), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n568), .A2(new_n569), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G57gat), .B(G64gat), .Z(new_n580));
  INV_X1    g379(.A(G71gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(new_n442), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(KEYINPUT9), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G71gat), .B(G78gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(new_n312), .ZN(new_n589));
  XOR2_X1   g388(.A(G183gat), .B(G211gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT21), .ZN(new_n592));
  INV_X1    g391(.A(new_n585), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n208), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT95), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(new_n373), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n595), .B(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n591), .A2(new_n598), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n579), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n561), .A2(new_n593), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n560), .A3(new_n558), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n585), .A2(KEYINPUT10), .ZN(new_n607));
  OAI22_X1  g406(.A1(new_n606), .A2(KEYINPUT10), .B1(new_n561), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G230gat), .ZN(new_n609));
  INV_X1    g408(.A(G233gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n606), .A2(new_n611), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G120gat), .B(G148gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT100), .ZN(new_n617));
  XOR2_X1   g416(.A(G176gat), .B(G204gat), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n615), .B(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n620), .A2(KEYINPUT101), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(KEYINPUT101), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n603), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n549), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(new_n482), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n204), .ZN(G1324gat));
  NAND3_X1  g426(.A1(new_n549), .A2(new_n519), .A3(new_n624), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n628), .A2(G8gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT16), .B(G8gat), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT42), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n632), .B1(KEYINPUT42), .B2(new_n631), .ZN(G1325gat));
  OAI21_X1  g432(.A(G15gat), .B1(new_n625), .B2(new_n369), .ZN(new_n634));
  INV_X1    g433(.A(new_n368), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n635), .A2(G15gat), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n625), .B2(new_n636), .ZN(G1326gat));
  NOR2_X1   g436(.A1(new_n625), .A2(new_n450), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT43), .B(G22gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(G1327gat));
  INV_X1    g439(.A(G29gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n576), .A2(new_n578), .ZN(new_n642));
  INV_X1    g441(.A(new_n539), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n545), .A2(KEYINPUT35), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT90), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n545), .A2(KEYINPUT90), .A3(KEYINPUT35), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n369), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n649), .A2(new_n531), .A3(new_n500), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n642), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n533), .A2(new_n548), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n579), .A2(new_n652), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n651), .A2(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n248), .A2(new_n602), .A3(new_n623), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n482), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n641), .B1(new_n659), .B2(KEYINPUT102), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(KEYINPUT102), .B2(new_n659), .ZN(new_n661));
  INV_X1    g460(.A(new_n623), .ZN(new_n662));
  AND4_X1   g461(.A1(new_n549), .A2(new_n601), .A3(new_n642), .A4(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n641), .A3(new_n508), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT45), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n665), .ZN(G1328gat));
  AOI21_X1  g465(.A(G36gat), .B1(KEYINPUT103), .B2(KEYINPUT46), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n519), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(G36gat), .B1(new_n657), .B2(new_n499), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(G1329gat));
  OAI21_X1  g471(.A(G43gat), .B1(new_n657), .B2(new_n369), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n635), .A2(G43gat), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT47), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n663), .A2(new_n674), .B1(KEYINPUT104), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n675), .A2(KEYINPUT104), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n677), .B(new_n678), .Z(G1330gat));
  NAND3_X1  g478(.A1(new_n655), .A2(new_n537), .A3(new_n656), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n450), .A2(G50gat), .ZN(new_n681));
  AOI22_X1  g480(.A1(new_n680), .A2(G50gat), .B1(new_n663), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g482(.A1(new_n248), .A2(new_n623), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n532), .A2(new_n501), .A3(new_n369), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n684), .B(new_n603), .C1(new_n548), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n508), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G57gat), .ZN(G1332gat));
  INV_X1    g487(.A(KEYINPUT49), .ZN(new_n689));
  INV_X1    g488(.A(G64gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n519), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT105), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1333gat));
  AOI21_X1  g494(.A(new_n581), .B1(new_n686), .B2(new_n649), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n635), .A2(G71gat), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n686), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g498(.A1(new_n686), .A2(new_n537), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(G78gat), .ZN(G1335gat));
  INV_X1    g500(.A(KEYINPUT51), .ZN(new_n702));
  OAI211_X1 g501(.A(KEYINPUT107), .B(new_n642), .C1(new_n648), .C2(new_n650), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n248), .A2(new_n601), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n579), .B1(new_n548), .B2(new_n685), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(KEYINPUT107), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n702), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n651), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n711), .A2(KEYINPUT51), .A3(new_n705), .A4(new_n703), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n662), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(new_n553), .A3(new_n508), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n502), .A2(new_n506), .A3(new_n531), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n654), .B1(new_n648), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n704), .A2(new_n662), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n716), .B(new_n717), .C1(new_n707), .C2(KEYINPUT44), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n651), .A2(new_n652), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n721), .A2(KEYINPUT106), .A3(new_n716), .A4(new_n717), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G85gat), .B1(new_n723), .B2(new_n482), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n714), .A2(new_n724), .ZN(G1336gat));
  NAND3_X1  g524(.A1(new_n713), .A2(new_n554), .A3(new_n519), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727));
  OAI21_X1  g526(.A(G92gat), .B1(new_n718), .B2(new_n499), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(G92gat), .B1(new_n723), .B2(new_n499), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n731), .B2(new_n727), .ZN(G1337gat));
  INV_X1    g531(.A(G99gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n713), .A2(new_n733), .A3(new_n368), .ZN(new_n734));
  OAI21_X1  g533(.A(G99gat), .B1(new_n723), .B2(new_n369), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1338gat));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n709), .A2(new_n712), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n623), .A2(new_n446), .A3(new_n537), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT109), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n718), .B2(new_n450), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n655), .A2(KEYINPUT110), .A3(new_n537), .A4(new_n717), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n745), .A3(G106gat), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n747));
  AND4_X1   g546(.A1(KEYINPUT111), .A2(new_n742), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT53), .B1(new_n738), .B2(new_n741), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT111), .B1(new_n749), .B2(new_n746), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n740), .B1(new_n709), .B2(new_n712), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n720), .A2(new_n537), .A3(new_n722), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G106gat), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n753), .A2(KEYINPUT108), .A3(G106gat), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n747), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n737), .B1(new_n751), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n754), .A2(new_n755), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n757), .A3(new_n742), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT53), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n742), .A2(new_n746), .A3(new_n747), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n749), .A2(KEYINPUT111), .A3(new_n746), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n762), .A2(KEYINPUT112), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n759), .A2(new_n768), .ZN(G1339gat));
  INV_X1    g568(.A(new_n242), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n231), .A2(new_n223), .ZN(new_n771));
  OR2_X1    g570(.A1(new_n222), .A2(new_n224), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n238), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n245), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n623), .ZN(new_n776));
  INV_X1    g575(.A(new_n613), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n612), .B2(new_n608), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n619), .B1(new_n777), .B2(new_n778), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n782), .A2(KEYINPUT55), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n780), .A2(KEYINPUT55), .A3(new_n781), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n776), .B1(new_n248), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n579), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n642), .A2(new_n775), .A3(new_n787), .A4(new_n783), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n602), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n603), .A2(new_n247), .A3(new_n623), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OR3_X1    g593(.A1(new_n794), .A2(KEYINPUT113), .A3(new_n537), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT113), .B1(new_n794), .B2(new_n537), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n635), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n519), .A2(new_n482), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n799), .A2(new_n303), .A3(new_n248), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n794), .A2(new_n482), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n542), .A2(new_n544), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n801), .A2(new_n499), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(G113gat), .B1(new_n803), .B2(new_n247), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n800), .A2(new_n804), .ZN(G1340gat));
  NAND3_X1  g604(.A1(new_n797), .A2(new_n623), .A3(new_n798), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n662), .A2(G120gat), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n806), .A2(G120gat), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT114), .ZN(G1341gat));
  OAI21_X1  g608(.A(G127gat), .B1(new_n799), .B2(new_n601), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n803), .A2(new_n312), .A3(new_n602), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(G1342gat));
  NAND3_X1  g611(.A1(new_n803), .A2(new_n310), .A3(new_n642), .ZN(new_n813));
  XOR2_X1   g612(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n814));
  XNOR2_X1  g613(.A(new_n813), .B(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G134gat), .B1(new_n799), .B2(new_n579), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1343gat));
  NOR3_X1   g616(.A1(new_n794), .A2(new_n482), .A3(new_n519), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(new_n649), .B2(new_n450), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n369), .A2(KEYINPUT119), .A3(new_n537), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n822), .A2(G141gat), .A3(new_n248), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(KEYINPUT58), .ZN(new_n824));
  XNOR2_X1  g623(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n782), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n786), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n828), .A2(new_n247), .B1(new_n775), .B2(new_n623), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n579), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n247), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n830), .A3(new_n776), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n791), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n601), .ZN(new_n836));
  INV_X1    g635(.A(new_n793), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n537), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT57), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n369), .A2(new_n798), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n794), .A2(new_n450), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G141gat), .B1(new_n845), .B2(new_n248), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n824), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n840), .A2(new_n844), .A3(KEYINPUT118), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n247), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n823), .B1(new_n851), .B2(G141gat), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n847), .B1(new_n852), .B2(new_n853), .ZN(G1344gat));
  NOR2_X1   g653(.A1(new_n378), .A2(KEYINPUT59), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n849), .A2(new_n850), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n662), .ZN(new_n857));
  XNOR2_X1  g656(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT57), .B(new_n537), .C1(new_n792), .C2(new_n793), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n450), .B1(new_n836), .B2(new_n837), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(KEYINPUT57), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(new_n662), .A3(new_n841), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n858), .B1(new_n863), .B2(new_n378), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n822), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n378), .A3(new_n623), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1345gat));
  NAND4_X1  g667(.A1(new_n849), .A2(G155gat), .A3(new_n850), .A4(new_n602), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n373), .B1(new_n822), .B2(new_n601), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n869), .A2(KEYINPUT121), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1346gat));
  OAI21_X1  g674(.A(G162gat), .B1(new_n856), .B2(new_n579), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n866), .A2(new_n374), .A3(new_n642), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n508), .A2(new_n499), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n802), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n794), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(G169gat), .B1(new_n881), .B2(new_n247), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n797), .A2(new_n879), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n248), .A2(new_n252), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(G1348gat));
  NAND3_X1  g684(.A1(new_n881), .A2(new_n253), .A3(new_n623), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n883), .A2(new_n623), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n253), .ZN(G1349gat));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(KEYINPUT60), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(KEYINPUT60), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n797), .A2(new_n602), .A3(new_n879), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G183gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n881), .A2(new_n273), .A3(new_n602), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n890), .B(new_n891), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  AND4_X1   g694(.A1(new_n889), .A2(new_n893), .A3(KEYINPUT60), .A4(new_n894), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(G1350gat));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n274), .A3(new_n642), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n642), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(G190gat), .ZN(new_n901));
  AOI211_X1 g700(.A(KEYINPUT61), .B(new_n274), .C1(new_n883), .C2(new_n642), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(G1351gat));
  AND2_X1   g702(.A1(new_n369), .A2(new_n879), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n842), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g704(.A(KEYINPUT123), .B(G197gat), .Z(new_n906));
  OR3_X1    g705(.A1(new_n905), .A2(new_n248), .A3(new_n906), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n904), .B(KEYINPUT124), .Z(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n862), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n911), .A3(new_n247), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n906), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n911), .B1(new_n910), .B2(new_n247), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n907), .B1(new_n913), .B2(new_n914), .ZN(G1352gat));
  NOR3_X1   g714(.A1(new_n905), .A2(G204gat), .A3(new_n662), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT62), .ZN(new_n923));
  INV_X1    g722(.A(G204gat), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n862), .A2(new_n662), .A3(new_n909), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n922), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(G1353gat));
  INV_X1    g725(.A(new_n905), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n399), .A3(new_n602), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n861), .A2(new_n602), .A3(new_n908), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT63), .B1(new_n929), .B2(G211gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g733(.A(KEYINPUT127), .B(new_n928), .C1(new_n930), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1354gat));
  NAND3_X1  g735(.A1(new_n927), .A2(new_n400), .A3(new_n642), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n862), .A2(new_n579), .A3(new_n909), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n400), .ZN(G1355gat));
endmodule


