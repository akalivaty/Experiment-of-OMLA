

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U553 ( .A1(n762), .A2(n755), .ZN(n519) );
  NOR2_X1 U554 ( .A1(n975), .A2(n692), .ZN(n701) );
  XNOR2_X1 U555 ( .A(n700), .B(n699), .ZN(n703) );
  OR2_X1 U556 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U557 ( .A1(n519), .A2(n972), .ZN(n756) );
  NAND2_X1 U558 ( .A1(n674), .A2(G40), .ZN(n679) );
  XOR2_X1 U559 ( .A(KEYINPUT17), .B(n526), .Z(n881) );
  NOR2_X1 U560 ( .A1(G651), .A2(n616), .ZN(n632) );
  NOR2_X1 U561 ( .A1(n530), .A2(n529), .ZN(n674) );
  BUF_X1 U562 ( .A(n674), .Z(G160) );
  INV_X1 U563 ( .A(G2104), .ZN(n522) );
  NOR2_X4 U564 ( .A1(G2105), .A2(n522), .ZN(n880) );
  NAND2_X1 U565 ( .A1(G101), .A2(n880), .ZN(n520) );
  XOR2_X1 U566 ( .A(n520), .B(KEYINPUT23), .Z(n521) );
  XNOR2_X1 U567 ( .A(n521), .B(KEYINPUT66), .ZN(n524) );
  AND2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n876) );
  NAND2_X1 U569 ( .A1(G113), .A2(n876), .ZN(n523) );
  NAND2_X1 U570 ( .A1(n524), .A2(n523), .ZN(n530) );
  NAND2_X1 U571 ( .A1(n522), .A2(G2105), .ZN(n525) );
  XNOR2_X1 U572 ( .A(n525), .B(KEYINPUT65), .ZN(n875) );
  NAND2_X1 U573 ( .A1(G125), .A2(n875), .ZN(n528) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  NAND2_X1 U575 ( .A1(G137), .A2(n881), .ZN(n527) );
  NAND2_X1 U576 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U577 ( .A1(G651), .A2(G543), .ZN(n635) );
  NAND2_X1 U578 ( .A1(G85), .A2(n635), .ZN(n532) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n616) );
  INV_X1 U580 ( .A(G651), .ZN(n533) );
  NOR2_X1 U581 ( .A1(n616), .A2(n533), .ZN(n629) );
  NAND2_X1 U582 ( .A1(G72), .A2(n629), .ZN(n531) );
  NAND2_X1 U583 ( .A1(n532), .A2(n531), .ZN(n538) );
  NOR2_X1 U584 ( .A1(G543), .A2(n533), .ZN(n534) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n534), .Z(n631) );
  NAND2_X1 U586 ( .A1(G60), .A2(n631), .ZN(n536) );
  NAND2_X1 U587 ( .A1(G47), .A2(n632), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n537) );
  OR2_X1 U589 ( .A1(n538), .A2(n537), .ZN(G290) );
  NAND2_X1 U590 ( .A1(G90), .A2(n635), .ZN(n540) );
  NAND2_X1 U591 ( .A1(G77), .A2(n629), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U593 ( .A(n541), .B(KEYINPUT9), .ZN(n543) );
  NAND2_X1 U594 ( .A1(G52), .A2(n632), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n543), .A2(n542), .ZN(n546) );
  NAND2_X1 U596 ( .A1(G64), .A2(n631), .ZN(n544) );
  XNOR2_X1 U597 ( .A(KEYINPUT67), .B(n544), .ZN(n545) );
  NOR2_X1 U598 ( .A1(n546), .A2(n545), .ZN(G171) );
  AND2_X1 U599 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U600 ( .A1(G99), .A2(n880), .ZN(n548) );
  NAND2_X1 U601 ( .A1(G111), .A2(n876), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U603 ( .A1(n875), .A2(G123), .ZN(n549) );
  XOR2_X1 U604 ( .A(KEYINPUT18), .B(n549), .Z(n550) );
  NOR2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n553) );
  NAND2_X1 U606 ( .A1(n881), .A2(G135), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n553), .A2(n552), .ZN(n923) );
  XNOR2_X1 U608 ( .A(G2096), .B(n923), .ZN(n554) );
  OR2_X1 U609 ( .A1(G2100), .A2(n554), .ZN(G156) );
  INV_X1 U610 ( .A(G57), .ZN(G237) );
  INV_X1 U611 ( .A(G69), .ZN(G235) );
  INV_X1 U612 ( .A(G108), .ZN(G238) );
  INV_X1 U613 ( .A(G120), .ZN(G236) );
  XNOR2_X1 U614 ( .A(KEYINPUT6), .B(KEYINPUT72), .ZN(n558) );
  NAND2_X1 U615 ( .A1(G63), .A2(n631), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G51), .A2(n632), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n558), .B(n557), .ZN(n564) );
  NAND2_X1 U619 ( .A1(n635), .A2(G89), .ZN(n559) );
  XNOR2_X1 U620 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U621 ( .A1(G76), .A2(n629), .ZN(n560) );
  NAND2_X1 U622 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U623 ( .A(KEYINPUT5), .B(n562), .Z(n563) );
  NOR2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n566) );
  XNOR2_X1 U625 ( .A(KEYINPUT7), .B(KEYINPUT73), .ZN(n565) );
  XNOR2_X1 U626 ( .A(n566), .B(n565), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U629 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U630 ( .A(G223), .ZN(n823) );
  NAND2_X1 U631 ( .A1(n823), .A2(G567), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  NAND2_X1 U633 ( .A1(G56), .A2(n631), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT14), .B(n569), .Z(n576) );
  NAND2_X1 U635 ( .A1(G81), .A2(n635), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT69), .B(n570), .Z(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G68), .A2(n629), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT13), .B(n574), .Z(n575) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n632), .A2(G43), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n975) );
  INV_X1 U644 ( .A(G860), .ZN(n604) );
  OR2_X1 U645 ( .A1(n975), .A2(n604), .ZN(G153) );
  XOR2_X1 U646 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U648 ( .A1(G79), .A2(n629), .ZN(n580) );
  NAND2_X1 U649 ( .A1(G54), .A2(n632), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G66), .A2(n631), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G92), .A2(n635), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U654 ( .A(KEYINPUT71), .B(n583), .Z(n584) );
  NOR2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U656 ( .A(KEYINPUT15), .B(n586), .Z(n990) );
  OR2_X1 U657 ( .A1(n990), .A2(G868), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U659 ( .A1(G65), .A2(n631), .ZN(n590) );
  NAND2_X1 U660 ( .A1(G78), .A2(n629), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U662 ( .A1(n635), .A2(G91), .ZN(n591) );
  XOR2_X1 U663 ( .A(KEYINPUT68), .B(n591), .Z(n592) );
  NOR2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n632), .A2(G53), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(G299) );
  INV_X1 U667 ( .A(G868), .ZN(n649) );
  NOR2_X1 U668 ( .A1(G286), .A2(n649), .ZN(n597) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U670 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U671 ( .A1(n604), .A2(G559), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n598), .A2(n990), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n599), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U674 ( .A1(G868), .A2(n975), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n990), .A2(G868), .ZN(n600) );
  NOR2_X1 U676 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U678 ( .A1(G559), .A2(n990), .ZN(n603) );
  XOR2_X1 U679 ( .A(n975), .B(n603), .Z(n646) );
  NAND2_X1 U680 ( .A1(n604), .A2(n646), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G93), .A2(n635), .ZN(n606) );
  NAND2_X1 U682 ( .A1(G80), .A2(n629), .ZN(n605) );
  NAND2_X1 U683 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n632), .A2(G55), .ZN(n607) );
  XOR2_X1 U685 ( .A(KEYINPUT74), .B(n607), .Z(n608) );
  NOR2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n631), .A2(G67), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n650) );
  XNOR2_X1 U689 ( .A(n612), .B(n650), .ZN(G145) );
  NAND2_X1 U690 ( .A1(G49), .A2(n632), .ZN(n614) );
  NAND2_X1 U691 ( .A1(G74), .A2(G651), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U693 ( .A1(n631), .A2(n615), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n616), .A2(G87), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(G288) );
  NAND2_X1 U696 ( .A1(G75), .A2(n629), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n619), .B(KEYINPUT78), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G62), .A2(n631), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G50), .A2(n632), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U701 ( .A(KEYINPUT76), .B(n622), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G88), .A2(n635), .ZN(n623) );
  XNOR2_X1 U703 ( .A(KEYINPUT77), .B(n623), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U706 ( .A(KEYINPUT79), .B(n628), .ZN(G166) );
  NAND2_X1 U707 ( .A1(G73), .A2(n629), .ZN(n630) );
  XNOR2_X1 U708 ( .A(n630), .B(KEYINPUT2), .ZN(n640) );
  NAND2_X1 U709 ( .A1(G61), .A2(n631), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G48), .A2(n632), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G86), .A2(n635), .ZN(n636) );
  XNOR2_X1 U713 ( .A(KEYINPUT75), .B(n636), .ZN(n637) );
  NOR2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(G305) );
  XNOR2_X1 U716 ( .A(KEYINPUT19), .B(G288), .ZN(n645) );
  INV_X1 U717 ( .A(G299), .ZN(n978) );
  XNOR2_X1 U718 ( .A(G166), .B(G305), .ZN(n641) );
  XNOR2_X1 U719 ( .A(n641), .B(n650), .ZN(n642) );
  XNOR2_X1 U720 ( .A(n978), .B(n642), .ZN(n643) );
  XNOR2_X1 U721 ( .A(n643), .B(G290), .ZN(n644) );
  XNOR2_X1 U722 ( .A(n645), .B(n644), .ZN(n898) );
  XNOR2_X1 U723 ( .A(n646), .B(n898), .ZN(n647) );
  XNOR2_X1 U724 ( .A(KEYINPUT80), .B(n647), .ZN(n648) );
  NOR2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n652) );
  NOR2_X1 U726 ( .A1(G868), .A2(n650), .ZN(n651) );
  NOR2_X1 U727 ( .A1(n652), .A2(n651), .ZN(G295) );
  NAND2_X1 U728 ( .A1(G2078), .A2(G2084), .ZN(n653) );
  XOR2_X1 U729 ( .A(KEYINPUT20), .B(n653), .Z(n654) );
  NAND2_X1 U730 ( .A1(G2090), .A2(n654), .ZN(n655) );
  XNOR2_X1 U731 ( .A(KEYINPUT21), .B(n655), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n656), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U733 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U734 ( .A(KEYINPUT22), .B(KEYINPUT81), .Z(n658) );
  NAND2_X1 U735 ( .A1(G132), .A2(G82), .ZN(n657) );
  XNOR2_X1 U736 ( .A(n658), .B(n657), .ZN(n659) );
  NOR2_X1 U737 ( .A1(n659), .A2(G218), .ZN(n660) );
  NAND2_X1 U738 ( .A1(G96), .A2(n660), .ZN(n827) );
  NAND2_X1 U739 ( .A1(n827), .A2(G2106), .ZN(n665) );
  NOR2_X1 U740 ( .A1(G236), .A2(G238), .ZN(n662) );
  NOR2_X1 U741 ( .A1(G235), .A2(G237), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U743 ( .A(KEYINPUT82), .B(n663), .ZN(n828) );
  NAND2_X1 U744 ( .A1(n828), .A2(G567), .ZN(n664) );
  NAND2_X1 U745 ( .A1(n665), .A2(n664), .ZN(n829) );
  NAND2_X1 U746 ( .A1(G661), .A2(G483), .ZN(n666) );
  NOR2_X1 U747 ( .A1(n829), .A2(n666), .ZN(n826) );
  NAND2_X1 U748 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U749 ( .A1(n881), .A2(G138), .ZN(n669) );
  NAND2_X1 U750 ( .A1(G102), .A2(n880), .ZN(n667) );
  XOR2_X1 U751 ( .A(KEYINPUT83), .B(n667), .Z(n668) );
  NAND2_X1 U752 ( .A1(n669), .A2(n668), .ZN(n673) );
  NAND2_X1 U753 ( .A1(G126), .A2(n875), .ZN(n671) );
  NAND2_X1 U754 ( .A1(G114), .A2(n876), .ZN(n670) );
  NAND2_X1 U755 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U756 ( .A1(n673), .A2(n672), .ZN(G164) );
  INV_X1 U757 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U758 ( .A(G1986), .B(G290), .ZN(n986) );
  NOR2_X1 U759 ( .A1(G164), .A2(G1384), .ZN(n680) );
  NOR2_X1 U760 ( .A1(n679), .A2(n680), .ZN(n675) );
  XNOR2_X1 U761 ( .A(n675), .B(KEYINPUT84), .ZN(n817) );
  NAND2_X1 U762 ( .A1(n986), .A2(n817), .ZN(n805) );
  NOR2_X1 U763 ( .A1(G1981), .A2(G305), .ZN(n676) );
  XOR2_X1 U764 ( .A(n676), .B(KEYINPUT93), .Z(n677) );
  XNOR2_X1 U765 ( .A(KEYINPUT24), .B(n677), .ZN(n682) );
  INV_X1 U766 ( .A(KEYINPUT92), .ZN(n678) );
  XNOR2_X1 U767 ( .A(n679), .B(n678), .ZN(n681) );
  NAND2_X2 U768 ( .A1(n681), .A2(n680), .ZN(n729) );
  NAND2_X1 U769 ( .A1(n729), .A2(G8), .ZN(n762) );
  INV_X1 U770 ( .A(n762), .ZN(n750) );
  AND2_X1 U771 ( .A1(n682), .A2(n750), .ZN(n768) );
  NOR2_X1 U772 ( .A1(G1976), .A2(G288), .ZN(n754) );
  NOR2_X1 U773 ( .A1(G1971), .A2(G303), .ZN(n683) );
  NOR2_X1 U774 ( .A1(n754), .A2(n683), .ZN(n984) );
  INV_X1 U775 ( .A(G1996), .ZN(n796) );
  NOR2_X1 U776 ( .A1(n729), .A2(n796), .ZN(n684) );
  XOR2_X1 U777 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n685) );
  NAND2_X1 U778 ( .A1(n684), .A2(n685), .ZN(n689) );
  OR2_X1 U779 ( .A1(n729), .A2(n796), .ZN(n687) );
  INV_X1 U780 ( .A(n685), .ZN(n686) );
  NAND2_X1 U781 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U782 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U783 ( .A1(n729), .A2(G1341), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U785 ( .A1(n990), .A2(n701), .ZN(n698) );
  INV_X1 U786 ( .A(KEYINPUT94), .ZN(n693) );
  XNOR2_X2 U787 ( .A(n729), .B(n693), .ZN(n717) );
  NAND2_X1 U788 ( .A1(G2067), .A2(n717), .ZN(n694) );
  XNOR2_X1 U789 ( .A(n694), .B(KEYINPUT96), .ZN(n696) );
  NAND2_X1 U790 ( .A1(G1348), .A2(n729), .ZN(n695) );
  NAND2_X1 U791 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U792 ( .A1(n698), .A2(n697), .ZN(n700) );
  INV_X1 U793 ( .A(KEYINPUT97), .ZN(n699) );
  OR2_X1 U794 ( .A1(n990), .A2(n701), .ZN(n702) );
  NAND2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n710) );
  NAND2_X1 U796 ( .A1(G2072), .A2(n717), .ZN(n704) );
  XNOR2_X1 U797 ( .A(KEYINPUT27), .B(n704), .ZN(n708) );
  INV_X1 U798 ( .A(n717), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n705), .A2(G1956), .ZN(n706) );
  XNOR2_X1 U800 ( .A(n706), .B(KEYINPUT95), .ZN(n707) );
  NOR2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n711), .A2(n978), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n714) );
  NOR2_X1 U804 ( .A1(n711), .A2(n978), .ZN(n712) );
  XOR2_X1 U805 ( .A(n712), .B(KEYINPUT28), .Z(n713) );
  NAND2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n716) );
  XOR2_X1 U807 ( .A(KEYINPUT29), .B(KEYINPUT98), .Z(n715) );
  XNOR2_X1 U808 ( .A(n716), .B(n715), .ZN(n721) );
  XNOR2_X1 U809 ( .A(KEYINPUT25), .B(G2078), .ZN(n952) );
  NAND2_X1 U810 ( .A1(n717), .A2(n952), .ZN(n719) );
  INV_X1 U811 ( .A(G1961), .ZN(n997) );
  NAND2_X1 U812 ( .A1(n997), .A2(n729), .ZN(n718) );
  NAND2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n725) );
  NAND2_X1 U814 ( .A1(n725), .A2(G171), .ZN(n720) );
  NAND2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n742) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n762), .ZN(n744) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n729), .ZN(n743) );
  NOR2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n722) );
  NAND2_X1 U819 ( .A1(G8), .A2(n722), .ZN(n723) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n723), .ZN(n724) );
  NOR2_X1 U821 ( .A1(G168), .A2(n724), .ZN(n727) );
  NOR2_X1 U822 ( .A1(G171), .A2(n725), .ZN(n726) );
  NOR2_X1 U823 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U824 ( .A(KEYINPUT31), .B(n728), .Z(n741) );
  INV_X1 U825 ( .A(G8), .ZN(n734) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n729), .ZN(n731) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n762), .ZN(n730) );
  NOR2_X1 U828 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U829 ( .A1(n732), .A2(G303), .ZN(n733) );
  OR2_X1 U830 ( .A1(n734), .A2(n733), .ZN(n736) );
  AND2_X1 U831 ( .A1(n741), .A2(n736), .ZN(n735) );
  NAND2_X1 U832 ( .A1(n742), .A2(n735), .ZN(n739) );
  INV_X1 U833 ( .A(n736), .ZN(n737) );
  OR2_X1 U834 ( .A1(n737), .A2(G286), .ZN(n738) );
  NAND2_X1 U835 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U836 ( .A(n740), .B(KEYINPUT32), .ZN(n749) );
  AND2_X1 U837 ( .A1(n742), .A2(n741), .ZN(n747) );
  AND2_X1 U838 ( .A1(G8), .A2(n743), .ZN(n745) );
  OR2_X1 U839 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U840 ( .A1(n749), .A2(n748), .ZN(n760) );
  AND2_X1 U841 ( .A1(n984), .A2(n760), .ZN(n752) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n979) );
  NAND2_X1 U843 ( .A1(n979), .A2(n750), .ZN(n751) );
  NOR2_X1 U844 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U845 ( .A1(KEYINPUT33), .A2(n753), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n754), .A2(KEYINPUT33), .ZN(n755) );
  XOR2_X1 U847 ( .A(G1981), .B(G305), .Z(n972) );
  OR2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n765) );
  NOR2_X1 U849 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U850 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U853 ( .A(KEYINPUT99), .B(n763), .Z(n764) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U855 ( .A(n766), .B(KEYINPUT100), .ZN(n767) );
  NOR2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n803) );
  XOR2_X1 U857 ( .A(G2067), .B(KEYINPUT37), .Z(n769) );
  XNOR2_X1 U858 ( .A(KEYINPUT85), .B(n769), .ZN(n814) );
  XNOR2_X1 U859 ( .A(KEYINPUT86), .B(KEYINPUT34), .ZN(n773) );
  NAND2_X1 U860 ( .A1(G104), .A2(n880), .ZN(n771) );
  NAND2_X1 U861 ( .A1(G140), .A2(n881), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U863 ( .A(n773), .B(n772), .ZN(n780) );
  XNOR2_X1 U864 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n875), .A2(G128), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n876), .A2(G116), .ZN(n774) );
  XOR2_X1 U867 ( .A(KEYINPUT87), .B(n774), .Z(n775) );
  NAND2_X1 U868 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U869 ( .A(n778), .B(n777), .Z(n779) );
  NOR2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U871 ( .A(KEYINPUT36), .B(n781), .ZN(n893) );
  NOR2_X1 U872 ( .A1(n814), .A2(n893), .ZN(n929) );
  NAND2_X1 U873 ( .A1(n929), .A2(n817), .ZN(n812) );
  NAND2_X1 U874 ( .A1(G95), .A2(n880), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G131), .A2(n881), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G119), .A2(n875), .ZN(n785) );
  NAND2_X1 U878 ( .A1(G107), .A2(n876), .ZN(n784) );
  NAND2_X1 U879 ( .A1(n785), .A2(n784), .ZN(n786) );
  OR2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n858) );
  XOR2_X1 U881 ( .A(KEYINPUT89), .B(G1991), .Z(n958) );
  AND2_X1 U882 ( .A1(n858), .A2(n958), .ZN(n799) );
  NAND2_X1 U883 ( .A1(G117), .A2(n876), .ZN(n794) );
  NAND2_X1 U884 ( .A1(G129), .A2(n875), .ZN(n789) );
  NAND2_X1 U885 ( .A1(G141), .A2(n881), .ZN(n788) );
  NAND2_X1 U886 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U887 ( .A1(n880), .A2(G105), .ZN(n790) );
  XOR2_X1 U888 ( .A(KEYINPUT38), .B(n790), .Z(n791) );
  NOR2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U891 ( .A(n795), .B(KEYINPUT90), .ZN(n872) );
  INV_X1 U892 ( .A(n872), .ZN(n797) );
  NOR2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n931) );
  XNOR2_X1 U895 ( .A(KEYINPUT91), .B(n817), .ZN(n800) );
  NOR2_X1 U896 ( .A1(n931), .A2(n800), .ZN(n809) );
  INV_X1 U897 ( .A(n809), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n812), .A2(n801), .ZN(n802) );
  NOR2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n820) );
  NOR2_X1 U901 ( .A1(G1996), .A2(n872), .ZN(n934) );
  NOR2_X1 U902 ( .A1(n958), .A2(n858), .ZN(n926) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n806) );
  XOR2_X1 U904 ( .A(n806), .B(KEYINPUT101), .Z(n807) );
  NOR2_X1 U905 ( .A1(n926), .A2(n807), .ZN(n808) );
  NOR2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U907 ( .A1(n934), .A2(n810), .ZN(n811) );
  XNOR2_X1 U908 ( .A(KEYINPUT39), .B(n811), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n893), .A2(n814), .ZN(n815) );
  XNOR2_X1 U911 ( .A(n815), .B(KEYINPUT102), .ZN(n941) );
  NAND2_X1 U912 ( .A1(n816), .A2(n941), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n822) );
  XOR2_X1 U915 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n821) );
  XNOR2_X1 U916 ( .A(n822), .B(n821), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U919 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U923 ( .A(G132), .ZN(G219) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G82), .ZN(G220) );
  NOR2_X1 U926 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  INV_X1 U928 ( .A(n829), .ZN(G319) );
  XOR2_X1 U929 ( .A(G2100), .B(G2096), .Z(n831) );
  XNOR2_X1 U930 ( .A(KEYINPUT42), .B(G2678), .ZN(n830) );
  XNOR2_X1 U931 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U932 ( .A(KEYINPUT43), .B(G2090), .Z(n833) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n832) );
  XNOR2_X1 U934 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U935 ( .A(n835), .B(n834), .Z(n837) );
  XNOR2_X1 U936 ( .A(G2078), .B(G2084), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(G227) );
  XOR2_X1 U938 ( .A(KEYINPUT106), .B(KEYINPUT109), .Z(n839) );
  XNOR2_X1 U939 ( .A(G2474), .B(KEYINPUT108), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U941 ( .A(n840), .B(KEYINPUT107), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n850) );
  XOR2_X1 U944 ( .A(G1956), .B(G1971), .Z(n844) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1976), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U947 ( .A(KEYINPUT41), .B(G1961), .Z(n846) );
  XNOR2_X1 U948 ( .A(G1981), .B(G1966), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U950 ( .A(n848), .B(n847), .Z(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(G229) );
  NAND2_X1 U952 ( .A1(G100), .A2(n880), .ZN(n852) );
  NAND2_X1 U953 ( .A1(G112), .A2(n876), .ZN(n851) );
  NAND2_X1 U954 ( .A1(n852), .A2(n851), .ZN(n857) );
  NAND2_X1 U955 ( .A1(n875), .A2(G124), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U957 ( .A1(G136), .A2(n881), .ZN(n854) );
  NAND2_X1 U958 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U959 ( .A1(n857), .A2(n856), .ZN(G162) );
  XOR2_X1 U960 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n860) );
  XOR2_X1 U961 ( .A(n858), .B(G162), .Z(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n923), .B(n861), .ZN(n874) );
  NAND2_X1 U964 ( .A1(G127), .A2(n875), .ZN(n863) );
  NAND2_X1 U965 ( .A1(G115), .A2(n876), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U967 ( .A(KEYINPUT47), .B(n864), .ZN(n870) );
  NAND2_X1 U968 ( .A1(G103), .A2(n880), .ZN(n865) );
  XOR2_X1 U969 ( .A(KEYINPUT112), .B(n865), .Z(n868) );
  NAND2_X1 U970 ( .A1(G139), .A2(n881), .ZN(n866) );
  XNOR2_X1 U971 ( .A(KEYINPUT113), .B(n866), .ZN(n867) );
  NOR2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U974 ( .A(KEYINPUT114), .B(n871), .ZN(n919) );
  XNOR2_X1 U975 ( .A(n872), .B(n919), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n889) );
  NAND2_X1 U977 ( .A1(G130), .A2(n875), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G118), .A2(n876), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U980 ( .A(KEYINPUT110), .B(n879), .ZN(n887) );
  NAND2_X1 U981 ( .A1(G106), .A2(n880), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G142), .A2(n881), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(KEYINPUT111), .B(n884), .ZN(n885) );
  XNOR2_X1 U985 ( .A(KEYINPUT45), .B(n885), .ZN(n886) );
  NOR2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U987 ( .A(n889), .B(n888), .Z(n891) );
  XNOR2_X1 U988 ( .A(G164), .B(G160), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U990 ( .A(n893), .B(n892), .Z(n894) );
  NOR2_X1 U991 ( .A1(G37), .A2(n894), .ZN(n895) );
  XOR2_X1 U992 ( .A(KEYINPUT115), .B(n895), .Z(G395) );
  XNOR2_X1 U993 ( .A(n975), .B(KEYINPUT116), .ZN(n897) );
  XNOR2_X1 U994 ( .A(G171), .B(n990), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n900) );
  XNOR2_X1 U996 ( .A(G286), .B(n898), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U998 ( .A1(G37), .A2(n901), .ZN(G397) );
  XNOR2_X1 U999 ( .A(G2446), .B(KEYINPUT104), .ZN(n911) );
  XOR2_X1 U1000 ( .A(KEYINPUT105), .B(G2427), .Z(n903) );
  XNOR2_X1 U1001 ( .A(G2435), .B(G2438), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1003 ( .A(G2454), .B(G2430), .Z(n905) );
  XNOR2_X1 U1004 ( .A(G1348), .B(G1341), .ZN(n904) );
  XNOR2_X1 U1005 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1006 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1007 ( .A(G2443), .B(G2451), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  NAND2_X1 U1010 ( .A1(n912), .A2(G14), .ZN(n918) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(n918), .ZN(G401) );
  XNOR2_X1 U1019 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1028) );
  INV_X1 U1020 ( .A(KEYINPUT55), .ZN(n947) );
  XOR2_X1 U1021 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n944) );
  XOR2_X1 U1022 ( .A(G164), .B(G2078), .Z(n921) );
  XNOR2_X1 U1023 ( .A(G2072), .B(n919), .ZN(n920) );
  NOR2_X1 U1024 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1025 ( .A(KEYINPUT50), .B(n922), .Z(n940) );
  XNOR2_X1 U1026 ( .A(G160), .B(G2084), .ZN(n924) );
  NAND2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1029 ( .A(KEYINPUT117), .B(n927), .ZN(n928) );
  NOR2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n937) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n932) );
  XNOR2_X1 U1033 ( .A(KEYINPUT118), .B(n932), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(KEYINPUT51), .B(n935), .ZN(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(KEYINPUT119), .B(n938), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1040 ( .A(n944), .B(n943), .ZN(n945) );
  XOR2_X1 U1041 ( .A(KEYINPUT52), .B(n945), .Z(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n948), .A2(G29), .ZN(n1026) );
  XOR2_X1 U1044 ( .A(G29), .B(KEYINPUT124), .Z(n970) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G32), .B(G1996), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n957) );
  XOR2_X1 U1048 ( .A(G2072), .B(G33), .Z(n951) );
  NAND2_X1 U1049 ( .A1(n951), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G27), .B(n952), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(KEYINPUT123), .B(n953), .ZN(n954) );
  NOR2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G25), .B(n958), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1056 ( .A(KEYINPUT53), .B(n961), .Z(n964) );
  XOR2_X1 U1057 ( .A(KEYINPUT54), .B(G34), .Z(n962) );
  XNOR2_X1 U1058 ( .A(G2084), .B(n962), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(KEYINPUT122), .B(G2090), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(G35), .B(n965), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n968), .B(KEYINPUT55), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n971), .ZN(n1024) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n996) );
  XNOR2_X1 U1067 ( .A(G1966), .B(G168), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n974), .B(KEYINPUT57), .ZN(n994) );
  XOR2_X1 U1070 ( .A(G171), .B(G1961), .Z(n977) );
  XNOR2_X1 U1071 ( .A(n975), .B(G1341), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n989) );
  XNOR2_X1 U1073 ( .A(G1956), .B(n978), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n982) );
  AND2_X1 U1075 ( .A1(G303), .A2(G1971), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1079 ( .A(KEYINPUT125), .B(n987), .Z(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n992) );
  XOR2_X1 U1081 ( .A(G1348), .B(n990), .Z(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n1022) );
  INV_X1 U1085 ( .A(G16), .ZN(n1020) );
  XNOR2_X1 U1086 ( .A(G5), .B(n997), .ZN(n1017) );
  XOR2_X1 U1087 ( .A(G1966), .B(G21), .Z(n1007) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(n998), .B(G4), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G1981), .B(G6), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G1341), .B(G19), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G20), .B(G1956), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(n1005), .B(KEYINPUT60), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT126), .B(n1008), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(G1976), .B(G23), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XOR2_X1 U1102 ( .A(G1986), .B(G24), .Z(n1011) );
  NAND2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1104 ( .A(KEYINPUT58), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1018), .Z(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(n1028), .B(n1027), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

