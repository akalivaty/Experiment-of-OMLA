//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT76), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n190), .A2(G221), .ZN(new_n191));
  INV_X1    g005(.A(G469), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT78), .A2(G107), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT78), .A2(G107), .ZN(new_n194));
  AOI21_X1  g008(.A(G104), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G107), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT79), .A3(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(G101), .B1(new_n195), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT80), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n206), .A2(G128), .B1(new_n207), .B2(G146), .ZN(new_n208));
  OAI22_X1  g022(.A1(new_n205), .A2(new_n208), .B1(G128), .B2(new_n204), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT80), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n210), .B(G101), .C1(new_n195), .C2(new_n201), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n199), .A2(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n199), .A2(G104), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n212), .B1(KEYINPUT3), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n193), .A2(new_n194), .ZN(new_n216));
  OR2_X1    g030(.A1(new_n197), .A2(KEYINPUT3), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n203), .A2(new_n209), .A3(new_n211), .A4(new_n218), .ZN(new_n219));
  XOR2_X1   g033(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G101), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n218), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n225), .A3(G101), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n207), .A2(G146), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  OAI22_X1  g047(.A1(new_n228), .A2(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n204), .A2(new_n231), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n221), .B1(new_n227), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G137), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(G137), .ZN(new_n243));
  INV_X1    g057(.A(G137), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT11), .A3(G134), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT64), .A2(G131), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n242), .A2(new_n245), .A3(new_n247), .A4(new_n243), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n203), .A2(new_n211), .A3(new_n218), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT82), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n203), .A2(KEYINPUT82), .A3(new_n211), .A4(new_n218), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n255), .A2(KEYINPUT10), .A3(new_n209), .A4(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n239), .A2(new_n252), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G110), .B(G140), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n260), .A2(G227), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n259), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n219), .A2(KEYINPUT83), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n229), .A2(G143), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n207), .A2(G146), .ZN(new_n267));
  AOI21_X1  g081(.A(G128), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n206), .B1(new_n228), .B2(new_n230), .ZN(new_n269));
  INV_X1    g083(.A(new_n208), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n253), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n253), .A2(KEYINPUT83), .A3(new_n271), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT12), .B1(new_n275), .B2(new_n251), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT12), .ZN(new_n277));
  AOI211_X1 g091(.A(new_n277), .B(new_n252), .C1(new_n273), .C2(new_n274), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(KEYINPUT84), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n275), .A2(KEYINPUT12), .A3(new_n251), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT84), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n264), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n257), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n251), .B1(new_n284), .B2(new_n238), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n263), .B1(new_n285), .B2(new_n258), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n192), .B(new_n189), .C1(new_n283), .C2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT85), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n284), .A2(new_n238), .A3(new_n251), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(new_n262), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n275), .A2(KEYINPUT84), .A3(KEYINPUT12), .A4(new_n251), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n252), .B1(new_n273), .B2(new_n274), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n292), .B1(KEYINPUT12), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n278), .A2(KEYINPUT84), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n286), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT85), .A3(new_n192), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n289), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n285), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n264), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n275), .A2(new_n251), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n277), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n282), .A2(new_n304), .A3(new_n292), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n258), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n262), .B(KEYINPUT77), .Z(new_n307));
  AOI21_X1  g121(.A(new_n302), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G469), .B1(new_n308), .B2(G902), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n191), .B1(new_n300), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT16), .ZN(new_n312));
  INV_X1    g126(.A(G140), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(G125), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(G125), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n314), .B1(new_n318), .B2(new_n312), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n229), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n316), .A2(KEYINPUT16), .A3(G140), .ZN(new_n321));
  XNOR2_X1  g135(.A(G125), .B(G140), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(KEYINPUT16), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G146), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G110), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT24), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT24), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G110), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT70), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT70), .B1(new_n327), .B2(new_n329), .ZN(new_n331));
  INV_X1    g145(.A(G128), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G119), .ZN(new_n333));
  INV_X1    g147(.A(G119), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G128), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OR3_X1    g150(.A1(new_n330), .A2(new_n331), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n334), .B2(G128), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n332), .A2(KEYINPUT23), .A3(G119), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n335), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n325), .B(new_n337), .C1(new_n326), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT72), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n322), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n346), .A3(new_n229), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n324), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n342), .A2(KEYINPUT71), .A3(new_n326), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n336), .B1(new_n330), .B2(new_n331), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT71), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n341), .B2(G110), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n348), .A2(new_n353), .A3(KEYINPUT73), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT73), .B1(new_n348), .B2(new_n353), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n343), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT22), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(G137), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n343), .B(new_n359), .C1(new_n354), .C2(new_n355), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n189), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT74), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(KEYINPUT25), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n365), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n361), .A2(new_n189), .A3(new_n367), .A4(new_n362), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT69), .B(G217), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(G234), .B2(new_n189), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n311), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n371), .ZN(new_n373));
  AOI211_X1 g187(.A(KEYINPUT75), .B(new_n373), .C1(new_n366), .C2(new_n368), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n361), .A2(new_n362), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n371), .A2(G902), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n380));
  NOR2_X1   g194(.A1(G116), .A2(G119), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(G116), .A2(G119), .ZN(new_n383));
  NAND2_X1  g197(.A1(KEYINPUT2), .A2(G113), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(KEYINPUT2), .A2(G113), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n382), .B(new_n383), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n386), .ZN(new_n388));
  INV_X1    g202(.A(new_n383), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n388), .B(new_n384), .C1(new_n389), .C2(new_n381), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G131), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n242), .A2(new_n245), .A3(new_n393), .A4(new_n243), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n241), .A2(G137), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n244), .A2(G134), .ZN(new_n396));
  OAI21_X1  g210(.A(G131), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n271), .A2(new_n398), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n249), .A2(new_n250), .B1(new_n234), .B2(new_n235), .ZN(new_n400));
  OAI211_X1 g214(.A(KEYINPUT65), .B(KEYINPUT30), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n251), .A2(new_n236), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n266), .A2(new_n267), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n208), .B1(new_n206), .B2(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n397), .B(new_n394), .C1(new_n404), .C2(new_n268), .ZN(new_n405));
  OR2_X1    g219(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n406));
  NAND2_X1  g220(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n402), .A2(new_n405), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n392), .B1(new_n401), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT26), .B(G101), .ZN(new_n410));
  NOR2_X1   g224(.A1(G237), .A2(G953), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G210), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n410), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT66), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n391), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n387), .A2(new_n390), .A3(KEYINPUT66), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n420), .A2(new_n399), .A3(new_n400), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n409), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(KEYINPUT28), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n402), .A2(new_n405), .A3(new_n418), .A4(new_n419), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT28), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n402), .A2(new_n405), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n424), .A2(new_n425), .B1(new_n426), .B2(new_n391), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n415), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n380), .B1(new_n422), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n424), .A2(new_n425), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n415), .A2(new_n380), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n426), .A2(new_n420), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT68), .A3(new_n424), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT68), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n426), .A2(new_n434), .A3(new_n420), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n430), .B(new_n431), .C1(new_n436), .C2(new_n425), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n429), .A2(new_n189), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G472), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n401), .A2(new_n408), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n391), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n416), .A3(new_n424), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT31), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n416), .B1(new_n423), .B2(new_n427), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n421), .B1(new_n440), .B2(new_n391), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT31), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(new_n416), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(G472), .A2(G902), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(KEYINPUT32), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n439), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT32), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n449), .A2(new_n450), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n379), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n370), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n188), .A2(new_n260), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G128), .B(G143), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT13), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n207), .A2(G128), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n460), .B(G134), .C1(KEYINPUT13), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n241), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G116), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT94), .ZN(new_n466));
  INV_X1    g280(.A(G122), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT94), .A2(G122), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(G122), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n216), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n193), .A2(new_n194), .ZN(new_n474));
  INV_X1    g288(.A(new_n469), .ZN(new_n475));
  NOR2_X1   g289(.A1(KEYINPUT94), .A2(G122), .ZN(new_n476));
  OAI21_X1  g290(.A(G116), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(new_n477), .A3(new_n471), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT95), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT95), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n473), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n464), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n471), .B(KEYINPUT14), .ZN(new_n484));
  OAI21_X1  g298(.A(G107), .B1(new_n484), .B2(new_n470), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT96), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n474), .A2(new_n477), .A3(KEYINPUT96), .A4(new_n471), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n459), .B(new_n241), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n485), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n458), .B1(new_n483), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT97), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n462), .A2(new_n463), .ZN(new_n494));
  INV_X1    g308(.A(new_n482), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n481), .B1(new_n473), .B2(new_n478), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n458), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n490), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n492), .A2(new_n493), .A3(new_n499), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n497), .A2(KEYINPUT97), .A3(new_n490), .A4(new_n498), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n189), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT98), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT98), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n500), .A2(new_n504), .A3(new_n189), .A4(new_n501), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G478), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n502), .A2(new_n508), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT20), .ZN(new_n512));
  INV_X1    g326(.A(G237), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n260), .A3(G214), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(new_n207), .ZN(new_n515));
  AOI21_X1  g329(.A(G143), .B1(new_n411), .B2(G214), .ZN(new_n516));
  OAI21_X1  g330(.A(G131), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n514), .A2(new_n207), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n411), .A2(G143), .A3(G214), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n393), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT92), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n320), .A2(new_n324), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n517), .A2(new_n525), .A3(new_n518), .A4(new_n521), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n517), .A2(new_n518), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n523), .A2(new_n524), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(G113), .B(G122), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(new_n197), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n318), .A2(G146), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n347), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(KEYINPUT18), .A2(G131), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n519), .A2(new_n520), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(KEYINPUT18), .B(G131), .C1(new_n515), .C2(new_n516), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n528), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n517), .A2(new_n521), .B1(G146), .B2(new_n323), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT19), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n344), .A2(new_n346), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n318), .A2(KEYINPUT19), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n229), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n536), .ZN(new_n544));
  INV_X1    g358(.A(new_n530), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n537), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(G475), .A2(G902), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n512), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n548), .ZN(new_n550));
  AOI211_X1 g364(.A(KEYINPUT20), .B(new_n550), .C1(new_n537), .C2(new_n546), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n528), .A2(new_n536), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n545), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n553), .B2(new_n537), .ZN(new_n554));
  INV_X1    g368(.A(G475), .ZN(new_n555));
  OAI22_X1  g369(.A1(new_n549), .A2(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT93), .ZN(new_n557));
  INV_X1    g371(.A(new_n537), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n530), .B1(new_n528), .B2(new_n536), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n189), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G475), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n561), .B(new_n562), .C1(new_n549), .C2(new_n551), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n260), .A2(G952), .ZN(new_n565));
  NAND2_X1  g379(.A1(G234), .A2(G237), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT21), .B(G898), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(G902), .A3(G953), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n511), .A2(new_n564), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n390), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT86), .B(KEYINPUT5), .Z(new_n575));
  NOR2_X1   g389(.A1(new_n389), .A2(new_n381), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(G113), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n465), .A2(G119), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n578), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n574), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n255), .A2(new_n256), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(G110), .B(G122), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n224), .A2(new_n391), .A3(new_n226), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT6), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n583), .B1(new_n582), .B2(new_n584), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT87), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n582), .A2(new_n584), .ZN(new_n589));
  INV_X1    g403(.A(new_n583), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT87), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n591), .A2(new_n592), .A3(KEYINPUT6), .A4(new_n585), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n237), .A2(G125), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(G125), .B2(new_n209), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n260), .A2(G224), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g411(.A(KEYINPUT6), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n587), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n588), .A2(new_n593), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n594), .A2(KEYINPUT90), .B1(KEYINPUT7), .B2(new_n596), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(new_n595), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT88), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT5), .ZN(new_n604));
  OAI22_X1  g418(.A1(new_n580), .A2(new_n603), .B1(new_n604), .B2(new_n576), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n580), .A2(new_n603), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n390), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT89), .ZN(new_n608));
  OR3_X1    g422(.A1(new_n607), .A2(new_n608), .A3(new_n253), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n608), .B1(new_n607), .B2(new_n253), .ZN(new_n610));
  INV_X1    g424(.A(new_n253), .ZN(new_n611));
  OR2_X1    g425(.A1(new_n611), .A2(new_n581), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n583), .B(KEYINPUT8), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n602), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n615), .B2(new_n585), .ZN(new_n616));
  OAI21_X1  g430(.A(G210), .B1(G237), .B2(G902), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n617), .B(KEYINPUT91), .Z(new_n618));
  NAND3_X1  g432(.A1(new_n600), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(G214), .B1(G237), .B2(G902), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n618), .B1(new_n600), .B2(new_n616), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n620), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n310), .A2(new_n456), .A3(new_n573), .A4(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT99), .B(G101), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G3));
  AOI21_X1  g441(.A(new_n447), .B1(new_n446), .B2(new_n416), .ZN(new_n628));
  NOR4_X1   g442(.A1(new_n409), .A2(KEYINPUT31), .A3(new_n415), .A4(new_n421), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n628), .A2(new_n629), .A3(new_n444), .ZN(new_n630));
  OAI21_X1  g444(.A(G472), .B1(new_n630), .B2(G902), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n454), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n379), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n310), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n506), .A2(new_n507), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n500), .A2(new_n636), .A3(new_n501), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n492), .A2(KEYINPUT33), .A3(new_n499), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(G478), .A3(new_n189), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n641), .A2(new_n564), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n624), .A2(new_n571), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  NAND2_X1  g460(.A1(new_n624), .A2(new_n571), .ZN(new_n647));
  INV_X1    g461(.A(new_n511), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n551), .A2(KEYINPUT100), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n649), .A2(new_n549), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n551), .A2(KEYINPUT100), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n561), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n647), .A2(new_n648), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n634), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NOR2_X1   g470(.A1(new_n360), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n356), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n377), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n632), .B1(new_n375), .B2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n310), .A2(new_n573), .A3(new_n624), .A4(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  AOI21_X1  g477(.A(KEYINPUT85), .B1(new_n298), .B2(new_n192), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n286), .B1(new_n305), .B2(new_n291), .ZN(new_n665));
  NOR4_X1   g479(.A1(new_n665), .A2(new_n288), .A3(G469), .A4(G902), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n309), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n191), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n439), .A2(new_n451), .ZN(new_n669));
  INV_X1    g483(.A(new_n450), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n453), .B1(new_n630), .B2(new_n670), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n375), .A2(new_n659), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n667), .A2(new_n668), .A3(new_n624), .A4(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n567), .B1(G900), .B2(new_n570), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n561), .B(new_n674), .C1(new_n650), .C2(new_n651), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n675), .A2(new_n648), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n332), .ZN(G30));
  NOR2_X1   g492(.A1(new_n620), .A2(new_n623), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT38), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n375), .A2(new_n659), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n509), .A2(new_n510), .B1(new_n557), .B2(new_n563), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n621), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT103), .B1(new_n681), .B2(new_n683), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n680), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(G472), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n436), .B2(new_n415), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n416), .B1(new_n409), .B2(new_n421), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n454), .B2(new_n453), .ZN(new_n693));
  AOI21_X1  g507(.A(KEYINPUT101), .B1(new_n693), .B2(new_n451), .ZN(new_n694));
  INV_X1    g508(.A(new_n692), .ZN(new_n695));
  AND4_X1   g509(.A1(KEYINPUT101), .A2(new_n671), .A3(new_n451), .A4(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n688), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n674), .B(KEYINPUT39), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT40), .B1(new_n310), .B2(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n310), .A2(KEYINPUT40), .A3(new_n701), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT104), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n700), .B(new_n706), .C1(new_n702), .C2(new_n703), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n207), .ZN(G45));
  NAND2_X1  g523(.A1(new_n642), .A2(new_n674), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n310), .A2(new_n624), .A3(new_n672), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  NAND2_X1  g527(.A1(new_n298), .A2(KEYINPUT105), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n665), .B2(G902), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(G469), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n300), .A2(new_n668), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n300), .A2(KEYINPUT106), .A3(new_n668), .A4(new_n717), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n456), .A3(new_n643), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND4_X1  g538(.A1(new_n720), .A2(new_n653), .A3(new_n456), .A4(new_n721), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND4_X1  g540(.A1(new_n300), .A2(new_n668), .A3(new_n624), .A4(new_n717), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n672), .A2(new_n573), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  NAND2_X1  g546(.A1(new_n600), .A2(new_n616), .ZN(new_n733));
  INV_X1    g547(.A(new_n618), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n682), .A2(new_n621), .A3(new_n735), .A4(new_n619), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n430), .B1(new_n436), .B2(new_n425), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n415), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n443), .A3(new_n448), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n450), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n631), .ZN(new_n741));
  NOR4_X1   g555(.A1(new_n736), .A2(new_n379), .A3(new_n572), .A4(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n720), .A2(new_n721), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  AND3_X1   g558(.A1(new_n300), .A2(new_n668), .A3(new_n717), .ZN(new_n745));
  INV_X1    g559(.A(new_n741), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n681), .A2(new_n642), .A3(new_n674), .A4(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n745), .A2(new_n748), .A3(KEYINPUT108), .A4(new_n624), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n727), .B2(new_n747), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  XNOR2_X1  g567(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n667), .A2(KEYINPUT109), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n309), .B(new_n756), .C1(new_n664), .C2(new_n666), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n668), .A2(new_n621), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n679), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n755), .A2(new_n456), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n754), .B1(new_n760), .B2(new_n710), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n755), .A2(new_n757), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n642), .A2(KEYINPUT42), .A3(new_n674), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n454), .A2(KEYINPUT111), .A3(new_n453), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT111), .B1(new_n454), .B2(new_n453), .ZN(new_n765));
  OR3_X1    g579(.A1(new_n764), .A2(new_n452), .A3(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n375), .A2(new_n378), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n764), .A2(new_n452), .A3(new_n765), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT112), .B1(new_n770), .B2(new_n379), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n763), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n762), .A2(new_n772), .A3(new_n759), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n761), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G131), .ZN(G33));
  NOR2_X1   g589(.A1(new_n760), .A2(new_n676), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n241), .ZN(G36));
  NAND3_X1  g591(.A1(new_n641), .A2(new_n563), .A3(new_n557), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT43), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n632), .A3(new_n681), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n679), .A2(new_n622), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(G469), .B1(new_n308), .B2(KEYINPUT45), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n308), .A2(KEYINPUT45), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n787), .B2(new_n788), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(G469), .A2(G902), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(KEYINPUT114), .A3(KEYINPUT46), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n793), .B1(new_n789), .B2(new_n791), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT46), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n795), .A2(new_n796), .B1(new_n289), .B2(new_n299), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n795), .B2(new_n796), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n794), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n786), .A2(new_n668), .A3(new_n701), .A4(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n668), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT47), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT47), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n800), .A2(new_n805), .A3(new_n668), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n711), .A2(new_n455), .A3(new_n379), .A4(new_n785), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n804), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  NOR2_X1   g624(.A1(new_n729), .A2(new_n730), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n727), .A2(KEYINPUT107), .A3(new_n728), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n722), .B(new_n725), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n648), .A2(new_n564), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n642), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n647), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n310), .A3(new_n633), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n743), .A2(new_n817), .A3(new_n625), .A4(new_n661), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n776), .B1(new_n761), .B2(new_n773), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n675), .A2(new_n511), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n785), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n785), .A2(KEYINPUT115), .A3(new_n821), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n310), .A3(new_n672), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n748), .A2(new_n755), .A3(new_n757), .A4(new_n759), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n819), .A2(KEYINPUT53), .A3(new_n820), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n830));
  INV_X1    g644(.A(new_n736), .ZN(new_n831));
  INV_X1    g645(.A(new_n372), .ZN(new_n832));
  INV_X1    g646(.A(new_n374), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n668), .A2(new_n674), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n832), .A2(new_n833), .A3(new_n659), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n696), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n693), .A2(new_n451), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT101), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n835), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n755), .A2(new_n831), .A3(new_n840), .A4(new_n757), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT116), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n697), .A2(new_n736), .A3(new_n835), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n755), .A4(new_n757), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n842), .A2(new_n712), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n677), .B1(new_n749), .B2(new_n751), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n845), .A2(new_n712), .ZN(new_n849));
  AND4_X1   g663(.A1(KEYINPUT52), .A2(new_n847), .A3(new_n849), .A4(new_n842), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n830), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  INV_X1    g666(.A(new_n677), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n752), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n842), .A2(new_n712), .A3(new_n845), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n847), .A2(new_n849), .A3(KEYINPUT52), .A4(new_n842), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(KEYINPUT117), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n829), .B1(new_n851), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n818), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n725), .A2(new_n722), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n731), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n820), .A2(new_n828), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n856), .A2(new_n857), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT53), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n859), .A2(KEYINPUT54), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n848), .A2(new_n850), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n819), .A2(new_n820), .A3(new_n828), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n856), .A2(KEYINPUT117), .A3(new_n857), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT117), .B1(new_n856), .B2(new_n857), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n864), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n872), .B1(new_n875), .B2(new_n871), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n868), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n300), .A2(new_n717), .ZN(new_n879));
  NOR4_X1   g693(.A1(new_n879), .A2(new_n567), .A3(new_n679), .A4(new_n758), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n780), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n769), .A2(new_n771), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n883), .A2(KEYINPUT119), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(KEYINPUT119), .ZN(new_n885));
  OR2_X1    g699(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n886));
  NAND2_X1  g700(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n887));
  AND4_X1   g701(.A1(new_n884), .A2(new_n885), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n886), .B1(new_n884), .B2(new_n885), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n699), .A2(new_n767), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n890), .A2(new_n880), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n642), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n767), .A2(new_n566), .A3(new_n565), .A4(new_n746), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n779), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n892), .B(new_n565), .C1(new_n727), .C2(new_n895), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n888), .A2(new_n889), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n894), .A2(new_n785), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n804), .A2(new_n806), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n300), .A2(new_n191), .A3(new_n717), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n641), .A2(new_n564), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n891), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n880), .A2(new_n681), .A3(new_n746), .A4(new_n780), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n680), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n894), .A2(new_n622), .A3(new_n907), .A4(new_n745), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT50), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n902), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n909), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(KEYINPUT118), .A3(new_n905), .A4(new_n904), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n912), .A3(KEYINPUT51), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n901), .A2(new_n909), .A3(new_n906), .ZN(new_n914));
  OAI221_X1 g728(.A(new_n897), .B1(new_n901), .B2(new_n913), .C1(new_n914), .C2(KEYINPUT51), .ZN(new_n915));
  OAI22_X1  g729(.A1(new_n878), .A2(new_n915), .B1(G952), .B2(G953), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n879), .B(KEYINPUT49), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n680), .A2(new_n758), .A3(new_n778), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n890), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(G75));
  NOR2_X1   g734(.A1(new_n859), .A2(new_n866), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n189), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT56), .B1(new_n922), .B2(new_n618), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n588), .A2(new_n593), .A3(new_n599), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n597), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT55), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n260), .A2(G952), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n923), .B2(new_n927), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n928), .A2(new_n931), .ZN(G51));
  NOR3_X1   g746(.A1(new_n921), .A2(new_n189), .A3(new_n792), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n793), .B(KEYINPUT57), .Z(new_n934));
  NOR3_X1   g748(.A1(new_n862), .A2(new_n863), .A3(new_n871), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n873), .B2(new_n874), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n871), .B1(new_n869), .B2(new_n870), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n877), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n934), .B1(new_n867), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n665), .B(KEYINPUT121), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n933), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n939), .A2(KEYINPUT122), .A3(new_n940), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n929), .B1(new_n943), .B2(new_n944), .ZN(G54));
  NAND3_X1  g759(.A1(new_n922), .A2(KEYINPUT58), .A3(G475), .ZN(new_n946));
  INV_X1    g760(.A(new_n547), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(new_n929), .ZN(G60));
  NAND2_X1  g764(.A1(G478), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT59), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n639), .B1(new_n878), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n639), .B(new_n952), .C1(new_n867), .C2(new_n938), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n930), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n953), .A2(new_n955), .ZN(G63));
  NAND2_X1  g770(.A1(G217), .A2(G902), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT60), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n921), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n658), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n376), .B(KEYINPUT123), .Z(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n921), .B2(new_n958), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n930), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n960), .A2(KEYINPUT61), .A3(new_n930), .A4(new_n962), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(G66));
  NAND3_X1  g781(.A1(new_n569), .A2(G224), .A3(G953), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n862), .B2(G953), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n924), .B1(G898), .B2(new_n260), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n969), .B(new_n970), .Z(G69));
  NOR2_X1   g785(.A1(new_n882), .A2(new_n736), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n800), .A2(new_n668), .A3(new_n701), .A4(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n847), .A2(new_n712), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n973), .A2(new_n820), .A3(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n809), .A2(new_n975), .A3(new_n801), .A4(new_n260), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n540), .A2(new_n541), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n440), .B(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(G900), .B2(G953), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  OR3_X1    g794(.A1(new_n814), .A2(new_n642), .A3(KEYINPUT125), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT125), .B1(new_n814), .B2(new_n642), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n981), .A2(new_n456), .A3(new_n785), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n310), .A2(new_n701), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n705), .A2(new_n974), .A3(new_n707), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT62), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n705), .A2(new_n974), .A3(new_n707), .A4(KEYINPUT62), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n809), .A2(new_n801), .ZN(new_n991));
  AOI21_X1  g805(.A(G953), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n978), .B(KEYINPUT124), .Z(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n980), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n260), .B1(G227), .B2(G900), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n997), .A2(KEYINPUT126), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n995), .A2(new_n999), .A3(new_n996), .ZN(new_n1000));
  AOI21_X1  g814(.A(KEYINPUT127), .B1(new_n995), .B2(new_n996), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n995), .A2(KEYINPUT127), .A3(new_n996), .ZN(new_n1002));
  OAI22_X1  g816(.A1(new_n998), .A2(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(G72));
  INV_X1    g817(.A(new_n422), .ZN(new_n1004));
  NAND2_X1  g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT63), .Z(new_n1006));
  NAND3_X1  g820(.A1(new_n1004), .A2(new_n691), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n876), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n990), .A2(new_n991), .A3(new_n819), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n691), .B1(new_n1009), .B2(new_n1006), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n991), .A2(new_n819), .A3(new_n975), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1004), .B1(new_n1011), .B2(new_n1006), .ZN(new_n1012));
  NOR4_X1   g826(.A1(new_n1008), .A2(new_n1010), .A3(new_n1012), .A4(new_n929), .ZN(G57));
endmodule


