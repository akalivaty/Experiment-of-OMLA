

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592;

  XNOR2_X1 U323 ( .A(n396), .B(n395), .ZN(n541) );
  XNOR2_X1 U324 ( .A(n394), .B(KEYINPUT64), .ZN(n395) );
  XNOR2_X1 U325 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U326 ( .A(n341), .B(n340), .Z(n291) );
  XNOR2_X1 U327 ( .A(KEYINPUT65), .B(KEYINPUT10), .ZN(n347) );
  XNOR2_X1 U328 ( .A(n427), .B(n347), .ZN(n348) );
  XNOR2_X1 U329 ( .A(n389), .B(KEYINPUT47), .ZN(n390) );
  XNOR2_X1 U330 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U331 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U332 ( .A(n356), .B(KEYINPUT9), .ZN(n357) );
  XNOR2_X1 U333 ( .A(n342), .B(n291), .ZN(n343) );
  XNOR2_X1 U334 ( .A(n375), .B(n374), .ZN(n378) );
  XNOR2_X1 U335 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U336 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U337 ( .A(n467), .B(n466), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(G1GAT), .B(KEYINPUT70), .Z(n371) );
  XOR2_X1 U339 ( .A(G15GAT), .B(G50GAT), .Z(n293) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(G36GAT), .ZN(n292) );
  XNOR2_X1 U341 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U342 ( .A(n371), .B(n294), .Z(n296) );
  NAND2_X1 U343 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U345 ( .A(n297), .B(KEYINPUT30), .Z(n300) );
  XNOR2_X1 U346 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n298) );
  XOR2_X1 U347 ( .A(n298), .B(KEYINPUT7), .Z(n361) );
  XOR2_X1 U348 ( .A(n361), .B(KEYINPUT29), .Z(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n308) );
  XOR2_X1 U350 ( .A(G141GAT), .B(G22GAT), .Z(n302) );
  XNOR2_X1 U351 ( .A(G169GAT), .B(G113GAT), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U353 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n304) );
  XNOR2_X1 U354 ( .A(G197GAT), .B(G8GAT), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U356 ( .A(n306), .B(n305), .Z(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n575) );
  XOR2_X1 U358 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n434) );
  XOR2_X1 U359 ( .A(G113GAT), .B(KEYINPUT0), .Z(n439) );
  XOR2_X1 U360 ( .A(G85GAT), .B(G162GAT), .Z(n310) );
  XNOR2_X1 U361 ( .A(G29GAT), .B(G134GAT), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U363 ( .A(n439), .B(n311), .Z(n313) );
  NAND2_X1 U364 ( .A1(G225GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U366 ( .A(n314), .B(KEYINPUT92), .Z(n317) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n315), .B(KEYINPUT2), .ZN(n422) );
  XNOR2_X1 U369 ( .A(n422), .B(KEYINPUT93), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U371 ( .A(G155GAT), .B(G148GAT), .Z(n319) );
  XNOR2_X1 U372 ( .A(G120GAT), .B(G127GAT), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U374 ( .A(n321), .B(n320), .Z(n329) );
  XOR2_X1 U375 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n323) );
  XNOR2_X1 U376 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U378 ( .A(KEYINPUT5), .B(G57GAT), .Z(n325) );
  XNOR2_X1 U379 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n505) );
  INV_X1 U383 ( .A(KEYINPUT54), .ZN(n414) );
  XOR2_X1 U384 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n331) );
  XNOR2_X1 U385 ( .A(G176GAT), .B(KEYINPUT76), .ZN(n330) );
  XOR2_X1 U386 ( .A(n331), .B(n330), .Z(n346) );
  XOR2_X1 U387 ( .A(G64GAT), .B(KEYINPUT71), .Z(n333) );
  XNOR2_X1 U388 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n376) );
  XOR2_X1 U390 ( .A(G120GAT), .B(G71GAT), .Z(n444) );
  XNOR2_X1 U391 ( .A(n376), .B(n444), .ZN(n335) );
  AND2_X1 U392 ( .A1(G230GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n344) );
  XOR2_X1 U394 ( .A(G78GAT), .B(G148GAT), .Z(n337) );
  XNOR2_X1 U395 ( .A(KEYINPUT72), .B(G204GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n421) );
  XOR2_X1 U397 ( .A(G92GAT), .B(G85GAT), .Z(n339) );
  XNOR2_X1 U398 ( .A(G99GAT), .B(G106GAT), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n360) );
  XNOR2_X1 U400 ( .A(n421), .B(n360), .ZN(n342) );
  XOR2_X1 U401 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n341) );
  XNOR2_X1 U402 ( .A(KEYINPUT75), .B(KEYINPUT33), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n384) );
  INV_X1 U404 ( .A(n384), .ZN(n383) );
  XOR2_X1 U405 ( .A(G50GAT), .B(G162GAT), .Z(n427) );
  XOR2_X1 U406 ( .A(G36GAT), .B(G218GAT), .Z(n409) );
  XNOR2_X1 U407 ( .A(n348), .B(n409), .ZN(n352) );
  INV_X1 U408 ( .A(n352), .ZN(n350) );
  AND2_X1 U409 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  INV_X1 U410 ( .A(n351), .ZN(n349) );
  NAND2_X1 U411 ( .A1(n350), .A2(n349), .ZN(n354) );
  NAND2_X1 U412 ( .A1(n352), .A2(n351), .ZN(n353) );
  NAND2_X1 U413 ( .A1(n354), .A2(n353), .ZN(n358) );
  XNOR2_X1 U414 ( .A(G43GAT), .B(G190GAT), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n355), .B(G134GAT), .ZN(n445) );
  XOR2_X1 U416 ( .A(n445), .B(KEYINPUT11), .Z(n356) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n566) );
  XNOR2_X1 U419 ( .A(KEYINPUT77), .B(n566), .ZN(n463) );
  XNOR2_X1 U420 ( .A(KEYINPUT36), .B(n463), .ZN(n588) );
  XOR2_X1 U421 ( .A(G8GAT), .B(G183GAT), .Z(n408) );
  XOR2_X1 U422 ( .A(G22GAT), .B(G155GAT), .Z(n428) );
  XOR2_X1 U423 ( .A(n408), .B(n428), .Z(n364) );
  NAND2_X1 U424 ( .A1(G231GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n369) );
  XOR2_X1 U426 ( .A(G15GAT), .B(G127GAT), .Z(n442) );
  XOR2_X1 U427 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n366) );
  XNOR2_X1 U428 ( .A(G211GAT), .B(KEYINPUT78), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n442), .B(n367), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U432 ( .A(n370), .B(G78GAT), .ZN(n375) );
  XOR2_X1 U433 ( .A(n371), .B(G71GAT), .Z(n373) );
  INV_X1 U434 ( .A(KEYINPUT14), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n376), .B(KEYINPUT12), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n500) );
  NAND2_X1 U437 ( .A1(n588), .A2(n500), .ZN(n380) );
  XNOR2_X1 U438 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n381) );
  INV_X1 U440 ( .A(n575), .ZN(n516) );
  NOR2_X1 U441 ( .A1(n381), .A2(n516), .ZN(n382) );
  NAND2_X1 U442 ( .A1(n383), .A2(n382), .ZN(n393) );
  XOR2_X1 U443 ( .A(n500), .B(KEYINPUT109), .Z(n569) );
  XNOR2_X1 U444 ( .A(n384), .B(KEYINPUT41), .ZN(n559) );
  NOR2_X1 U445 ( .A1(n575), .A2(n559), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n385), .B(KEYINPUT46), .ZN(n386) );
  NOR2_X1 U447 ( .A1(n569), .A2(n386), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n387), .B(KEYINPUT110), .ZN(n388) );
  NAND2_X1 U449 ( .A1(n388), .A2(n566), .ZN(n391) );
  XNOR2_X1 U450 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n389) );
  NAND2_X1 U451 ( .A1(n393), .A2(n392), .ZN(n396) );
  INV_X1 U452 ( .A(KEYINPUT48), .ZN(n394) );
  XOR2_X1 U453 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n398) );
  XNOR2_X1 U454 ( .A(KEYINPUT17), .B(G176GAT), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U456 ( .A(G169GAT), .B(n399), .Z(n452) );
  XOR2_X1 U457 ( .A(G211GAT), .B(KEYINPUT21), .Z(n401) );
  XNOR2_X1 U458 ( .A(G197GAT), .B(KEYINPUT89), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n425) );
  XOR2_X1 U460 ( .A(KEYINPUT94), .B(n425), .Z(n403) );
  NAND2_X1 U461 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U463 ( .A(G64GAT), .B(G92GAT), .Z(n405) );
  XNOR2_X1 U464 ( .A(G190GAT), .B(G204GAT), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U466 ( .A(n407), .B(n406), .Z(n411) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n452), .B(n412), .ZN(n532) );
  NOR2_X1 U470 ( .A1(n541), .A2(n532), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n415) );
  NOR2_X1 U472 ( .A1(n505), .A2(n415), .ZN(n574) );
  XOR2_X1 U473 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n417) );
  XNOR2_X1 U474 ( .A(G218GAT), .B(G106GAT), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n432) );
  XOR2_X1 U476 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n419) );
  NAND2_X1 U477 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U478 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U479 ( .A(n420), .B(KEYINPUT88), .Z(n424) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U482 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U485 ( .A(n432), .B(n431), .Z(n479) );
  NAND2_X1 U486 ( .A1(n574), .A2(n479), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n435), .B(KEYINPUT55), .ZN(n455) );
  XOR2_X1 U489 ( .A(KEYINPUT81), .B(KEYINPUT85), .Z(n437) );
  XNOR2_X1 U490 ( .A(G183GAT), .B(KEYINPUT84), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n438), .B(KEYINPUT20), .Z(n441) );
  XNOR2_X1 U493 ( .A(n439), .B(G99GAT), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U495 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U496 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U497 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U498 ( .A(KEYINPUT83), .B(KEYINPUT80), .Z(n449) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U501 ( .A(n451), .B(n450), .Z(n454) );
  XNOR2_X1 U502 ( .A(n452), .B(KEYINPUT82), .ZN(n453) );
  XNOR2_X1 U503 ( .A(n454), .B(n453), .ZN(n542) );
  NAND2_X1 U504 ( .A1(n455), .A2(n542), .ZN(n462) );
  NOR2_X1 U505 ( .A1(n575), .A2(n462), .ZN(n458) );
  INV_X1 U506 ( .A(KEYINPUT120), .ZN(n456) );
  XNOR2_X1 U507 ( .A(n456), .B(G169GAT), .ZN(n457) );
  XNOR2_X1 U508 ( .A(n458), .B(n457), .ZN(G1348GAT) );
  NOR2_X1 U509 ( .A1(n559), .A2(n462), .ZN(n461) );
  XNOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n459), .B(G176GAT), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  INV_X1 U513 ( .A(n462), .ZN(n570) );
  NAND2_X1 U514 ( .A1(n570), .A2(n463), .ZN(n467) );
  XOR2_X1 U515 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n465) );
  INV_X1 U516 ( .A(G190GAT), .ZN(n464) );
  INV_X1 U517 ( .A(n505), .ZN(n529) );
  NOR2_X1 U518 ( .A1(n384), .A2(n575), .ZN(n503) );
  INV_X1 U519 ( .A(n500), .ZN(n586) );
  NOR2_X1 U520 ( .A1(n463), .A2(n586), .ZN(n468) );
  XNOR2_X1 U521 ( .A(KEYINPUT16), .B(n468), .ZN(n484) );
  NOR2_X1 U522 ( .A1(n479), .A2(n542), .ZN(n469) );
  XNOR2_X1 U523 ( .A(n469), .B(KEYINPUT26), .ZN(n573) );
  XOR2_X1 U524 ( .A(KEYINPUT27), .B(n532), .Z(n477) );
  NAND2_X1 U525 ( .A1(n573), .A2(n477), .ZN(n474) );
  INV_X1 U526 ( .A(n532), .ZN(n509) );
  NAND2_X1 U527 ( .A1(n509), .A2(n542), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n470), .A2(n479), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT25), .ZN(n472) );
  XNOR2_X1 U530 ( .A(KEYINPUT95), .B(n472), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n475), .A2(n529), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n476), .B(KEYINPUT96), .ZN(n483) );
  NAND2_X1 U534 ( .A1(n505), .A2(n477), .ZN(n540) );
  XNOR2_X1 U535 ( .A(KEYINPUT86), .B(n542), .ZN(n478) );
  NOR2_X1 U536 ( .A1(n540), .A2(n478), .ZN(n481) );
  XOR2_X1 U537 ( .A(n479), .B(KEYINPUT67), .Z(n480) );
  XNOR2_X1 U538 ( .A(KEYINPUT28), .B(n480), .ZN(n544) );
  NAND2_X1 U539 ( .A1(n481), .A2(n544), .ZN(n482) );
  NAND2_X1 U540 ( .A1(n483), .A2(n482), .ZN(n498) );
  NAND2_X1 U541 ( .A1(n484), .A2(n498), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n485), .B(KEYINPUT97), .ZN(n517) );
  NAND2_X1 U543 ( .A1(n503), .A2(n517), .ZN(n496) );
  NOR2_X1 U544 ( .A1(n529), .A2(n496), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT34), .B(KEYINPUT98), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U547 ( .A(G1GAT), .B(n488), .Z(G1324GAT) );
  NOR2_X1 U548 ( .A1(n532), .A2(n496), .ZN(n490) );
  XNOR2_X1 U549 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G8GAT), .B(n491), .ZN(G1325GAT) );
  INV_X1 U552 ( .A(n542), .ZN(n535) );
  NOR2_X1 U553 ( .A1(n496), .A2(n535), .ZN(n495) );
  XOR2_X1 U554 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n493) );
  XNOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NOR2_X1 U558 ( .A1(n544), .A2(n496), .ZN(n497) );
  XOR2_X1 U559 ( .A(G22GAT), .B(n497), .Z(G1327GAT) );
  NAND2_X1 U560 ( .A1(n588), .A2(n498), .ZN(n499) );
  NOR2_X1 U561 ( .A1(n500), .A2(n499), .ZN(n501) );
  XOR2_X1 U562 ( .A(n501), .B(KEYINPUT104), .Z(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT37), .B(n502), .ZN(n527) );
  NAND2_X1 U564 ( .A1(n527), .A2(n503), .ZN(n504) );
  XOR2_X1 U565 ( .A(KEYINPUT38), .B(n504), .Z(n513) );
  NAND2_X1 U566 ( .A1(n513), .A2(n505), .ZN(n508) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n506), .B(KEYINPUT39), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n508), .B(n507), .ZN(G1328GAT) );
  NAND2_X1 U570 ( .A1(n513), .A2(n509), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n510), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U572 ( .A1(n513), .A2(n542), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(KEYINPUT40), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G43GAT), .B(n512), .ZN(G1330GAT) );
  INV_X1 U575 ( .A(n544), .ZN(n514) );
  NAND2_X1 U576 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U577 ( .A(G50GAT), .B(n515), .ZN(G1331GAT) );
  NOR2_X1 U578 ( .A1(n516), .A2(n559), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n517), .A2(n528), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n529), .A2(n523), .ZN(n518) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n518), .Z(n519) );
  XNOR2_X1 U582 ( .A(KEYINPUT42), .B(n519), .ZN(G1332GAT) );
  NOR2_X1 U583 ( .A1(n532), .A2(n523), .ZN(n521) );
  XNOR2_X1 U584 ( .A(G64GAT), .B(KEYINPUT105), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(G1333GAT) );
  NOR2_X1 U586 ( .A1(n535), .A2(n523), .ZN(n522) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n522), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n544), .A2(n523), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G78GAT), .B(n526), .ZN(G1335GAT) );
  NAND2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n537) );
  NOR2_X1 U593 ( .A1(n529), .A2(n537), .ZN(n531) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1336GAT) );
  NOR2_X1 U596 ( .A1(n532), .A2(n537), .ZN(n533) );
  XOR2_X1 U597 ( .A(KEYINPUT108), .B(n533), .Z(n534) );
  XNOR2_X1 U598 ( .A(G92GAT), .B(n534), .ZN(G1337GAT) );
  NOR2_X1 U599 ( .A1(n535), .A2(n537), .ZN(n536) );
  XOR2_X1 U600 ( .A(G99GAT), .B(n536), .Z(G1338GAT) );
  NOR2_X1 U601 ( .A1(n544), .A2(n537), .ZN(n538) );
  XOR2_X1 U602 ( .A(KEYINPUT44), .B(n538), .Z(n539) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  NOR2_X1 U604 ( .A1(n541), .A2(n540), .ZN(n557) );
  NAND2_X1 U605 ( .A1(n542), .A2(n557), .ZN(n543) );
  XNOR2_X1 U606 ( .A(n543), .B(KEYINPUT113), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n550) );
  NOR2_X1 U608 ( .A1(n575), .A2(n550), .ZN(n546) );
  XOR2_X1 U609 ( .A(n546), .B(KEYINPUT114), .Z(n547) );
  XNOR2_X1 U610 ( .A(G113GAT), .B(n547), .ZN(G1340GAT) );
  NOR2_X1 U611 ( .A1(n559), .A2(n550), .ZN(n549) );
  XNOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  INV_X1 U614 ( .A(n550), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n553), .A2(n569), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n551), .B(KEYINPUT50), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n552), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U619 ( .A1(n553), .A2(n463), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U621 ( .A(G134GAT), .B(n556), .Z(G1343GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n573), .ZN(n565) );
  NOR2_X1 U623 ( .A1(n575), .A2(n565), .ZN(n558) );
  XOR2_X1 U624 ( .A(G141GAT), .B(n558), .Z(G1344GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n565), .ZN(n561) );
  XNOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U629 ( .A1(n586), .A2(n565), .ZN(n563) );
  XOR2_X1 U630 ( .A(KEYINPUT116), .B(n563), .Z(n564) );
  XNOR2_X1 U631 ( .A(G155GAT), .B(n564), .ZN(G1346GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1347GAT) );
  XOR2_X1 U635 ( .A(G183GAT), .B(KEYINPUT121), .Z(n572) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1350GAT) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n585) );
  NOR2_X1 U639 ( .A1(n575), .A2(n585), .ZN(n580) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n577) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(KEYINPUT59), .B(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  INV_X1 U645 ( .A(n585), .ZN(n589) );
  AND2_X1 U646 ( .A1(n589), .A2(n384), .ZN(n584) );
  XOR2_X1 U647 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n582) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n587), .Z(G1354GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n591) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

