

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U554 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  OR2_X1 U555 ( .A1(n606), .A2(n605), .ZN(n619) );
  OR2_X1 U556 ( .A1(n638), .A2(n961), .ZN(n637) );
  INV_X1 U557 ( .A(KEYINPUT105), .ZN(n680) );
  OR2_X1 U558 ( .A1(G2105), .A2(n521), .ZN(n522) );
  XOR2_X2 U559 ( .A(KEYINPUT17), .B(n520), .Z(n893) );
  INV_X1 U560 ( .A(KEYINPUT29), .ZN(n648) );
  NAND2_X1 U561 ( .A1(n593), .A2(n687), .ZN(n604) );
  BUF_X1 U562 ( .A(n604), .Z(n668) );
  NOR2_X2 U563 ( .A1(G543), .A2(G651), .ZN(n799) );
  INV_X1 U564 ( .A(KEYINPUT109), .ZN(n757) );
  NOR2_X1 U565 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U566 ( .A1(G2105), .A2(n530), .ZN(n892) );
  XNOR2_X1 U567 ( .A(n758), .B(n757), .ZN(n772) );
  NOR2_X1 U568 ( .A1(n529), .A2(n528), .ZN(G160) );
  NAND2_X1 U569 ( .A1(n893), .A2(G137), .ZN(n525) );
  INV_X1 U570 ( .A(KEYINPUT23), .ZN(n523) );
  NAND2_X1 U571 ( .A1(G2104), .A2(G101), .ZN(n521) );
  XNOR2_X1 U572 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n529) );
  INV_X1 U574 ( .A(G2104), .ZN(n530) );
  AND2_X1 U575 ( .A1(n530), .A2(G2105), .ZN(n888) );
  NAND2_X1 U576 ( .A1(G125), .A2(n888), .ZN(n527) );
  AND2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n889) );
  NAND2_X1 U578 ( .A1(G113), .A2(n889), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U580 ( .A1(G102), .A2(n892), .ZN(n532) );
  NAND2_X1 U581 ( .A1(G138), .A2(n893), .ZN(n531) );
  NAND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n536) );
  NAND2_X1 U583 ( .A1(G126), .A2(n888), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G114), .A2(n889), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U586 ( .A1(n536), .A2(n535), .ZN(G164) );
  INV_X1 U587 ( .A(G651), .ZN(n544) );
  NOR2_X1 U588 ( .A1(G543), .A2(n544), .ZN(n537) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n537), .Z(n607) );
  BUF_X1 U590 ( .A(n607), .Z(n803) );
  NAND2_X1 U591 ( .A1(n803), .A2(G63), .ZN(n538) );
  XNOR2_X1 U592 ( .A(n538), .B(KEYINPUT78), .ZN(n541) );
  XOR2_X1 U593 ( .A(G543), .B(KEYINPUT0), .Z(n539) );
  XNOR2_X1 U594 ( .A(KEYINPUT66), .B(n539), .ZN(n573) );
  NOR2_X1 U595 ( .A1(G651), .A2(n573), .ZN(n623) );
  BUF_X1 U596 ( .A(n623), .Z(n804) );
  NAND2_X1 U597 ( .A1(G51), .A2(n804), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U599 ( .A(KEYINPUT6), .B(n542), .ZN(n550) );
  NAND2_X1 U600 ( .A1(n799), .A2(G89), .ZN(n543) );
  XNOR2_X1 U601 ( .A(n543), .B(KEYINPUT4), .ZN(n546) );
  NOR2_X1 U602 ( .A1(n573), .A2(n544), .ZN(n624) );
  BUF_X1 U603 ( .A(n624), .Z(n800) );
  NAND2_X1 U604 ( .A1(G76), .A2(n800), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U606 ( .A(KEYINPUT5), .B(n547), .ZN(n548) );
  XNOR2_X1 U607 ( .A(KEYINPUT77), .B(n548), .ZN(n549) );
  NOR2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U609 ( .A(KEYINPUT7), .B(n551), .Z(G168) );
  XOR2_X1 U610 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U611 ( .A1(n800), .A2(G77), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n552), .B(KEYINPUT68), .ZN(n554) );
  NAND2_X1 U613 ( .A1(G90), .A2(n799), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n556) );
  XOR2_X1 U615 ( .A(KEYINPUT9), .B(KEYINPUT69), .Z(n555) );
  XNOR2_X1 U616 ( .A(n556), .B(n555), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G64), .A2(n803), .ZN(n558) );
  NAND2_X1 U618 ( .A1(G52), .A2(n804), .ZN(n557) );
  AND2_X1 U619 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(G301) );
  INV_X1 U621 ( .A(G301), .ZN(G171) );
  NAND2_X1 U622 ( .A1(n800), .A2(G75), .ZN(n561) );
  XNOR2_X1 U623 ( .A(n561), .B(KEYINPUT86), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G88), .A2(n799), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U626 ( .A(KEYINPUT87), .B(n564), .ZN(n568) );
  NAND2_X1 U627 ( .A1(G62), .A2(n803), .ZN(n566) );
  NAND2_X1 U628 ( .A1(G50), .A2(n804), .ZN(n565) );
  AND2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n568), .A2(n567), .ZN(G303) );
  NAND2_X1 U631 ( .A1(G49), .A2(n804), .ZN(n570) );
  NAND2_X1 U632 ( .A1(G74), .A2(G651), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U634 ( .A1(n803), .A2(n571), .ZN(n572) );
  XOR2_X1 U635 ( .A(KEYINPUT83), .B(n572), .Z(n575) );
  NAND2_X1 U636 ( .A1(G87), .A2(n573), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(G288) );
  NAND2_X1 U638 ( .A1(G73), .A2(n800), .ZN(n576) );
  XNOR2_X1 U639 ( .A(n576), .B(KEYINPUT2), .ZN(n584) );
  NAND2_X1 U640 ( .A1(G61), .A2(n803), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G86), .A2(n799), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT84), .B(n579), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G48), .A2(n804), .ZN(n580) );
  XNOR2_X1 U645 ( .A(KEYINPUT85), .B(n580), .ZN(n581) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U647 ( .A1(n584), .A2(n583), .ZN(G305) );
  NAND2_X1 U648 ( .A1(n804), .A2(G47), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n803), .A2(G60), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT67), .B(n587), .Z(n590) );
  NAND2_X1 U652 ( .A1(G85), .A2(n799), .ZN(n588) );
  XNOR2_X1 U653 ( .A(KEYINPUT65), .B(n588), .ZN(n589) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U655 ( .A1(n800), .A2(G72), .ZN(n591) );
  NAND2_X1 U656 ( .A1(n592), .A2(n591), .ZN(G290) );
  NAND2_X1 U657 ( .A1(G160), .A2(G40), .ZN(n686) );
  INV_X1 U658 ( .A(n686), .ZN(n593) );
  NOR2_X2 U659 ( .A1(G164), .A2(G1384), .ZN(n687) );
  INV_X1 U660 ( .A(n668), .ZN(n651) );
  NAND2_X1 U661 ( .A1(n651), .A2(G2072), .ZN(n594) );
  XNOR2_X1 U662 ( .A(n594), .B(KEYINPUT27), .ZN(n596) );
  INV_X1 U663 ( .A(G1956), .ZN(n997) );
  NOR2_X1 U664 ( .A1(n997), .A2(n651), .ZN(n595) );
  NOR2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n644) );
  NAND2_X1 U666 ( .A1(G65), .A2(n803), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G53), .A2(n804), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U669 ( .A1(G91), .A2(n799), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G78), .A2(n800), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n964) );
  NAND2_X1 U673 ( .A1(n644), .A2(n964), .ZN(n643) );
  INV_X1 U674 ( .A(G1996), .ZN(n936) );
  NOR2_X1 U675 ( .A1(n604), .A2(n936), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n603), .B(KEYINPUT26), .ZN(n606) );
  AND2_X1 U677 ( .A1(n604), .A2(G1341), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n607), .A2(G56), .ZN(n608) );
  XOR2_X1 U679 ( .A(n608), .B(KEYINPUT14), .Z(n615) );
  INV_X1 U680 ( .A(KEYINPUT13), .ZN(n613) );
  NAND2_X1 U681 ( .A1(n799), .A2(G81), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n609), .B(KEYINPUT12), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G68), .A2(n624), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n616), .B(KEYINPUT74), .ZN(n618) );
  NAND2_X1 U687 ( .A1(G43), .A2(n804), .ZN(n617) );
  NAND2_X1 U688 ( .A1(n618), .A2(n617), .ZN(n976) );
  NOR2_X1 U689 ( .A1(n619), .A2(n976), .ZN(n620) );
  XOR2_X1 U690 ( .A(n620), .B(KEYINPUT64), .Z(n638) );
  INV_X1 U691 ( .A(KEYINPUT15), .ZN(n632) );
  NAND2_X1 U692 ( .A1(G66), .A2(n803), .ZN(n622) );
  NAND2_X1 U693 ( .A1(G92), .A2(n799), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n630) );
  NAND2_X1 U695 ( .A1(G54), .A2(n623), .ZN(n626) );
  NAND2_X1 U696 ( .A1(G79), .A2(n624), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n628) );
  INV_X1 U698 ( .A(KEYINPUT75), .ZN(n627) );
  XNOR2_X1 U699 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X1 U700 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U702 ( .A(KEYINPUT76), .B(n633), .ZN(n818) );
  INV_X1 U703 ( .A(n818), .ZN(n961) );
  NOR2_X1 U704 ( .A1(n651), .A2(G1348), .ZN(n635) );
  NOR2_X1 U705 ( .A1(G2067), .A2(n668), .ZN(n634) );
  NOR2_X1 U706 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U708 ( .A1(n961), .A2(n638), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U710 ( .A(KEYINPUT101), .B(n641), .Z(n642) );
  NAND2_X1 U711 ( .A1(n643), .A2(n642), .ZN(n647) );
  NOR2_X1 U712 ( .A1(n644), .A2(n964), .ZN(n645) );
  XOR2_X1 U713 ( .A(n645), .B(KEYINPUT28), .Z(n646) );
  NAND2_X1 U714 ( .A1(n647), .A2(n646), .ZN(n649) );
  XNOR2_X1 U715 ( .A(n649), .B(n648), .ZN(n655) );
  NOR2_X1 U716 ( .A1(n651), .A2(G1961), .ZN(n650) );
  XOR2_X1 U717 ( .A(KEYINPUT100), .B(n650), .Z(n653) );
  XNOR2_X1 U718 ( .A(G2078), .B(KEYINPUT25), .ZN(n937) );
  NAND2_X1 U719 ( .A1(n651), .A2(n937), .ZN(n652) );
  NAND2_X1 U720 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U721 ( .A1(n656), .A2(G171), .ZN(n654) );
  NAND2_X1 U722 ( .A1(n655), .A2(n654), .ZN(n667) );
  NOR2_X1 U723 ( .A1(G171), .A2(n656), .ZN(n657) );
  XOR2_X1 U724 ( .A(KEYINPUT103), .B(n657), .Z(n663) );
  NOR2_X1 U725 ( .A1(G2084), .A2(n668), .ZN(n682) );
  NAND2_X1 U726 ( .A1(G8), .A2(n668), .ZN(n737) );
  NOR2_X1 U727 ( .A1(G1966), .A2(n737), .ZN(n679) );
  NOR2_X1 U728 ( .A1(n682), .A2(n679), .ZN(n658) );
  NAND2_X1 U729 ( .A1(G8), .A2(n658), .ZN(n659) );
  XNOR2_X1 U730 ( .A(KEYINPUT30), .B(n659), .ZN(n660) );
  NOR2_X1 U731 ( .A1(G168), .A2(n660), .ZN(n661) );
  XNOR2_X1 U732 ( .A(KEYINPUT102), .B(n661), .ZN(n662) );
  NOR2_X1 U733 ( .A1(n663), .A2(n662), .ZN(n665) );
  XOR2_X1 U734 ( .A(KEYINPUT104), .B(KEYINPUT31), .Z(n664) );
  XNOR2_X1 U735 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n677) );
  NAND2_X1 U737 ( .A1(G286), .A2(n677), .ZN(n673) );
  NOR2_X1 U738 ( .A1(G1971), .A2(n737), .ZN(n670) );
  NOR2_X1 U739 ( .A1(G2090), .A2(n668), .ZN(n669) );
  NOR2_X1 U740 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U741 ( .A1(n671), .A2(G303), .ZN(n672) );
  NAND2_X1 U742 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U743 ( .A(n674), .B(KEYINPUT106), .ZN(n675) );
  NAND2_X1 U744 ( .A1(n675), .A2(G8), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n676), .B(KEYINPUT32), .ZN(n740) );
  INV_X1 U746 ( .A(n677), .ZN(n678) );
  NOR2_X1 U747 ( .A1(n679), .A2(n678), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n681), .B(n680), .ZN(n684) );
  NAND2_X1 U749 ( .A1(G8), .A2(n682), .ZN(n683) );
  NAND2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n738) );
  NAND2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n966) );
  AND2_X1 U752 ( .A1(n738), .A2(n966), .ZN(n719) );
  NOR2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n723) );
  NAND2_X1 U754 ( .A1(n723), .A2(KEYINPUT33), .ZN(n685) );
  NOR2_X1 U755 ( .A1(n685), .A2(n737), .ZN(n718) );
  XOR2_X1 U756 ( .A(G1981), .B(G305), .Z(n958) );
  NOR2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n769) );
  XNOR2_X1 U758 ( .A(G2067), .B(KEYINPUT37), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT94), .ZN(n767) );
  NAND2_X1 U760 ( .A1(G104), .A2(n892), .ZN(n690) );
  NAND2_X1 U761 ( .A1(G140), .A2(n893), .ZN(n689) );
  NAND2_X1 U762 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U763 ( .A(KEYINPUT34), .B(n691), .ZN(n696) );
  NAND2_X1 U764 ( .A1(G128), .A2(n888), .ZN(n693) );
  NAND2_X1 U765 ( .A1(G116), .A2(n889), .ZN(n692) );
  NAND2_X1 U766 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U767 ( .A(KEYINPUT35), .B(n694), .Z(n695) );
  NOR2_X1 U768 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U769 ( .A(KEYINPUT36), .B(n697), .ZN(n910) );
  NOR2_X1 U770 ( .A1(n767), .A2(n910), .ZN(n1018) );
  NAND2_X1 U771 ( .A1(n769), .A2(n1018), .ZN(n765) );
  NAND2_X1 U772 ( .A1(G119), .A2(n888), .ZN(n699) );
  NAND2_X1 U773 ( .A1(G131), .A2(n893), .ZN(n698) );
  NAND2_X1 U774 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U775 ( .A1(G95), .A2(n892), .ZN(n701) );
  NAND2_X1 U776 ( .A1(G107), .A2(n889), .ZN(n700) );
  NAND2_X1 U777 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U778 ( .A1(n703), .A2(n702), .ZN(n901) );
  INV_X1 U779 ( .A(G1991), .ZN(n759) );
  NOR2_X1 U780 ( .A1(n901), .A2(n759), .ZN(n713) );
  NAND2_X1 U781 ( .A1(G105), .A2(n892), .ZN(n704) );
  XOR2_X1 U782 ( .A(KEYINPUT38), .B(n704), .Z(n709) );
  NAND2_X1 U783 ( .A1(G129), .A2(n888), .ZN(n706) );
  NAND2_X1 U784 ( .A1(G117), .A2(n889), .ZN(n705) );
  NAND2_X1 U785 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U786 ( .A(KEYINPUT95), .B(n707), .Z(n708) );
  NOR2_X1 U787 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U788 ( .A1(n893), .A2(G141), .ZN(n710) );
  NAND2_X1 U789 ( .A1(n711), .A2(n710), .ZN(n887) );
  AND2_X1 U790 ( .A1(n887), .A2(G1996), .ZN(n712) );
  NOR2_X1 U791 ( .A1(n713), .A2(n712), .ZN(n1020) );
  XOR2_X1 U792 ( .A(n769), .B(KEYINPUT96), .Z(n714) );
  NOR2_X1 U793 ( .A1(n1020), .A2(n714), .ZN(n762) );
  INV_X1 U794 ( .A(n762), .ZN(n715) );
  NAND2_X1 U795 ( .A1(n765), .A2(n715), .ZN(n716) );
  XNOR2_X1 U796 ( .A(KEYINPUT97), .B(n716), .ZN(n751) );
  NAND2_X1 U797 ( .A1(n958), .A2(n751), .ZN(n717) );
  NOR2_X1 U798 ( .A1(n718), .A2(n717), .ZN(n721) );
  AND2_X1 U799 ( .A1(n719), .A2(n721), .ZN(n720) );
  NAND2_X1 U800 ( .A1(n740), .A2(n720), .ZN(n732) );
  INV_X1 U801 ( .A(n721), .ZN(n730) );
  INV_X1 U802 ( .A(KEYINPUT33), .ZN(n728) );
  INV_X1 U803 ( .A(n966), .ZN(n725) );
  NOR2_X1 U804 ( .A1(G1971), .A2(G303), .ZN(n722) );
  NOR2_X1 U805 ( .A1(n723), .A2(n722), .ZN(n971) );
  XOR2_X1 U806 ( .A(n971), .B(KEYINPUT107), .Z(n724) );
  OR2_X1 U807 ( .A1(n725), .A2(n724), .ZN(n726) );
  OR2_X1 U808 ( .A1(n737), .A2(n726), .ZN(n727) );
  AND2_X1 U809 ( .A1(n728), .A2(n727), .ZN(n729) );
  OR2_X1 U810 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U811 ( .A1(n732), .A2(n731), .ZN(n753) );
  NOR2_X1 U812 ( .A1(G1981), .A2(G305), .ZN(n733) );
  XOR2_X1 U813 ( .A(n733), .B(KEYINPUT98), .Z(n734) );
  XNOR2_X1 U814 ( .A(KEYINPUT24), .B(n734), .ZN(n735) );
  NOR2_X1 U815 ( .A1(n737), .A2(n735), .ZN(n736) );
  XOR2_X1 U816 ( .A(KEYINPUT99), .B(n736), .Z(n743) );
  OR2_X1 U817 ( .A1(n743), .A2(n737), .ZN(n741) );
  AND2_X1 U818 ( .A1(n738), .A2(n741), .ZN(n739) );
  NAND2_X1 U819 ( .A1(n740), .A2(n739), .ZN(n749) );
  INV_X1 U820 ( .A(n741), .ZN(n747) );
  NOR2_X1 U821 ( .A1(G2090), .A2(G303), .ZN(n742) );
  NAND2_X1 U822 ( .A1(G8), .A2(n742), .ZN(n745) );
  INV_X1 U823 ( .A(n743), .ZN(n744) );
  AND2_X1 U824 ( .A1(n745), .A2(n744), .ZN(n746) );
  OR2_X1 U825 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U826 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U827 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U828 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U829 ( .A(n754), .B(KEYINPUT108), .ZN(n756) );
  XNOR2_X1 U830 ( .A(G1986), .B(G290), .ZN(n973) );
  NAND2_X1 U831 ( .A1(n769), .A2(n973), .ZN(n755) );
  NAND2_X1 U832 ( .A1(n756), .A2(n755), .ZN(n758) );
  NOR2_X1 U833 ( .A1(G1996), .A2(n887), .ZN(n1028) );
  AND2_X1 U834 ( .A1(n759), .A2(n901), .ZN(n1014) );
  NOR2_X1 U835 ( .A1(G1986), .A2(G290), .ZN(n760) );
  NOR2_X1 U836 ( .A1(n1014), .A2(n760), .ZN(n761) );
  NOR2_X1 U837 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U838 ( .A1(n1028), .A2(n763), .ZN(n764) );
  XNOR2_X1 U839 ( .A(n764), .B(KEYINPUT39), .ZN(n766) );
  NAND2_X1 U840 ( .A1(n766), .A2(n765), .ZN(n768) );
  NAND2_X1 U841 ( .A1(n767), .A2(n910), .ZN(n1032) );
  NAND2_X1 U842 ( .A1(n768), .A2(n1032), .ZN(n770) );
  NAND2_X1 U843 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U844 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U845 ( .A(n773), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U846 ( .A(G132), .ZN(G219) );
  INV_X1 U847 ( .A(G82), .ZN(G220) );
  INV_X1 U848 ( .A(G120), .ZN(G236) );
  INV_X1 U849 ( .A(G69), .ZN(G235) );
  NAND2_X1 U850 ( .A1(G94), .A2(G452), .ZN(n774) );
  XOR2_X1 U851 ( .A(KEYINPUT70), .B(n774), .Z(G173) );
  NAND2_X1 U852 ( .A1(G7), .A2(G661), .ZN(n775) );
  XNOR2_X1 U853 ( .A(n775), .B(KEYINPUT10), .ZN(n776) );
  XNOR2_X1 U854 ( .A(KEYINPUT72), .B(n776), .ZN(G223) );
  XNOR2_X1 U855 ( .A(KEYINPUT73), .B(G223), .ZN(n840) );
  NAND2_X1 U856 ( .A1(n840), .A2(G567), .ZN(n777) );
  XOR2_X1 U857 ( .A(KEYINPUT11), .B(n777), .Z(G234) );
  INV_X1 U858 ( .A(G860), .ZN(n783) );
  OR2_X1 U859 ( .A1(n976), .A2(n783), .ZN(G153) );
  NOR2_X1 U860 ( .A1(n961), .A2(G868), .ZN(n779) );
  INV_X1 U861 ( .A(G868), .ZN(n780) );
  NOR2_X1 U862 ( .A1(n780), .A2(G301), .ZN(n778) );
  NOR2_X1 U863 ( .A1(n779), .A2(n778), .ZN(G284) );
  INV_X1 U864 ( .A(n964), .ZN(G299) );
  NOR2_X1 U865 ( .A1(G286), .A2(n780), .ZN(n782) );
  NOR2_X1 U866 ( .A1(G868), .A2(G299), .ZN(n781) );
  NOR2_X1 U867 ( .A1(n782), .A2(n781), .ZN(G297) );
  NAND2_X1 U868 ( .A1(n783), .A2(G559), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n784), .A2(n818), .ZN(n785) );
  XNOR2_X1 U870 ( .A(n785), .B(KEYINPUT79), .ZN(n786) );
  XOR2_X1 U871 ( .A(KEYINPUT16), .B(n786), .Z(G148) );
  NOR2_X1 U872 ( .A1(G868), .A2(n976), .ZN(n789) );
  NAND2_X1 U873 ( .A1(n818), .A2(G868), .ZN(n787) );
  NOR2_X1 U874 ( .A1(G559), .A2(n787), .ZN(n788) );
  NOR2_X1 U875 ( .A1(n789), .A2(n788), .ZN(G282) );
  NAND2_X1 U876 ( .A1(G123), .A2(n888), .ZN(n790) );
  XNOR2_X1 U877 ( .A(n790), .B(KEYINPUT18), .ZN(n792) );
  NAND2_X1 U878 ( .A1(n892), .A2(G99), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G135), .A2(n893), .ZN(n794) );
  NAND2_X1 U881 ( .A1(G111), .A2(n889), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n1013) );
  XNOR2_X1 U884 ( .A(n1013), .B(G2096), .ZN(n798) );
  INV_X1 U885 ( .A(G2100), .ZN(n797) );
  NAND2_X1 U886 ( .A1(n798), .A2(n797), .ZN(G156) );
  NAND2_X1 U887 ( .A1(G93), .A2(n799), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G80), .A2(n800), .ZN(n801) );
  NAND2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n809) );
  NAND2_X1 U890 ( .A1(G67), .A2(n803), .ZN(n806) );
  NAND2_X1 U891 ( .A1(G55), .A2(n804), .ZN(n805) );
  NAND2_X1 U892 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U893 ( .A(KEYINPUT81), .B(n807), .Z(n808) );
  NOR2_X1 U894 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U895 ( .A(KEYINPUT82), .B(n810), .ZN(n848) );
  NOR2_X1 U896 ( .A1(G868), .A2(n848), .ZN(n811) );
  XNOR2_X1 U897 ( .A(n811), .B(KEYINPUT89), .ZN(n823) );
  INV_X1 U898 ( .A(n848), .ZN(n812) );
  XNOR2_X1 U899 ( .A(n812), .B(G290), .ZN(n813) );
  XNOR2_X1 U900 ( .A(n813), .B(G288), .ZN(n814) );
  XNOR2_X1 U901 ( .A(KEYINPUT19), .B(n814), .ZN(n816) );
  XNOR2_X1 U902 ( .A(G305), .B(n964), .ZN(n815) );
  XNOR2_X1 U903 ( .A(n816), .B(n815), .ZN(n817) );
  XNOR2_X1 U904 ( .A(n817), .B(G303), .ZN(n913) );
  XNOR2_X1 U905 ( .A(n913), .B(KEYINPUT88), .ZN(n820) );
  NAND2_X1 U906 ( .A1(n818), .A2(G559), .ZN(n819) );
  XNOR2_X1 U907 ( .A(n819), .B(n976), .ZN(n846) );
  XNOR2_X1 U908 ( .A(n820), .B(n846), .ZN(n821) );
  NAND2_X1 U909 ( .A1(G868), .A2(n821), .ZN(n822) );
  NAND2_X1 U910 ( .A1(n823), .A2(n822), .ZN(G295) );
  NAND2_X1 U911 ( .A1(G2084), .A2(G2078), .ZN(n824) );
  XOR2_X1 U912 ( .A(KEYINPUT20), .B(n824), .Z(n825) );
  NAND2_X1 U913 ( .A1(G2090), .A2(n825), .ZN(n826) );
  XNOR2_X1 U914 ( .A(KEYINPUT21), .B(n826), .ZN(n827) );
  NAND2_X1 U915 ( .A1(n827), .A2(G2072), .ZN(n828) );
  XNOR2_X1 U916 ( .A(KEYINPUT90), .B(n828), .ZN(G158) );
  XNOR2_X1 U917 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  XNOR2_X1 U918 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U919 ( .A1(G235), .A2(G236), .ZN(n829) );
  XOR2_X1 U920 ( .A(KEYINPUT92), .B(n829), .Z(n830) );
  NOR2_X1 U921 ( .A1(G237), .A2(n830), .ZN(n831) );
  NAND2_X1 U922 ( .A1(G108), .A2(n831), .ZN(n850) );
  NAND2_X1 U923 ( .A1(G567), .A2(n850), .ZN(n832) );
  XOR2_X1 U924 ( .A(KEYINPUT93), .B(n832), .Z(n838) );
  NOR2_X1 U925 ( .A1(G220), .A2(G219), .ZN(n833) );
  XOR2_X1 U926 ( .A(KEYINPUT22), .B(n833), .Z(n834) );
  NOR2_X1 U927 ( .A1(G218), .A2(n834), .ZN(n835) );
  NAND2_X1 U928 ( .A1(G96), .A2(n835), .ZN(n851) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n851), .ZN(n836) );
  XOR2_X1 U930 ( .A(KEYINPUT91), .B(n836), .Z(n837) );
  NAND2_X1 U931 ( .A1(n838), .A2(n837), .ZN(n852) );
  NAND2_X1 U932 ( .A1(G483), .A2(G661), .ZN(n839) );
  NOR2_X1 U933 ( .A1(n852), .A2(n839), .ZN(n845) );
  NAND2_X1 U934 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n840), .ZN(G217) );
  INV_X1 U936 ( .A(G661), .ZN(n842) );
  NAND2_X1 U937 ( .A1(G2), .A2(G15), .ZN(n841) );
  NOR2_X1 U938 ( .A1(n842), .A2(n841), .ZN(n843) );
  XOR2_X1 U939 ( .A(KEYINPUT110), .B(n843), .Z(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U941 ( .A1(n845), .A2(n844), .ZN(G188) );
  XNOR2_X1 U943 ( .A(KEYINPUT80), .B(n846), .ZN(n847) );
  NOR2_X1 U944 ( .A1(G860), .A2(n847), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(G145) );
  INV_X1 U946 ( .A(G108), .ZN(G238) );
  INV_X1 U947 ( .A(G96), .ZN(G221) );
  NOR2_X1 U948 ( .A1(n851), .A2(n850), .ZN(G325) );
  INV_X1 U949 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U950 ( .A(KEYINPUT111), .B(n852), .ZN(G319) );
  XOR2_X1 U951 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n854) );
  XNOR2_X1 U952 ( .A(G2678), .B(KEYINPUT43), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(G2090), .Z(n856) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U957 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U958 ( .A(G2096), .B(G2100), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n862) );
  XOR2_X1 U960 ( .A(G2084), .B(G2078), .Z(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(G227) );
  XOR2_X1 U962 ( .A(G1971), .B(G1961), .Z(n864) );
  XNOR2_X1 U963 ( .A(G1976), .B(G1966), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(n865), .B(KEYINPUT41), .Z(n867) );
  XNOR2_X1 U966 ( .A(G1996), .B(G1991), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U968 ( .A(G2474), .B(G1956), .Z(n869) );
  XNOR2_X1 U969 ( .A(G1986), .B(G1981), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U972 ( .A1(G124), .A2(n888), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n872), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n892), .A2(G100), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G136), .A2(n893), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G112), .A2(n889), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U979 ( .A1(n878), .A2(n877), .ZN(G162) );
  NAND2_X1 U980 ( .A1(G127), .A2(n888), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G115), .A2(n889), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n881), .B(KEYINPUT47), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G139), .A2(n893), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n892), .A2(G103), .ZN(n884) );
  XOR2_X1 U987 ( .A(KEYINPUT114), .B(n884), .Z(n885) );
  NOR2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n1021) );
  XOR2_X1 U989 ( .A(n887), .B(n1021), .Z(n909) );
  NAND2_X1 U990 ( .A1(G130), .A2(n888), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G118), .A2(n889), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n898) );
  NAND2_X1 U993 ( .A1(G106), .A2(n892), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G142), .A2(n893), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U996 ( .A(KEYINPUT45), .B(n896), .Z(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n905) );
  XNOR2_X1 U998 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n899), .B(KEYINPUT46), .ZN(n900) );
  XOR2_X1 U1000 ( .A(n900), .B(n1013), .Z(n903) );
  XNOR2_X1 U1001 ( .A(G164), .B(n901), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1003 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1004 ( .A(G160), .B(G162), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n911) );
  XOR2_X1 U1007 ( .A(n911), .B(n910), .Z(n912) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n912), .ZN(G395) );
  XOR2_X1 U1009 ( .A(n913), .B(G286), .Z(n915) );
  XNOR2_X1 U1010 ( .A(G171), .B(n961), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1012 ( .A(n916), .B(n976), .Z(n917) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n917), .ZN(G397) );
  XOR2_X1 U1014 ( .A(G2451), .B(G2430), .Z(n919) );
  XNOR2_X1 U1015 ( .A(G2438), .B(G2443), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(n925) );
  XOR2_X1 U1017 ( .A(G2435), .B(G2454), .Z(n921) );
  XNOR2_X1 U1018 ( .A(G1341), .B(G1348), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(n921), .B(n920), .ZN(n923) );
  XOR2_X1 U1020 ( .A(G2446), .B(G2427), .Z(n922) );
  XNOR2_X1 U1021 ( .A(n923), .B(n922), .ZN(n924) );
  XOR2_X1 U1022 ( .A(n925), .B(n924), .Z(n926) );
  NAND2_X1 U1023 ( .A1(G14), .A2(n926), .ZN(n932) );
  NAND2_X1 U1024 ( .A1(G319), .A2(n932), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(G227), .A2(G229), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(KEYINPUT49), .B(n927), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(G395), .A2(G397), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(G225) );
  INV_X1 U1030 ( .A(G225), .ZN(G308) );
  INV_X1 U1031 ( .A(G303), .ZN(G166) );
  INV_X1 U1032 ( .A(n932), .ZN(G401) );
  XOR2_X1 U1033 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n1043) );
  INV_X1 U1034 ( .A(KEYINPUT55), .ZN(n1037) );
  XOR2_X1 U1035 ( .A(G34), .B(KEYINPUT120), .Z(n934) );
  XNOR2_X1 U1036 ( .A(G2084), .B(KEYINPUT54), .ZN(n933) );
  XNOR2_X1 U1037 ( .A(n934), .B(n933), .ZN(n952) );
  XNOR2_X1 U1038 ( .A(G2090), .B(G35), .ZN(n950) );
  XOR2_X1 U1039 ( .A(G2072), .B(G33), .Z(n935) );
  NAND2_X1 U1040 ( .A1(n935), .A2(G28), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(n936), .B(G32), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(G27), .B(KEYINPUT118), .ZN(n938) );
  XNOR2_X1 U1043 ( .A(n938), .B(n937), .ZN(n939) );
  NAND2_X1 U1044 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1045 ( .A(n941), .B(KEYINPUT119), .ZN(n945) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n943) );
  XNOR2_X1 U1047 ( .A(G1991), .B(G25), .ZN(n942) );
  NOR2_X1 U1048 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1049 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1050 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1051 ( .A(KEYINPUT53), .B(n948), .ZN(n949) );
  NOR2_X1 U1052 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1054 ( .A(n1037), .B(n953), .ZN(n955) );
  INV_X1 U1055 ( .A(G29), .ZN(n954) );
  NAND2_X1 U1056 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n956), .ZN(n1012) );
  INV_X1 U1058 ( .A(G16), .ZN(n1008) );
  XNOR2_X1 U1059 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n957) );
  XNOR2_X1 U1060 ( .A(n1008), .B(n957), .ZN(n982) );
  XNOR2_X1 U1061 ( .A(G1966), .B(G168), .ZN(n959) );
  NAND2_X1 U1062 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1063 ( .A(n960), .B(KEYINPUT57), .ZN(n980) );
  XNOR2_X1 U1064 ( .A(G301), .B(G1961), .ZN(n963) );
  XNOR2_X1 U1065 ( .A(n961), .B(G1348), .ZN(n962) );
  NOR2_X1 U1066 ( .A1(n963), .A2(n962), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n964), .B(G1956), .ZN(n965) );
  XNOR2_X1 U1068 ( .A(n965), .B(KEYINPUT122), .ZN(n967) );
  NAND2_X1 U1069 ( .A1(n967), .A2(n966), .ZN(n969) );
  AND2_X1 U1070 ( .A1(G303), .A2(G1971), .ZN(n968) );
  NOR2_X1 U1071 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1072 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1073 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1074 ( .A1(n975), .A2(n974), .ZN(n978) );
  XNOR2_X1 U1075 ( .A(G1341), .B(n976), .ZN(n977) );
  NOR2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n1010) );
  XNOR2_X1 U1079 ( .A(KEYINPUT125), .B(G1966), .ZN(n983) );
  XNOR2_X1 U1080 ( .A(n983), .B(G21), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(G1961), .B(G5), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(G1986), .B(G24), .ZN(n985) );
  XNOR2_X1 U1083 ( .A(G1971), .B(G22), .ZN(n984) );
  NOR2_X1 U1084 ( .A1(n985), .A2(n984), .ZN(n987) );
  XOR2_X1 U1085 ( .A(G1976), .B(G23), .Z(n986) );
  NAND2_X1 U1086 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1087 ( .A(KEYINPUT58), .B(n988), .ZN(n989) );
  NOR2_X1 U1088 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1089 ( .A1(n992), .A2(n991), .ZN(n1005) );
  XOR2_X1 U1090 ( .A(G1981), .B(G6), .Z(n993) );
  XNOR2_X1 U1091 ( .A(KEYINPUT123), .B(n993), .ZN(n995) );
  XNOR2_X1 U1092 ( .A(G19), .B(G1341), .ZN(n994) );
  NOR2_X1 U1093 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1094 ( .A(KEYINPUT124), .B(n996), .ZN(n999) );
  XNOR2_X1 U1095 ( .A(n997), .B(G20), .ZN(n998) );
  NAND2_X1 U1096 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XOR2_X1 U1097 ( .A(KEYINPUT59), .B(G1348), .Z(n1000) );
  XNOR2_X1 U1098 ( .A(G4), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1099 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1100 ( .A(KEYINPUT60), .B(n1003), .Z(n1004) );
  NOR2_X1 U1101 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1103 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1104 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1105 ( .A1(n1012), .A2(n1011), .ZN(n1041) );
  XNOR2_X1 U1106 ( .A(G160), .B(G2084), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1035) );
  XNOR2_X1 U1111 ( .A(G2072), .B(n1021), .ZN(n1024) );
  XNOR2_X1 U1112 ( .A(G164), .B(G2078), .ZN(n1022) );
  XNOR2_X1 U1113 ( .A(n1022), .B(KEYINPUT116), .ZN(n1023) );
  NAND2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1115 ( .A(n1025), .B(KEYINPUT50), .ZN(n1026) );
  XOR2_X1 U1116 ( .A(KEYINPUT117), .B(n1026), .Z(n1031) );
  XOR2_X1 U1117 ( .A(G2090), .B(G162), .Z(n1027) );
  NOR2_X1 U1118 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1119 ( .A(KEYINPUT51), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1033) );
  NAND2_X1 U1121 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1123 ( .A(KEYINPUT52), .B(n1036), .ZN(n1038) );
  NAND2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1125 ( .A1(n1039), .A2(G29), .ZN(n1040) );
  NAND2_X1 U1126 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1127 ( .A(n1043), .B(n1042), .ZN(G311) );
  XNOR2_X1 U1128 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

