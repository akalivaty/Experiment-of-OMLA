

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(G2104), .ZN(n522) );
  NOR2_X2 U553 ( .A1(n603), .A2(n898), .ZN(n613) );
  AND2_X1 U554 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n587) );
  INV_X1 U556 ( .A(KEYINPUT91), .ZN(n631) );
  NOR2_X1 U557 ( .A1(n652), .A2(n651), .ZN(n653) );
  AND2_X2 U558 ( .A1(n705), .A2(n588), .ZN(n639) );
  NAND2_X1 U559 ( .A1(n677), .A2(n676), .ZN(n696) );
  XNOR2_X1 U560 ( .A(n669), .B(KEYINPUT32), .ZN(n677) );
  INV_X1 U561 ( .A(n520), .ZN(n982) );
  NOR2_X1 U562 ( .A1(n738), .A2(n518), .ZN(n739) );
  NOR2_X1 U563 ( .A1(n567), .A2(G651), .ZN(n784) );
  AND2_X1 U564 ( .A1(n704), .A2(n703), .ZN(n515) );
  AND2_X1 U565 ( .A1(n693), .A2(n692), .ZN(n516) );
  XNOR2_X1 U566 ( .A(n635), .B(n634), .ZN(n517) );
  AND2_X1 U567 ( .A1(n908), .A2(n752), .ZN(n518) );
  XNOR2_X1 U568 ( .A(KEYINPUT30), .B(KEYINPUT92), .ZN(n648) );
  XNOR2_X1 U569 ( .A(n649), .B(n648), .ZN(n650) );
  AND2_X1 U570 ( .A1(n646), .A2(n701), .ZN(n673) );
  INV_X1 U571 ( .A(n639), .ZN(n659) );
  AND2_X1 U572 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U573 ( .A(n589), .B(KEYINPUT87), .ZN(n701) );
  XNOR2_X1 U574 ( .A(KEYINPUT17), .B(n519), .ZN(n520) );
  NOR2_X1 U575 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U576 ( .A1(n567), .A2(n542), .ZN(n788) );
  NOR2_X2 U577 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  INV_X1 U578 ( .A(n520), .ZN(n530) );
  NAND2_X1 U579 ( .A1(G138), .A2(n530), .ZN(n521) );
  XNOR2_X1 U580 ( .A(n521), .B(KEYINPUT81), .ZN(n526) );
  BUF_X1 U581 ( .A(G2105), .Z(n527) );
  NOR2_X4 U582 ( .A1(n527), .A2(n522), .ZN(n984) );
  NAND2_X1 U583 ( .A1(G102), .A2(n984), .ZN(n524) );
  AND2_X2 U584 ( .A1(n522), .A2(n527), .ZN(n992) );
  NAND2_X1 U585 ( .A1(G126), .A2(n992), .ZN(n523) );
  NAND2_X1 U586 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U587 ( .A1(n526), .A2(n525), .ZN(n529) );
  AND2_X1 U588 ( .A1(G2104), .A2(n527), .ZN(n989) );
  NAND2_X1 U589 ( .A1(n989), .A2(G114), .ZN(n528) );
  AND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(G164) );
  NAND2_X1 U591 ( .A1(n982), .A2(G137), .ZN(n533) );
  NAND2_X1 U592 ( .A1(G101), .A2(n984), .ZN(n531) );
  XOR2_X1 U593 ( .A(KEYINPUT23), .B(n531), .Z(n532) );
  NAND2_X1 U594 ( .A1(n533), .A2(n532), .ZN(n537) );
  NAND2_X1 U595 ( .A1(G113), .A2(n989), .ZN(n535) );
  NAND2_X1 U596 ( .A1(G125), .A2(n992), .ZN(n534) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U598 ( .A1(n537), .A2(n536), .ZN(G160) );
  INV_X1 U599 ( .A(G651), .ZN(n542) );
  NOR2_X1 U600 ( .A1(G543), .A2(n542), .ZN(n539) );
  XNOR2_X1 U601 ( .A(KEYINPUT1), .B(KEYINPUT65), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(n783) );
  NAND2_X1 U603 ( .A1(G64), .A2(n783), .ZN(n541) );
  XOR2_X1 U604 ( .A(KEYINPUT0), .B(G543), .Z(n567) );
  NAND2_X1 U605 ( .A1(G52), .A2(n784), .ZN(n540) );
  NAND2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n788), .A2(G77), .ZN(n543) );
  XNOR2_X1 U608 ( .A(KEYINPUT67), .B(n543), .ZN(n546) );
  NOR2_X1 U609 ( .A1(G543), .A2(G651), .ZN(n787) );
  NAND2_X1 U610 ( .A1(n787), .A2(G90), .ZN(n544) );
  XOR2_X1 U611 ( .A(KEYINPUT66), .B(n544), .Z(n545) );
  NOR2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(KEYINPUT9), .ZN(n548) );
  NOR2_X1 U614 ( .A1(n549), .A2(n548), .ZN(G171) );
  INV_X1 U615 ( .A(G171), .ZN(G301) );
  NAND2_X1 U616 ( .A1(n787), .A2(G89), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U618 ( .A1(G76), .A2(n788), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT5), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G63), .A2(n783), .ZN(n555) );
  NAND2_X1 U622 ( .A1(G51), .A2(n784), .ZN(n554) );
  NAND2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n556), .Z(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G88), .A2(n787), .ZN(n561) );
  NAND2_X1 U629 ( .A1(G75), .A2(n788), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U631 ( .A1(G62), .A2(n783), .ZN(n563) );
  NAND2_X1 U632 ( .A1(G50), .A2(n784), .ZN(n562) );
  NAND2_X1 U633 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U634 ( .A1(n565), .A2(n564), .ZN(G166) );
  INV_X1 U635 ( .A(G166), .ZN(G303) );
  NAND2_X1 U636 ( .A1(G49), .A2(n784), .ZN(n566) );
  XNOR2_X1 U637 ( .A(n566), .B(KEYINPUT74), .ZN(n572) );
  NAND2_X1 U638 ( .A1(G74), .A2(G651), .ZN(n569) );
  NAND2_X1 U639 ( .A1(G87), .A2(n567), .ZN(n568) );
  NAND2_X1 U640 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U641 ( .A1(n783), .A2(n570), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n572), .A2(n571), .ZN(G288) );
  NAND2_X1 U643 ( .A1(G86), .A2(n787), .ZN(n574) );
  NAND2_X1 U644 ( .A1(G61), .A2(n783), .ZN(n573) );
  NAND2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U646 ( .A1(G73), .A2(n788), .ZN(n575) );
  XNOR2_X1 U647 ( .A(n575), .B(KEYINPUT75), .ZN(n576) );
  XNOR2_X1 U648 ( .A(n576), .B(KEYINPUT2), .ZN(n577) );
  NOR2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U650 ( .A1(n784), .A2(G48), .ZN(n579) );
  NAND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(G305) );
  NAND2_X1 U652 ( .A1(G85), .A2(n787), .ZN(n582) );
  NAND2_X1 U653 ( .A1(G60), .A2(n783), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U655 ( .A1(G72), .A2(n788), .ZN(n584) );
  NAND2_X1 U656 ( .A1(G47), .A2(n784), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  OR2_X1 U658 ( .A1(n586), .A2(n585), .ZN(G290) );
  XNOR2_X1 U659 ( .A(n587), .B(KEYINPUT64), .ZN(n705) );
  NAND2_X1 U660 ( .A1(G160), .A2(G40), .ZN(n706) );
  INV_X1 U661 ( .A(n706), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n659), .A2(G8), .ZN(n589) );
  INV_X1 U663 ( .A(n701), .ZN(n698) );
  AND2_X2 U664 ( .A1(n639), .A2(G1996), .ZN(n590) );
  XOR2_X1 U665 ( .A(KEYINPUT26), .B(n590), .Z(n592) );
  NAND2_X1 U666 ( .A1(n659), .A2(G1341), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n603) );
  NAND2_X1 U668 ( .A1(n787), .A2(G81), .ZN(n593) );
  XNOR2_X1 U669 ( .A(n593), .B(KEYINPUT12), .ZN(n595) );
  NAND2_X1 U670 ( .A1(G68), .A2(n788), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U672 ( .A(KEYINPUT13), .B(n596), .ZN(n602) );
  NAND2_X1 U673 ( .A1(G56), .A2(n783), .ZN(n597) );
  XOR2_X1 U674 ( .A(KEYINPUT14), .B(n597), .Z(n600) );
  NAND2_X1 U675 ( .A1(G43), .A2(n784), .ZN(n598) );
  XNOR2_X1 U676 ( .A(KEYINPUT69), .B(n598), .ZN(n599) );
  NOR2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n898) );
  NAND2_X1 U679 ( .A1(G54), .A2(n784), .ZN(n610) );
  NAND2_X1 U680 ( .A1(G92), .A2(n787), .ZN(n605) );
  NAND2_X1 U681 ( .A1(G66), .A2(n783), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n788), .A2(G79), .ZN(n606) );
  XOR2_X1 U684 ( .A(KEYINPUT70), .B(n606), .Z(n607) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X2 U686 ( .A(n611), .B(KEYINPUT15), .ZN(n1015) );
  OR2_X1 U687 ( .A1(n613), .A2(n1015), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n612), .B(KEYINPUT90), .ZN(n619) );
  NAND2_X1 U689 ( .A1(n613), .A2(n1015), .ZN(n617) );
  NOR2_X1 U690 ( .A1(n639), .A2(G1348), .ZN(n615) );
  NOR2_X1 U691 ( .A1(G2067), .A2(n659), .ZN(n614) );
  NOR2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n630) );
  NAND2_X1 U695 ( .A1(G65), .A2(n783), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G53), .A2(n784), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G91), .A2(n787), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G78), .A2(n788), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n757) );
  NAND2_X1 U702 ( .A1(n639), .A2(G2072), .ZN(n626) );
  XNOR2_X1 U703 ( .A(n626), .B(KEYINPUT27), .ZN(n628) );
  INV_X1 U704 ( .A(G1956), .ZN(n924) );
  NOR2_X1 U705 ( .A1(n924), .A2(n639), .ZN(n627) );
  NOR2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n757), .A2(n633), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(n631), .ZN(n636) );
  OR2_X1 U710 ( .A1(n633), .A2(n757), .ZN(n635) );
  XOR2_X1 U711 ( .A(KEYINPUT28), .B(KEYINPUT89), .Z(n634) );
  NAND2_X1 U712 ( .A1(n636), .A2(n517), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n637), .B(KEYINPUT29), .ZN(n643) );
  NAND2_X1 U714 ( .A1(G1961), .A2(n659), .ZN(n641) );
  XOR2_X1 U715 ( .A(G2078), .B(KEYINPUT88), .Z(n638) );
  XNOR2_X1 U716 ( .A(KEYINPUT25), .B(n638), .ZN(n844) );
  NAND2_X1 U717 ( .A1(n639), .A2(n844), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n644) );
  NOR2_X1 U719 ( .A1(G301), .A2(n644), .ZN(n642) );
  NOR2_X1 U720 ( .A1(n643), .A2(n642), .ZN(n655) );
  NAND2_X1 U721 ( .A1(G301), .A2(n644), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n645), .B(KEYINPUT93), .ZN(n652) );
  INV_X1 U723 ( .A(G1966), .ZN(n646) );
  NOR2_X1 U724 ( .A1(G2084), .A2(n659), .ZN(n670) );
  NOR2_X1 U725 ( .A1(n673), .A2(n670), .ZN(n647) );
  NAND2_X1 U726 ( .A1(G8), .A2(n647), .ZN(n649) );
  NOR2_X1 U727 ( .A1(n650), .A2(G168), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n653), .B(KEYINPUT31), .ZN(n654) );
  NOR2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n657) );
  INV_X1 U730 ( .A(KEYINPUT94), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n657), .B(n656), .ZN(n671) );
  AND2_X1 U732 ( .A1(G286), .A2(G8), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n671), .A2(n658), .ZN(n668) );
  INV_X1 U734 ( .A(G8), .ZN(n666) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XOR2_X1 U736 ( .A(KEYINPUT95), .B(n660), .Z(n662) );
  NOR2_X1 U737 ( .A1(G1971), .A2(n698), .ZN(n661) );
  NOR2_X1 U738 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(KEYINPUT96), .ZN(n664) );
  NAND2_X1 U740 ( .A1(n664), .A2(G303), .ZN(n665) );
  OR2_X1 U741 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U742 ( .A1(G8), .A2(n670), .ZN(n675) );
  INV_X1 U743 ( .A(n671), .ZN(n672) );
  NOR2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U745 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n681) );
  NOR2_X1 U747 ( .A1(G1971), .A2(G303), .ZN(n678) );
  NOR2_X1 U748 ( .A1(n681), .A2(n678), .ZN(n906) );
  NAND2_X1 U749 ( .A1(n696), .A2(n906), .ZN(n679) );
  XNOR2_X1 U750 ( .A(n679), .B(KEYINPUT97), .ZN(n680) );
  NOR2_X1 U751 ( .A1(n698), .A2(n680), .ZN(n687) );
  NAND2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n902) );
  INV_X1 U753 ( .A(KEYINPUT33), .ZN(n689) );
  NAND2_X1 U754 ( .A1(n701), .A2(n681), .ZN(n682) );
  NOR2_X1 U755 ( .A1(n689), .A2(n682), .ZN(n683) );
  XOR2_X1 U756 ( .A(n683), .B(KEYINPUT98), .Z(n688) );
  AND2_X1 U757 ( .A1(n902), .A2(n688), .ZN(n685) );
  XNOR2_X1 U758 ( .A(G1981), .B(G305), .ZN(n896) );
  INV_X1 U759 ( .A(n896), .ZN(n684) );
  AND2_X1 U760 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U761 ( .A1(n687), .A2(n686), .ZN(n693) );
  INV_X1 U762 ( .A(n688), .ZN(n690) );
  OR2_X1 U763 ( .A1(n690), .A2(n689), .ZN(n691) );
  OR2_X1 U764 ( .A1(n896), .A2(n691), .ZN(n692) );
  NOR2_X1 U765 ( .A1(G2090), .A2(G303), .ZN(n694) );
  NAND2_X1 U766 ( .A1(G8), .A2(n694), .ZN(n695) );
  XNOR2_X1 U767 ( .A(KEYINPUT99), .B(n697), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n704) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n700) );
  XNOR2_X1 U770 ( .A(KEYINPUT24), .B(n700), .ZN(n702) );
  NAND2_X1 U771 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U772 ( .A1(n516), .A2(n515), .ZN(n740) );
  NOR2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n752) );
  XNOR2_X1 U774 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n719) );
  NAND2_X1 U775 ( .A1(n984), .A2(G104), .ZN(n707) );
  XNOR2_X1 U776 ( .A(n707), .B(KEYINPUT82), .ZN(n709) );
  NAND2_X1 U777 ( .A1(G140), .A2(n982), .ZN(n708) );
  NAND2_X1 U778 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U779 ( .A(KEYINPUT34), .B(n710), .ZN(n716) );
  NAND2_X1 U780 ( .A1(n989), .A2(G116), .ZN(n711) );
  XOR2_X1 U781 ( .A(KEYINPUT83), .B(n711), .Z(n713) );
  NAND2_X1 U782 ( .A1(n992), .A2(G128), .ZN(n712) );
  NAND2_X1 U783 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U784 ( .A(n714), .B(KEYINPUT35), .Z(n715) );
  NOR2_X1 U785 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U786 ( .A(KEYINPUT36), .B(n717), .Z(n718) );
  XNOR2_X1 U787 ( .A(n719), .B(n718), .ZN(n999) );
  XNOR2_X1 U788 ( .A(G2067), .B(KEYINPUT37), .ZN(n749) );
  NOR2_X1 U789 ( .A1(n999), .A2(n749), .ZN(n874) );
  NAND2_X1 U790 ( .A1(n752), .A2(n874), .ZN(n747) );
  NAND2_X1 U791 ( .A1(G95), .A2(n984), .ZN(n721) );
  NAND2_X1 U792 ( .A1(G131), .A2(n982), .ZN(n720) );
  NAND2_X1 U793 ( .A1(n721), .A2(n720), .ZN(n725) );
  NAND2_X1 U794 ( .A1(G107), .A2(n989), .ZN(n723) );
  NAND2_X1 U795 ( .A1(G119), .A2(n992), .ZN(n722) );
  NAND2_X1 U796 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U797 ( .A1(n725), .A2(n724), .ZN(n1002) );
  INV_X1 U798 ( .A(G1991), .ZN(n837) );
  NOR2_X1 U799 ( .A1(n1002), .A2(n837), .ZN(n735) );
  NAND2_X1 U800 ( .A1(G117), .A2(n989), .ZN(n727) );
  NAND2_X1 U801 ( .A1(G129), .A2(n992), .ZN(n726) );
  NAND2_X1 U802 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U803 ( .A1(n984), .A2(G105), .ZN(n728) );
  XOR2_X1 U804 ( .A(KEYINPUT38), .B(n728), .Z(n729) );
  NOR2_X1 U805 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U806 ( .A(n731), .B(KEYINPUT86), .ZN(n733) );
  NAND2_X1 U807 ( .A1(G141), .A2(n982), .ZN(n732) );
  NAND2_X1 U808 ( .A1(n733), .A2(n732), .ZN(n998) );
  AND2_X1 U809 ( .A1(G1996), .A2(n998), .ZN(n734) );
  NOR2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n876) );
  INV_X1 U811 ( .A(n752), .ZN(n736) );
  NOR2_X1 U812 ( .A1(n876), .A2(n736), .ZN(n744) );
  INV_X1 U813 ( .A(n744), .ZN(n737) );
  NAND2_X1 U814 ( .A1(n747), .A2(n737), .ZN(n738) );
  XNOR2_X1 U815 ( .A(G1986), .B(G290), .ZN(n908) );
  NAND2_X1 U816 ( .A1(n740), .A2(n739), .ZN(n755) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n998), .ZN(n881) );
  AND2_X1 U818 ( .A1(n837), .A2(n1002), .ZN(n870) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n741) );
  NOR2_X1 U820 ( .A1(n870), .A2(n741), .ZN(n742) );
  XNOR2_X1 U821 ( .A(n742), .B(KEYINPUT100), .ZN(n743) );
  NOR2_X1 U822 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U823 ( .A1(n881), .A2(n745), .ZN(n746) );
  XNOR2_X1 U824 ( .A(n746), .B(KEYINPUT39), .ZN(n748) );
  NAND2_X1 U825 ( .A1(n748), .A2(n747), .ZN(n750) );
  NAND2_X1 U826 ( .A1(n999), .A2(n749), .ZN(n878) );
  NAND2_X1 U827 ( .A1(n750), .A2(n878), .ZN(n751) );
  XOR2_X1 U828 ( .A(KEYINPUT101), .B(n751), .Z(n753) );
  NAND2_X1 U829 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U830 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U831 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U832 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U833 ( .A(G120), .ZN(G236) );
  INV_X1 U834 ( .A(G82), .ZN(G220) );
  INV_X1 U835 ( .A(n757), .ZN(G299) );
  NAND2_X1 U836 ( .A1(G7), .A2(G661), .ZN(n758) );
  XNOR2_X1 U837 ( .A(n758), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U838 ( .A(G223), .ZN(n823) );
  NAND2_X1 U839 ( .A1(n823), .A2(G567), .ZN(n759) );
  XOR2_X1 U840 ( .A(KEYINPUT11), .B(n759), .Z(G234) );
  INV_X1 U841 ( .A(G860), .ZN(n765) );
  OR2_X1 U842 ( .A1(n898), .A2(n765), .ZN(G153) );
  NAND2_X1 U843 ( .A1(G868), .A2(G301), .ZN(n761) );
  OR2_X1 U844 ( .A1(n1015), .A2(G868), .ZN(n760) );
  NAND2_X1 U845 ( .A1(n761), .A2(n760), .ZN(G284) );
  INV_X1 U846 ( .A(G868), .ZN(n762) );
  NOR2_X1 U847 ( .A1(G286), .A2(n762), .ZN(n764) );
  NOR2_X1 U848 ( .A1(G868), .A2(G299), .ZN(n763) );
  NOR2_X1 U849 ( .A1(n764), .A2(n763), .ZN(G297) );
  NAND2_X1 U850 ( .A1(n765), .A2(G559), .ZN(n766) );
  NAND2_X1 U851 ( .A1(n766), .A2(n1015), .ZN(n767) );
  XNOR2_X1 U852 ( .A(n767), .B(KEYINPUT71), .ZN(n768) );
  XOR2_X1 U853 ( .A(KEYINPUT16), .B(n768), .Z(G148) );
  NAND2_X1 U854 ( .A1(n1015), .A2(G868), .ZN(n769) );
  NOR2_X1 U855 ( .A1(G559), .A2(n769), .ZN(n770) );
  XNOR2_X1 U856 ( .A(n770), .B(KEYINPUT72), .ZN(n772) );
  NOR2_X1 U857 ( .A1(n898), .A2(G868), .ZN(n771) );
  NOR2_X1 U858 ( .A1(n772), .A2(n771), .ZN(G282) );
  NAND2_X1 U859 ( .A1(G123), .A2(n992), .ZN(n773) );
  XNOR2_X1 U860 ( .A(n773), .B(KEYINPUT18), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n989), .A2(G111), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n779) );
  NAND2_X1 U863 ( .A1(G99), .A2(n984), .ZN(n777) );
  NAND2_X1 U864 ( .A1(G135), .A2(n982), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n1005) );
  XNOR2_X1 U867 ( .A(n1005), .B(G2096), .ZN(n781) );
  INV_X1 U868 ( .A(G2100), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(G156) );
  NAND2_X1 U870 ( .A1(n1015), .A2(G559), .ZN(n804) );
  XNOR2_X1 U871 ( .A(n898), .B(n804), .ZN(n782) );
  NOR2_X1 U872 ( .A1(n782), .A2(G860), .ZN(n794) );
  NAND2_X1 U873 ( .A1(G67), .A2(n783), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G55), .A2(n784), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n793) );
  NAND2_X1 U876 ( .A1(G93), .A2(n787), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G80), .A2(n788), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U879 ( .A(KEYINPUT73), .B(n791), .Z(n792) );
  NOR2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n798) );
  XNOR2_X1 U881 ( .A(n794), .B(n798), .ZN(G145) );
  NOR2_X1 U882 ( .A1(G868), .A2(n798), .ZN(n795) );
  XNOR2_X1 U883 ( .A(n795), .B(KEYINPUT77), .ZN(n807) );
  XNOR2_X1 U884 ( .A(G166), .B(KEYINPUT19), .ZN(n796) );
  XNOR2_X1 U885 ( .A(n796), .B(KEYINPUT76), .ZN(n797) );
  XNOR2_X1 U886 ( .A(n798), .B(n797), .ZN(n801) );
  XOR2_X1 U887 ( .A(G290), .B(G305), .Z(n799) );
  XNOR2_X1 U888 ( .A(n898), .B(n799), .ZN(n800) );
  XNOR2_X1 U889 ( .A(n801), .B(n800), .ZN(n802) );
  XNOR2_X1 U890 ( .A(n802), .B(G299), .ZN(n803) );
  XNOR2_X1 U891 ( .A(n803), .B(G288), .ZN(n1014) );
  XNOR2_X1 U892 ( .A(n1014), .B(n804), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G868), .A2(n805), .ZN(n806) );
  NAND2_X1 U894 ( .A1(n807), .A2(n806), .ZN(G295) );
  NAND2_X1 U895 ( .A1(G2078), .A2(G2084), .ZN(n809) );
  XOR2_X1 U896 ( .A(KEYINPUT20), .B(KEYINPUT78), .Z(n808) );
  XNOR2_X1 U897 ( .A(n809), .B(n808), .ZN(n810) );
  NAND2_X1 U898 ( .A1(G2090), .A2(n810), .ZN(n811) );
  XNOR2_X1 U899 ( .A(KEYINPUT21), .B(n811), .ZN(n812) );
  NAND2_X1 U900 ( .A1(n812), .A2(G2072), .ZN(G158) );
  XOR2_X1 U901 ( .A(KEYINPUT68), .B(G132), .Z(G219) );
  XNOR2_X1 U902 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U903 ( .A1(G661), .A2(G483), .ZN(n821) );
  NOR2_X1 U904 ( .A1(G219), .A2(G220), .ZN(n814) );
  XNOR2_X1 U905 ( .A(KEYINPUT79), .B(KEYINPUT22), .ZN(n813) );
  XNOR2_X1 U906 ( .A(n814), .B(n813), .ZN(n815) );
  NOR2_X1 U907 ( .A1(n815), .A2(G218), .ZN(n816) );
  NAND2_X1 U908 ( .A1(G96), .A2(n816), .ZN(n952) );
  NAND2_X1 U909 ( .A1(n952), .A2(G2106), .ZN(n820) );
  NAND2_X1 U910 ( .A1(G69), .A2(G108), .ZN(n817) );
  NOR2_X1 U911 ( .A1(G236), .A2(n817), .ZN(n818) );
  NAND2_X1 U912 ( .A1(G57), .A2(n818), .ZN(n953) );
  NAND2_X1 U913 ( .A1(n953), .A2(G567), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n1024) );
  NOR2_X1 U915 ( .A1(n821), .A2(n1024), .ZN(n822) );
  XNOR2_X1 U916 ( .A(n822), .B(KEYINPUT80), .ZN(n827) );
  NAND2_X1 U917 ( .A1(G36), .A2(n827), .ZN(G176) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n823), .ZN(G217) );
  NAND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n824) );
  XOR2_X1 U920 ( .A(KEYINPUT104), .B(n824), .Z(n825) );
  NAND2_X1 U921 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(G188) );
  XNOR2_X1 U924 ( .A(G69), .B(KEYINPUT105), .ZN(G235) );
  XOR2_X1 U925 ( .A(G108), .B(KEYINPUT112), .Z(G238) );
  NAND2_X1 U927 ( .A1(G124), .A2(n992), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n828), .B(KEYINPUT44), .ZN(n830) );
  NAND2_X1 U929 ( .A1(n989), .A2(G112), .ZN(n829) );
  NAND2_X1 U930 ( .A1(n830), .A2(n829), .ZN(n834) );
  NAND2_X1 U931 ( .A1(G100), .A2(n984), .ZN(n832) );
  NAND2_X1 U932 ( .A1(G136), .A2(n982), .ZN(n831) );
  NAND2_X1 U933 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U934 ( .A1(n834), .A2(n833), .ZN(G162) );
  XNOR2_X1 U935 ( .A(KEYINPUT54), .B(KEYINPUT118), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n835), .B(G34), .ZN(n836) );
  XNOR2_X1 U937 ( .A(G2084), .B(n836), .ZN(n855) );
  XNOR2_X1 U938 ( .A(G2090), .B(G35), .ZN(n852) );
  XNOR2_X1 U939 ( .A(n837), .B(G25), .ZN(n838) );
  NAND2_X1 U940 ( .A1(n838), .A2(G28), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n839), .B(KEYINPUT115), .ZN(n843) );
  XNOR2_X1 U942 ( .A(G2067), .B(G26), .ZN(n841) );
  XNOR2_X1 U943 ( .A(G33), .B(G2072), .ZN(n840) );
  NOR2_X1 U944 ( .A1(n841), .A2(n840), .ZN(n842) );
  NAND2_X1 U945 ( .A1(n843), .A2(n842), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n844), .B(G27), .ZN(n846) );
  XNOR2_X1 U947 ( .A(G32), .B(G1996), .ZN(n845) );
  NOR2_X1 U948 ( .A1(n846), .A2(n845), .ZN(n847) );
  XOR2_X1 U949 ( .A(KEYINPUT116), .B(n847), .Z(n848) );
  NOR2_X1 U950 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U951 ( .A(KEYINPUT53), .B(n850), .ZN(n851) );
  NOR2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U953 ( .A(KEYINPUT117), .B(n853), .ZN(n854) );
  NOR2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(KEYINPUT55), .B(n856), .Z(n857) );
  NOR2_X1 U956 ( .A1(G29), .A2(n857), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n858), .B(KEYINPUT119), .ZN(n893) );
  NAND2_X1 U958 ( .A1(G103), .A2(n984), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G139), .A2(n982), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n866) );
  NAND2_X1 U961 ( .A1(n989), .A2(G115), .ZN(n861) );
  XOR2_X1 U962 ( .A(KEYINPUT109), .B(n861), .Z(n863) );
  NAND2_X1 U963 ( .A1(n992), .A2(G127), .ZN(n862) );
  NAND2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U965 ( .A(KEYINPUT47), .B(n864), .Z(n865) );
  NOR2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n996) );
  XOR2_X1 U967 ( .A(G2072), .B(n996), .Z(n868) );
  XOR2_X1 U968 ( .A(G164), .B(G2078), .Z(n867) );
  NOR2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U970 ( .A(KEYINPUT50), .B(n869), .Z(n887) );
  XNOR2_X1 U971 ( .A(G160), .B(G2084), .ZN(n872) );
  NOR2_X1 U972 ( .A1(n870), .A2(n1005), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U976 ( .A(n877), .B(KEYINPUT113), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n884) );
  XOR2_X1 U978 ( .A(G2090), .B(G162), .Z(n880) );
  NOR2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U980 ( .A(n882), .B(KEYINPUT51), .ZN(n883) );
  NOR2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(KEYINPUT114), .B(n885), .Z(n886) );
  NOR2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U984 ( .A(n888), .B(KEYINPUT52), .ZN(n890) );
  INV_X1 U985 ( .A(KEYINPUT55), .ZN(n889) );
  NAND2_X1 U986 ( .A1(n890), .A2(n889), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G29), .A2(n891), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n949) );
  INV_X1 U989 ( .A(G16), .ZN(n944) );
  XOR2_X1 U990 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n894) );
  XNOR2_X1 U991 ( .A(n944), .B(n894), .ZN(n917) );
  XOR2_X1 U992 ( .A(G168), .B(G1966), .Z(n895) );
  NOR2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U994 ( .A(KEYINPUT57), .B(n897), .Z(n915) );
  XOR2_X1 U995 ( .A(G1348), .B(n1015), .Z(n900) );
  XNOR2_X1 U996 ( .A(n898), .B(G1341), .ZN(n899) );
  NOR2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n910) );
  NAND2_X1 U998 ( .A1(G1971), .A2(G303), .ZN(n901) );
  NAND2_X1 U999 ( .A1(n902), .A2(n901), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(G1956), .B(G299), .ZN(n903) );
  NOR2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(n905) );
  NAND2_X1 U1002 ( .A1(n906), .A2(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(n908), .A2(n907), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(n910), .A2(n909), .ZN(n913) );
  XOR2_X1 U1005 ( .A(G1961), .B(G301), .Z(n911) );
  XNOR2_X1 U1006 ( .A(KEYINPUT121), .B(n911), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1008 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1009 ( .A1(n917), .A2(n916), .ZN(n946) );
  XOR2_X1 U1010 ( .A(G1986), .B(G24), .Z(n921) );
  XNOR2_X1 U1011 ( .A(G1971), .B(G22), .ZN(n919) );
  XNOR2_X1 U1012 ( .A(G23), .B(G1976), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1014 ( .A1(n921), .A2(n920), .ZN(n923) );
  XNOR2_X1 U1015 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n922) );
  XNOR2_X1 U1016 ( .A(n923), .B(n922), .ZN(n938) );
  XNOR2_X1 U1017 ( .A(G1966), .B(G21), .ZN(n936) );
  XNOR2_X1 U1018 ( .A(G20), .B(n924), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(G1341), .B(G19), .ZN(n926) );
  XNOR2_X1 U1020 ( .A(G1981), .B(G6), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n931) );
  XOR2_X1 U1023 ( .A(KEYINPUT59), .B(G1348), .Z(n929) );
  XNOR2_X1 U1024 ( .A(G4), .B(n929), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n934) );
  XNOR2_X1 U1026 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n932) );
  XNOR2_X1 U1027 ( .A(n932), .B(KEYINPUT60), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(n934), .B(n933), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n941) );
  XNOR2_X1 U1031 ( .A(KEYINPUT122), .B(G1961), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(G5), .B(n939), .ZN(n940) );
  NOR2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(KEYINPUT61), .B(n942), .ZN(n943) );
  NAND2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1036 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1037 ( .A(n947), .B(KEYINPUT126), .ZN(n948) );
  NOR2_X1 U1038 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1039 ( .A1(n950), .A2(G11), .ZN(n951) );
  XOR2_X1 U1040 ( .A(KEYINPUT62), .B(n951), .Z(G311) );
  XNOR2_X1 U1041 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1042 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1043 ( .A1(n953), .A2(n952), .ZN(G325) );
  INV_X1 U1044 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1045 ( .A(G2443), .B(G1341), .ZN(n962) );
  XNOR2_X1 U1046 ( .A(G2430), .B(G2446), .ZN(n960) );
  XOR2_X1 U1047 ( .A(G2454), .B(G2451), .Z(n955) );
  XNOR2_X1 U1048 ( .A(G2427), .B(G2435), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(n955), .B(n954), .ZN(n956) );
  XOR2_X1 U1050 ( .A(n956), .B(G2438), .Z(n958) );
  XNOR2_X1 U1051 ( .A(G1348), .B(KEYINPUT102), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(n958), .B(n957), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(n960), .B(n959), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n962), .B(n961), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n963), .A2(G14), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(KEYINPUT103), .B(n964), .ZN(G401) );
  XOR2_X1 U1057 ( .A(G2100), .B(G2096), .Z(n966) );
  XNOR2_X1 U1058 ( .A(G2067), .B(G2090), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(n966), .B(n965), .ZN(n970) );
  XOR2_X1 U1060 ( .A(G2678), .B(KEYINPUT42), .Z(n968) );
  XNOR2_X1 U1061 ( .A(G2072), .B(KEYINPUT43), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n968), .B(n967), .ZN(n969) );
  XOR2_X1 U1063 ( .A(n970), .B(n969), .Z(n972) );
  XNOR2_X1 U1064 ( .A(G2078), .B(G2084), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(n972), .B(n971), .ZN(G227) );
  XOR2_X1 U1066 ( .A(G1981), .B(G1971), .Z(n974) );
  XNOR2_X1 U1067 ( .A(G1996), .B(G1961), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(n974), .B(n973), .ZN(n975) );
  XOR2_X1 U1069 ( .A(n975), .B(KEYINPUT41), .Z(n977) );
  XNOR2_X1 U1070 ( .A(G1966), .B(G1976), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(n977), .B(n976), .ZN(n981) );
  XOR2_X1 U1072 ( .A(G2474), .B(G1956), .Z(n979) );
  XNOR2_X1 U1073 ( .A(G1991), .B(G1986), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(n979), .B(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n981), .B(n980), .ZN(G229) );
  NAND2_X1 U1076 ( .A1(n982), .A2(G142), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT108), .B(n983), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n984), .A2(G106), .ZN(n985) );
  XOR2_X1 U1079 ( .A(KEYINPUT107), .B(n985), .Z(n986) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(n988), .B(KEYINPUT45), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(G118), .A2(n989), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n992), .A2(G130), .ZN(n993) );
  XOR2_X1 U1085 ( .A(KEYINPUT106), .B(n993), .Z(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n997) );
  XOR2_X1 U1087 ( .A(n997), .B(n996), .Z(n1001) );
  XOR2_X1 U1088 ( .A(n999), .B(n998), .Z(n1000) );
  XNOR2_X1 U1089 ( .A(n1001), .B(n1000), .ZN(n1011) );
  XOR2_X1 U1090 ( .A(KEYINPUT48), .B(KEYINPUT110), .Z(n1004) );
  XNOR2_X1 U1091 ( .A(n1002), .B(KEYINPUT46), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1004), .B(n1003), .ZN(n1006) );
  XOR2_X1 U1093 ( .A(n1006), .B(n1005), .Z(n1008) );
  XNOR2_X1 U1094 ( .A(G160), .B(G162), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1008), .B(n1007), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(G164), .B(n1009), .Z(n1010) );
  XNOR2_X1 U1097 ( .A(n1011), .B(n1010), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(G37), .A2(n1012), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(KEYINPUT111), .B(n1013), .Z(G395) );
  XOR2_X1 U1100 ( .A(n1014), .B(G286), .Z(n1017) );
  XNOR2_X1 U1101 ( .A(G171), .B(n1015), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(n1017), .B(n1016), .ZN(n1018) );
  NOR2_X1 U1103 ( .A1(G37), .A2(n1018), .ZN(G397) );
  OR2_X1 U1104 ( .A1(n1024), .A2(G401), .ZN(n1021) );
  NOR2_X1 U1105 ( .A1(G227), .A2(G229), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(KEYINPUT49), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(G395), .A2(G397), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(G225) );
  INV_X1 U1110 ( .A(G225), .ZN(G308) );
  INV_X1 U1111 ( .A(n1024), .ZN(G319) );
  INV_X1 U1112 ( .A(G57), .ZN(G237) );
endmodule

