//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974;
  INV_X1    g000(.A(KEYINPUT26), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  AOI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(KEYINPUT69), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT69), .B1(new_n203), .B2(KEYINPUT70), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n204), .A2(new_n206), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT28), .ZN(new_n219));
  OR2_X1    g018(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n220));
  NAND2_X1  g019(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(G183gat), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT65), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G183gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n226), .A3(KEYINPUT27), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n219), .A2(new_n222), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n218), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n223), .A2(KEYINPUT27), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT27), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G183gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n229), .A2(new_n230), .A3(new_n232), .A4(new_n216), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n233), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n228), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT23), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n203), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n237), .A2(new_n238), .B1(new_n211), .B2(new_n212), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT25), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n229), .A2(new_n224), .A3(new_n226), .A4(new_n216), .ZN(new_n241));
  NAND2_X1  g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT24), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT24), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(G183gat), .A3(G190gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n241), .A2(KEYINPUT67), .A3(new_n246), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n240), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n246), .B1(G183gat), .B2(G190gat), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT25), .B1(new_n252), .B2(new_n239), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n235), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(G226gat), .A2(G233gat), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT29), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n255), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G197gat), .B(G204gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT22), .ZN(new_n261));
  INV_X1    g060(.A(G211gat), .ZN(new_n262));
  INV_X1    g061(.A(G218gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n259), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G8gat), .B(G36gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(G64gat), .B(G92gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  OAI21_X1  g071(.A(new_n267), .B1(new_n256), .B2(new_n258), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n274), .B(KEYINPUT30), .Z(new_n275));
  NAND2_X1  g074(.A1(new_n269), .A2(new_n273), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n272), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n269), .A2(KEYINPUT75), .A3(new_n273), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n239), .A2(KEYINPUT25), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n241), .A2(new_n246), .A3(KEYINPUT67), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT67), .B1(new_n241), .B2(new_n246), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n253), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n233), .A2(KEYINPUT28), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n228), .A2(new_n288), .A3(new_n242), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n286), .A2(new_n287), .B1(new_n289), .B2(new_n215), .ZN(new_n290));
  INV_X1    g089(.A(G127gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G134gat), .ZN(new_n292));
  INV_X1    g091(.A(G134gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G127gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n297));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G113gat), .B(G120gat), .Z(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT72), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n302), .A2(new_n293), .A3(G127gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(G127gat), .B(G134gat), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n303), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n295), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n299), .A2(new_n301), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT74), .B1(new_n290), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n299), .A2(new_n301), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n305), .A2(new_n306), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n254), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(new_n254), .B2(new_n312), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n290), .A2(KEYINPUT73), .A3(new_n307), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G227gat), .A2(G233gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT34), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n308), .A2(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT34), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n320), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT33), .B1(new_n319), .B2(new_n321), .ZN(new_n326));
  XOR2_X1   g125(.A(G15gat), .B(G43gat), .Z(new_n327));
  XNOR2_X1  g126(.A(G71gat), .B(G99gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n322), .B(new_n325), .C1(new_n326), .C2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT33), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(new_n323), .B2(new_n320), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n324), .B1(new_n323), .B2(new_n320), .ZN(new_n334));
  AND4_X1   g133(.A1(new_n324), .A2(new_n314), .A3(new_n318), .A4(new_n320), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n333), .B(new_n329), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT32), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n331), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n339), .B1(new_n331), .B2(new_n336), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT88), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n331), .A2(new_n336), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n338), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n331), .A2(new_n336), .A3(new_n339), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT88), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n282), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(G148gat), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n352));
  INV_X1    g151(.A(G148gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(G141gat), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT78), .ZN(new_n358));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT79), .B1(new_n359), .B2(KEYINPUT2), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(KEYINPUT79), .A3(KEYINPUT2), .ZN(new_n362));
  OR2_X1    g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n361), .A2(new_n362), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n351), .A2(new_n356), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n358), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G155gat), .B(G162gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(G141gat), .A2(G148gat), .ZN(new_n369));
  INV_X1    g168(.A(G141gat), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT2), .B1(new_n370), .B2(new_n353), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n368), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT3), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT3), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n367), .A2(new_n376), .A3(new_n373), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n312), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT5), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n374), .A2(KEYINPUT80), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n384), .A3(new_n373), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n382), .A2(new_n383), .A3(new_n307), .A4(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n307), .A2(new_n367), .A3(new_n373), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT4), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n380), .A2(new_n381), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n351), .A2(new_n356), .A3(new_n365), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n365), .B1(new_n351), .B2(new_n356), .ZN(new_n393));
  INV_X1    g192(.A(new_n362), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n368), .B1(new_n394), .B2(new_n360), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n312), .B1(new_n396), .B2(new_n372), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n387), .ZN(new_n398));
  INV_X1    g197(.A(new_n379), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n391), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI211_X1 g199(.A(KEYINPUT81), .B(new_n379), .C1(new_n397), .C2(new_n387), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT5), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n307), .A4(new_n385), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n383), .ZN(new_n404));
  AND4_X1   g203(.A1(new_n403), .A2(new_n378), .A3(new_n379), .A4(new_n404), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n402), .A2(new_n405), .A3(KEYINPUT82), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n307), .A2(new_n367), .A3(new_n373), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n307), .B1(new_n373), .B2(new_n367), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n399), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT81), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n398), .A2(new_n391), .A3(new_n399), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n381), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n403), .A2(new_n378), .A3(new_n379), .A4(new_n404), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n407), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n390), .B1(new_n406), .B2(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(G1gat), .B(G29gat), .Z(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G57gat), .B(G85gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n424));
  INV_X1    g223(.A(new_n390), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT82), .B1(new_n402), .B2(new_n405), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n412), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n427), .A2(new_n407), .A3(KEYINPUT5), .A4(new_n414), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n425), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n421), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n426), .A2(new_n428), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n421), .B1(new_n433), .B2(new_n390), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n434), .B2(KEYINPUT6), .ZN(new_n435));
  NOR4_X1   g234(.A1(new_n429), .A2(KEYINPUT84), .A3(new_n424), .A4(new_n421), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(G22gat), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n376), .B1(new_n267), .B2(KEYINPUT29), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n374), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT85), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n377), .A2(new_n257), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n267), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(new_n446), .A3(new_n374), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(G228gat), .A3(G233gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(G228gat), .A2(G233gat), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n382), .A2(new_n385), .ZN(new_n451));
  INV_X1    g250(.A(new_n441), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n450), .B(new_n445), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT31), .B(G50gat), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n449), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n449), .B2(new_n453), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n440), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n449), .A2(new_n453), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n454), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n439), .A3(new_n456), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n437), .A2(new_n467), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n348), .A2(new_n468), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n340), .A2(new_n341), .A3(new_n463), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n437), .A2(new_n282), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT35), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n471), .B2(KEYINPUT35), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n437), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n275), .A2(new_n281), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n463), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n379), .B1(new_n389), .B2(new_n378), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT39), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n422), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT86), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT39), .B1(new_n398), .B2(new_n399), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n484), .B(KEYINPUT87), .Z(new_n485));
  OR2_X1    g284(.A1(new_n485), .A2(new_n479), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT40), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n483), .A2(KEYINPUT40), .A3(new_n486), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n477), .A2(new_n489), .A3(new_n423), .A4(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT38), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n278), .A2(KEYINPUT37), .A3(new_n280), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT37), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n269), .A2(new_n494), .A3(new_n273), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n495), .A2(new_n279), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n492), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n276), .A2(KEYINPUT37), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n498), .A2(new_n492), .A3(new_n279), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n274), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n501), .B(new_n431), .C1(new_n435), .C2(new_n436), .ZN(new_n502));
  INV_X1    g301(.A(new_n463), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n491), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n340), .A2(new_n341), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT36), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(new_n340), .B2(new_n341), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n478), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n475), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G113gat), .B(G141gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(G197gat), .ZN(new_n513));
  XOR2_X1   g312(.A(KEYINPUT11), .B(G169gat), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT12), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT15), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT91), .B(G29gat), .ZN(new_n519));
  INV_X1    g318(.A(G36gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(G29gat), .A2(G36gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT14), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n518), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT14), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n522), .B(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n526), .B(KEYINPUT15), .C1(new_n520), .C2(new_n519), .ZN(new_n527));
  XNOR2_X1  g326(.A(G43gat), .B(G50gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n521), .A2(new_n523), .ZN(new_n530));
  INV_X1    g329(.A(new_n528), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(KEYINPUT15), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT93), .ZN(new_n535));
  INV_X1    g334(.A(G1gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(KEYINPUT93), .A3(G1gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT16), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G8gat), .ZN(new_n542));
  INV_X1    g341(.A(G8gat), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n537), .A2(new_n543), .A3(new_n538), .A4(new_n540), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n533), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n547), .B(KEYINPUT13), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n547), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n533), .A2(new_n545), .ZN(new_n551));
  NAND2_X1  g350(.A1(KEYINPUT92), .A2(KEYINPUT17), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT92), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n533), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n529), .A2(new_n532), .A3(new_n553), .A4(new_n554), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n542), .A2(new_n559), .A3(new_n544), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n559), .B1(new_n542), .B2(new_n544), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI211_X1 g361(.A(new_n550), .B(new_n551), .C1(new_n558), .C2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n549), .B1(new_n563), .B2(KEYINPUT18), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n551), .B1(new_n558), .B2(new_n562), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n547), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT18), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n517), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n567), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n563), .A2(KEYINPUT18), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n570), .A2(new_n571), .A3(new_n516), .A4(new_n549), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n574));
  INV_X1    g373(.A(G64gat), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n575), .A2(G57gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(G57gat), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G71gat), .ZN(new_n579));
  INV_X1    g378(.A(G78gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT95), .ZN(new_n583));
  OAI22_X1  g382(.A1(new_n581), .A2(new_n582), .B1(new_n574), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n578), .B(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n545), .B1(KEYINPUT21), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT97), .ZN(new_n587));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT96), .ZN(new_n589));
  XOR2_X1   g388(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n587), .B(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n593));
  XOR2_X1   g392(.A(G127gat), .B(G155gat), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n592), .A2(new_n598), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n603));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT8), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT99), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT7), .ZN(new_n613));
  OAI211_X1 g412(.A(G85gat), .B(G92gat), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G99gat), .B(G106gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n611), .A2(new_n616), .A3(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n558), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n624), .A2(new_n533), .B1(KEYINPUT41), .B2(new_n602), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G190gat), .B(G218gat), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n606), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n632), .A2(new_n605), .A3(new_n628), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n601), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G230gat), .A2(G233gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n585), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n611), .A2(new_n618), .A3(new_n616), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n618), .B1(new_n611), .B2(new_n616), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n620), .A2(new_n585), .A3(new_n621), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT100), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n622), .A2(new_n643), .A3(new_n637), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT10), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n636), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(G120gat), .B(G148gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT101), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n642), .A2(new_n644), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n648), .B(new_n653), .C1(new_n636), .C2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n636), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n648), .A2(KEYINPUT102), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n658), .B(new_n636), .C1(new_n645), .C2(new_n647), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n656), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n655), .B1(new_n660), .B2(new_n653), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n635), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n511), .A2(new_n573), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n437), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n536), .ZN(G1324gat));
  NOR2_X1   g466(.A1(new_n665), .A2(new_n282), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n543), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n669), .B1(new_n673), .B2(KEYINPUT42), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(KEYINPUT42), .B2(new_n673), .ZN(G1325gat));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n509), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n506), .A2(KEYINPUT104), .A3(new_n508), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n665), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n343), .A2(new_n347), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n683), .A2(G15gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n681), .B1(new_n665), .B2(new_n684), .ZN(G1326gat));
  NOR2_X1   g484(.A1(new_n665), .A2(new_n503), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT43), .B(G22gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  INV_X1    g487(.A(new_n601), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n631), .A2(new_n633), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n689), .A2(new_n690), .A3(new_n661), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n511), .A2(new_n573), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n476), .A3(new_n519), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n511), .B2(new_n634), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n478), .A2(new_n677), .A3(new_n504), .A4(new_n678), .ZN(new_n700));
  AOI211_X1 g499(.A(new_n690), .B(new_n699), .C1(new_n475), .C2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n573), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n689), .A2(new_n704), .A3(new_n661), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n437), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n694), .B1(new_n707), .B2(new_n519), .ZN(G1328gat));
  NAND3_X1  g507(.A1(new_n511), .A2(new_n573), .A3(new_n691), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(G36gat), .A3(new_n282), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT46), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n706), .B2(new_n282), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G36gat), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n706), .A2(new_n712), .A3(new_n282), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(G1329gat));
  NOR3_X1   g515(.A1(new_n709), .A2(G43gat), .A3(new_n683), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n679), .B(new_n705), .C1(new_n696), .C2(new_n701), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(G43gat), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(KEYINPUT107), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(KEYINPUT47), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n719), .A2(KEYINPUT107), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(G1330gat));
  OAI211_X1 g523(.A(new_n463), .B(new_n705), .C1(new_n696), .C2(new_n701), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(G50gat), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n503), .A2(G50gat), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n692), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n709), .A2(KEYINPUT109), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(KEYINPUT108), .B(KEYINPUT48), .C1(new_n726), .C2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734));
  AOI22_X1  g533(.A1(G50gat), .A2(new_n725), .B1(new_n730), .B2(new_n731), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n733), .A2(new_n737), .ZN(G1331gat));
  NAND2_X1  g537(.A1(new_n475), .A2(new_n700), .ZN(new_n739));
  NOR4_X1   g538(.A1(new_n601), .A2(new_n662), .A3(new_n573), .A4(new_n634), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n476), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g543(.A1(new_n741), .A2(new_n282), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n745), .B2(new_n746), .ZN(G1333gat));
  OAI21_X1  g548(.A(G71gat), .B1(new_n741), .B2(new_n680), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n682), .A2(new_n579), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n741), .B2(new_n751), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g552(.A1(new_n741), .A2(new_n503), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(new_n580), .ZN(G1335gat));
  NOR3_X1   g554(.A1(new_n689), .A2(new_n573), .A3(new_n662), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n703), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757), .B2(new_n437), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n689), .A2(new_n573), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n348), .A2(new_n468), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n471), .A2(KEYINPUT35), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT90), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT35), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n760), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND4_X1   g563(.A1(new_n478), .A2(new_n677), .A3(new_n504), .A4(new_n678), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n634), .B(new_n759), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n739), .A2(KEYINPUT51), .A3(new_n634), .A4(new_n759), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n662), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n608), .A3(new_n476), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n758), .A2(new_n771), .ZN(G1336gat));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n768), .A2(new_n769), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n282), .A2(new_n662), .A3(G92gat), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT52), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n477), .B(new_n756), .C1(new_n696), .C2(new_n701), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G92gat), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n775), .B(KEYINPUT110), .Z(new_n781));
  NAND2_X1  g580(.A1(new_n774), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n773), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n776), .A2(new_n778), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n777), .A2(G92gat), .B1(new_n774), .B2(new_n781), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n785), .B(KEYINPUT111), .C1(new_n780), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(G1337gat));
  OAI21_X1  g587(.A(G99gat), .B1(new_n757), .B2(new_n680), .ZN(new_n789));
  INV_X1    g588(.A(new_n770), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n683), .A2(G99gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(G1338gat));
  NOR2_X1   g591(.A1(new_n503), .A2(G106gat), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n770), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n463), .B(new_n756), .C1(new_n696), .C2(new_n701), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n795), .A2(G106gat), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT53), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n798), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n799), .A2(G106gat), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n794), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n797), .B1(new_n801), .B2(new_n803), .ZN(G1339gat));
  NOR2_X1   g603(.A1(new_n565), .A2(new_n547), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n546), .A2(new_n548), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n515), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n572), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n661), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n657), .A2(new_n812), .A3(new_n659), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n654), .A2(new_n646), .ZN(new_n814));
  INV_X1    g613(.A(new_n636), .ZN(new_n815));
  INV_X1    g614(.A(new_n647), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(KEYINPUT54), .A3(new_n648), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n813), .A2(KEYINPUT55), .A3(new_n652), .A4(new_n818), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n819), .A2(new_n573), .A3(new_n655), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n657), .A2(new_n812), .A3(new_n659), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n652), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n634), .B1(new_n811), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n824), .A2(new_n634), .A3(new_n655), .A4(new_n819), .ZN(new_n827));
  INV_X1    g626(.A(new_n808), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n601), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n663), .A2(new_n573), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n463), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(new_n476), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n505), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n477), .ZN(new_n836));
  AOI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n573), .ZN(new_n837));
  INV_X1    g636(.A(new_n348), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT115), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n573), .A2(G113gat), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n837), .B1(new_n840), .B2(new_n841), .ZN(G1340gat));
  AOI21_X1  g641(.A(G120gat), .B1(new_n836), .B2(new_n661), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n661), .A2(G120gat), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n840), .B2(new_n844), .ZN(G1341gat));
  NAND3_X1  g644(.A1(new_n836), .A2(new_n291), .A3(new_n689), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n840), .A2(new_n689), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n291), .ZN(G1342gat));
  NAND2_X1  g647(.A1(new_n282), .A2(new_n634), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT116), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n835), .A2(G134gat), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT56), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n840), .A2(new_n634), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n293), .ZN(G1343gat));
  NAND2_X1  g653(.A1(new_n824), .A2(KEYINPUT117), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n856), .B(new_n821), .C1(new_n822), .C2(new_n823), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n820), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n634), .B1(new_n858), .B2(new_n809), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n601), .B1(new_n859), .B2(new_n829), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n832), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(KEYINPUT57), .A3(new_n463), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n503), .B1(new_n830), .B2(new_n832), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(KEYINPUT57), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n680), .A2(new_n476), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n477), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n573), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n349), .A2(new_n350), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n866), .A2(new_n863), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n573), .A2(new_n370), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT118), .Z(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT58), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n354), .A2(new_n355), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n870), .A2(new_n877), .A3(new_n661), .ZN(new_n878));
  XOR2_X1   g677(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n879));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n808), .B1(new_n827), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n819), .A2(new_n655), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n813), .A2(new_n652), .A3(new_n818), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n690), .B1(new_n821), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT120), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n601), .B1(new_n886), .B2(new_n859), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n503), .B1(new_n887), .B2(new_n832), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT121), .B1(new_n888), .B2(KEYINPUT57), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  INV_X1    g690(.A(new_n809), .ZN(new_n892));
  INV_X1    g691(.A(new_n857), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n856), .B1(new_n883), .B2(new_n821), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n892), .B1(new_n895), .B2(new_n820), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n896), .A2(new_n634), .B1(new_n885), .B2(new_n881), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n831), .B1(new_n897), .B2(new_n601), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n890), .B(new_n891), .C1(new_n898), .C2(new_n503), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n830), .A2(new_n832), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(KEYINPUT57), .A3(new_n463), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n889), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n865), .A2(new_n477), .A3(new_n662), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n879), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  AOI211_X1 g704(.A(KEYINPUT59), .B(new_n877), .C1(new_n864), .C2(new_n903), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n878), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT122), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n909), .B(new_n878), .C1(new_n905), .C2(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1345gat));
  AOI21_X1  g710(.A(G155gat), .B1(new_n870), .B2(new_n689), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n864), .A2(new_n866), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n689), .A2(G155gat), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(G1346gat));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n634), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G162gat), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n865), .A2(G162gat), .A3(new_n850), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n863), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1347gat));
  NAND2_X1  g719(.A1(new_n437), .A2(new_n477), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n683), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n833), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G169gat), .B1(new_n923), .B2(new_n704), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n476), .B1(new_n830), .B2(new_n832), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n470), .A2(new_n477), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n704), .A2(G169gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT123), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n923), .B2(new_n662), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n662), .A2(G176gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n928), .B2(new_n933), .ZN(G1349gat));
  NAND2_X1  g733(.A1(new_n224), .A2(new_n226), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n935), .B1(new_n923), .B2(new_n601), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n689), .A2(new_n230), .A3(new_n232), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n928), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g738(.A1(new_n927), .A2(new_n229), .A3(new_n216), .A4(new_n634), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n833), .A2(new_n634), .A3(new_n922), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT61), .ZN(new_n943));
  AND4_X1   g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .A4(G190gat), .ZN(new_n944));
  INV_X1    g743(.A(G190gat), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n946));
  AOI22_X1  g745(.A1(new_n942), .A2(new_n946), .B1(new_n941), .B2(new_n943), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n940), .B1(new_n944), .B2(new_n947), .ZN(G1351gat));
  AND4_X1   g747(.A1(new_n477), .A2(new_n925), .A3(new_n463), .A4(new_n680), .ZN(new_n949));
  AOI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n573), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n679), .A2(new_n921), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT125), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n902), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n573), .A2(G197gat), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(G1352gat));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957));
  AOI21_X1  g756(.A(G204gat), .B1(new_n957), .B2(KEYINPUT62), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n949), .A2(new_n661), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n959), .B(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(G204gat), .B1(new_n953), .B2(new_n662), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1353gat));
  NAND3_X1  g762(.A1(new_n949), .A2(new_n262), .A3(new_n689), .ZN(new_n964));
  INV_X1    g763(.A(new_n951), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n902), .A2(new_n689), .A3(new_n965), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n966), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT63), .B1(new_n966), .B2(G211gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(G1354gat));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n634), .B1(new_n954), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n972));
  OAI21_X1  g771(.A(G218gat), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n949), .A2(new_n263), .A3(new_n634), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1355gat));
endmodule


