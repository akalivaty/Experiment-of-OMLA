//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT77), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  AND3_X1   g007(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT77), .B1(new_n191), .B2(KEYINPUT16), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n189), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G128), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G128), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT24), .B(G110), .Z(new_n205));
  XNOR2_X1  g019(.A(G119), .B(G128), .ZN(new_n206));
  OAI22_X1  g020(.A1(new_n204), .A2(G110), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OR2_X1    g021(.A1(KEYINPUT64), .A2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT64), .A2(G146), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n208), .A2(new_n191), .A3(new_n193), .A4(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n197), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n204), .A2(KEYINPUT75), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT75), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n200), .A2(new_n202), .A3(new_n213), .A4(new_n203), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(G110), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(KEYINPUT76), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n205), .A2(new_n206), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n218));
  OR3_X1    g032(.A1(new_n192), .A2(KEYINPUT16), .A3(G140), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT77), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(new_n189), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n221), .B1(new_n220), .B2(new_n189), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n217), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n211), .B1(new_n216), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G137), .ZN(new_n227));
  INV_X1    g041(.A(G221), .ZN(new_n228));
  INV_X1    g042(.A(G234), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n228), .A2(new_n229), .A3(G953), .ZN(new_n230));
  XOR2_X1   g044(.A(new_n227), .B(new_n230), .Z(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n211), .B(new_n231), .C1(new_n216), .C2(new_n225), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT73), .B(G217), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n229), .B2(G902), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  OR2_X1    g055(.A1(new_n241), .A2(KEYINPUT78), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n233), .A2(new_n238), .A3(new_n234), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT25), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n233), .A2(new_n245), .A3(new_n238), .A4(new_n234), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n237), .B(KEYINPUT74), .Z(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n241), .A2(KEYINPUT78), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n242), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n251), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT11), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(G137), .ZN(new_n259));
  INV_X1    g073(.A(G137), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT11), .A3(G134), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(G137), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT65), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G131), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n263), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n262), .A2(new_n268), .A3(KEYINPUT66), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n259), .A2(new_n261), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n263), .A2(new_n265), .A3(new_n267), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n262), .A2(new_n263), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G131), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n274), .A2(KEYINPUT68), .A3(new_n276), .ZN(new_n280));
  INV_X1    g094(.A(G143), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(G146), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(KEYINPUT64), .A2(G146), .ZN(new_n284));
  NOR2_X1   g098(.A1(KEYINPUT64), .A2(G146), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n283), .B1(new_n286), .B2(G143), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT0), .A2(G128), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(KEYINPUT0), .A2(G128), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n221), .A2(G143), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n286), .B2(G143), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n287), .A2(new_n291), .B1(new_n293), .B2(new_n289), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n279), .A2(new_n280), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n260), .A2(G134), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n263), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G131), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT66), .B1(new_n262), .B2(new_n268), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n271), .A2(new_n272), .A3(new_n270), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT69), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n269), .A2(new_n273), .B1(G131), .B2(new_n297), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n306), .B1(new_n286), .B2(G143), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n287), .B1(new_n307), .B2(new_n201), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n208), .A2(G143), .A3(new_n209), .ZN(new_n309));
  INV_X1    g123(.A(new_n292), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n302), .A2(new_n305), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n199), .A2(G116), .ZN(new_n316));
  INV_X1    g130(.A(G116), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G119), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT2), .B(G113), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n319), .A2(new_n320), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n315), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OR2_X1    g138(.A1(new_n319), .A2(new_n320), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(KEYINPUT67), .A3(new_n321), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n295), .A2(new_n314), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n277), .A2(new_n294), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n313), .A2(new_n303), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n326), .A3(new_n324), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n329), .B1(new_n328), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n256), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n295), .A2(new_n314), .A3(KEYINPUT30), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n327), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n256), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n328), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT31), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n340), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT31), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n328), .A4(new_n342), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n337), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT32), .B1(new_n348), .B2(new_n349), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(new_n328), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n353), .B2(new_n256), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n330), .A2(new_n342), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT71), .B1(new_n355), .B2(new_n336), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n328), .A2(new_n335), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT28), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT71), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n342), .A4(new_n330), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n354), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n295), .A2(new_n314), .A3(new_n327), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n327), .B1(new_n295), .B2(new_n314), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT28), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n330), .A2(KEYINPUT72), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT72), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n328), .A2(new_n366), .A3(new_n329), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n342), .A2(KEYINPUT29), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n364), .A2(new_n365), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n238), .ZN(new_n370));
  OAI21_X1  g184(.A(G472), .B1(new_n361), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n250), .B1(new_n352), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(G110), .B(G140), .ZN(new_n373));
  INV_X1    g187(.A(G227), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(G953), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n373), .B(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n279), .A2(new_n280), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n379));
  INV_X1    g193(.A(G104), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT80), .A2(G104), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(G107), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n380), .A2(KEYINPUT3), .A3(G107), .ZN(new_n387));
  INV_X1    g201(.A(G107), .ZN(new_n388));
  AND2_X1   g202(.A1(KEYINPUT80), .A2(G104), .ZN(new_n389));
  NOR2_X1   g203(.A1(KEYINPUT80), .A2(G104), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n387), .B1(new_n391), .B2(KEYINPUT3), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n378), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n387), .ZN(new_n394));
  AOI21_X1  g208(.A(G107), .B1(new_n381), .B2(new_n382), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n383), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G101), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n384), .A2(KEYINPUT4), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT81), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n397), .A2(KEYINPUT81), .A3(new_n400), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n399), .B(new_n294), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n388), .A2(G104), .ZN(new_n404));
  OAI21_X1  g218(.A(G101), .B1(new_n395), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT82), .ZN(new_n406));
  INV_X1    g220(.A(new_n404), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n384), .B1(new_n391), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT82), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n406), .A2(new_n410), .B1(new_n392), .B2(new_n386), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT10), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n308), .B2(new_n312), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G128), .B1(new_n282), .B2(new_n306), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n284), .A2(new_n285), .A3(new_n281), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n415), .B1(new_n416), .B2(new_n292), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n312), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n386), .A2(new_n392), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n408), .A2(new_n409), .ZN(new_n420));
  AOI211_X1 g234(.A(KEYINPUT82), .B(new_n384), .C1(new_n391), .C2(new_n407), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n418), .B(new_n419), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n412), .ZN(new_n423));
  AND4_X1   g237(.A1(new_n377), .A2(new_n403), .A3(new_n414), .A4(new_n423), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n412), .A2(new_n422), .B1(new_n411), .B2(new_n413), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n377), .B1(new_n425), .B2(new_n403), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n376), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT85), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n377), .A2(new_n403), .A3(new_n414), .A4(new_n423), .ZN(new_n430));
  INV_X1    g244(.A(new_n376), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n274), .A2(KEYINPUT68), .A3(new_n276), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT68), .B1(new_n274), .B2(new_n276), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n422), .B1(new_n411), .B2(new_n313), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT12), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n201), .B1(new_n309), .B2(KEYINPUT1), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n440), .A2(new_n287), .B1(new_n293), .B2(new_n311), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n312), .A2(new_n417), .B1(new_n386), .B2(new_n392), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n406), .A2(new_n410), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n438), .A2(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n277), .A2(KEYINPUT12), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT84), .B1(new_n437), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT12), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n377), .B2(new_n444), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n436), .A2(KEYINPUT12), .A3(new_n277), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n432), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(KEYINPUT85), .B(new_n376), .C1(new_n424), .C2(new_n426), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n429), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G469), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n238), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n430), .B1(new_n437), .B2(new_n446), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n376), .B(KEYINPUT79), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n426), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n430), .A3(new_n431), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT83), .B1(new_n463), .B2(new_n456), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT83), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n432), .A2(new_n461), .B1(new_n458), .B2(new_n459), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n465), .B(G469), .C1(new_n466), .C2(G902), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n457), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  XOR2_X1   g282(.A(KEYINPUT9), .B(G234), .Z(new_n469));
  AOI21_X1  g283(.A(new_n228), .B1(new_n469), .B2(new_n238), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G214), .B1(G237), .B2(G902), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G122), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT8), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT5), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n316), .A2(KEYINPUT5), .ZN(new_n477));
  INV_X1    g291(.A(G113), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n323), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n480), .B(new_n419), .C1(new_n420), .C2(new_n421), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n480), .B1(new_n443), .B2(new_n419), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n475), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT87), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT87), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n486), .B(new_n475), .C1(new_n482), .C2(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n208), .A2(new_n209), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n282), .B1(new_n489), .B2(new_n281), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n192), .B(new_n312), .C1(new_n439), .C2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT88), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT7), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n491), .B(new_n493), .C1(new_n294), .C2(new_n192), .ZN(new_n494));
  INV_X1    g308(.A(G953), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G224), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT7), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n287), .A2(new_n291), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n293), .A2(new_n289), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G125), .ZN(new_n502));
  INV_X1    g316(.A(new_n497), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n502), .A2(new_n491), .A3(new_n503), .A4(new_n493), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT4), .B1(new_n506), .B2(new_n385), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n384), .B1(new_n392), .B2(new_n383), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n326), .B(new_n324), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n402), .A2(new_n401), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n482), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n505), .B1(new_n512), .B2(new_n474), .ZN(new_n513));
  AOI21_X1  g327(.A(G902), .B1(new_n488), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n402), .A2(new_n401), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n481), .B1(new_n515), .B2(new_n509), .ZN(new_n516));
  INV_X1    g330(.A(new_n474), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n481), .B(new_n474), .C1(new_n515), .C2(new_n509), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(KEYINPUT6), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n502), .A2(new_n491), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n496), .B(KEYINPUT86), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT6), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n516), .A2(new_n524), .A3(new_n517), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(G210), .B1(G237), .B2(G902), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n514), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n514), .B2(new_n526), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n473), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n191), .A2(new_n193), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n531), .ZN(new_n533));
  NOR2_X1   g347(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n532), .B(new_n286), .C1(new_n535), .C2(new_n187), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n224), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n265), .A2(new_n267), .ZN(new_n539));
  OR2_X1    g353(.A1(KEYINPUT89), .A2(G143), .ZN(new_n540));
  NAND2_X1  g354(.A1(KEYINPUT89), .A2(G143), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n540), .A2(new_n541), .B1(new_n252), .B2(G214), .ZN(new_n542));
  INV_X1    g356(.A(G237), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n495), .A3(G214), .ZN(new_n544));
  NOR2_X1   g358(.A1(KEYINPUT89), .A2(G143), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n539), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n541), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n544), .B1(new_n548), .B2(new_n545), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n265), .A2(new_n267), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n540), .A2(G214), .A3(new_n252), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(KEYINPUT18), .A2(G131), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n549), .B2(new_n551), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n192), .A2(G140), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n190), .A2(G125), .ZN(new_n557));
  OAI21_X1  g371(.A(G146), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n210), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n555), .B1(KEYINPUT90), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT90), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(new_n210), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n549), .A2(new_n554), .A3(new_n551), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n538), .A2(new_n553), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G113), .B(G122), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(new_n380), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT92), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n547), .A2(new_n569), .A3(new_n552), .ZN(new_n570));
  OAI211_X1 g384(.A(KEYINPUT17), .B(new_n539), .C1(new_n542), .C2(new_n546), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n197), .A2(new_n570), .A3(new_n222), .A4(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n555), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n559), .A2(KEYINPUT90), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n573), .A2(new_n574), .A3(new_n563), .A4(new_n562), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(new_n567), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n197), .A2(new_n553), .A3(new_n536), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n575), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT92), .ZN(new_n579));
  INV_X1    g393(.A(new_n567), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n568), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(G475), .A2(G902), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n572), .A2(new_n575), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n567), .B1(new_n577), .B2(new_n575), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n585), .A2(new_n567), .B1(new_n586), .B2(new_n579), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT93), .B1(new_n587), .B2(new_n568), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n584), .B1(new_n588), .B2(KEYINPUT20), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT20), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n582), .A2(KEYINPUT93), .A3(new_n590), .A4(new_n583), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(G116), .B(G122), .Z(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G107), .ZN(new_n594));
  XNOR2_X1  g408(.A(G116), .B(G122), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n388), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n281), .A2(G128), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n201), .A2(G143), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n594), .A2(new_n596), .B1(new_n258), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT13), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n281), .A2(KEYINPUT13), .A3(G128), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n604), .A2(new_n605), .A3(G134), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n605), .B1(new_n604), .B2(G134), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n600), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n599), .B(new_n258), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n317), .A2(KEYINPUT14), .A3(G122), .ZN(new_n610));
  OAI211_X1 g424(.A(G107), .B(new_n610), .C1(new_n593), .C2(KEYINPUT14), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n596), .A3(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n469), .A2(new_n495), .A3(new_n236), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n608), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n613), .B1(new_n608), .B2(new_n612), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n238), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT96), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n608), .A2(new_n612), .ZN(new_n619));
  INV_X1    g433(.A(new_n613), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(G902), .B1(new_n621), .B2(new_n614), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(G478), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(KEYINPUT15), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n618), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n622), .B1(KEYINPUT15), .B2(new_n625), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT94), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n572), .A2(new_n575), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n631), .B1(new_n632), .B2(new_n580), .ZN(new_n633));
  AOI211_X1 g447(.A(KEYINPUT94), .B(new_n567), .C1(new_n572), .C2(new_n575), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n576), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n238), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G475), .ZN(new_n637));
  INV_X1    g451(.A(G952), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(G953), .ZN(new_n639));
  NAND2_X1  g453(.A1(G234), .A2(G237), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n640), .A2(G902), .A3(G953), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT21), .B(G898), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n592), .A2(new_n630), .A3(new_n637), .A4(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n530), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n372), .A2(new_n472), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT97), .B(G101), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G3));
  NAND2_X1  g466(.A1(new_n348), .A2(new_n349), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(G472), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n348), .B2(new_n238), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n250), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n657), .A2(new_n658), .A3(new_n471), .A4(new_n468), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n614), .A2(KEYINPUT98), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n660), .B(KEYINPUT33), .C1(new_n615), .C2(new_n616), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT33), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n621), .B(new_n614), .C1(KEYINPUT98), .C2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n625), .A2(G902), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n618), .A2(new_n624), .A3(new_n625), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n592), .B2(new_n637), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n514), .A2(new_n526), .ZN(new_n670));
  INV_X1    g484(.A(new_n527), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n514), .A2(new_n526), .A3(new_n527), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n669), .A2(new_n674), .A3(new_n473), .A4(new_n647), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n659), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT34), .B(G104), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  NOR3_X1   g492(.A1(new_n654), .A2(new_n656), .A3(new_n250), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n473), .B(new_n647), .C1(new_n528), .C2(new_n529), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n584), .A2(new_n590), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n582), .A2(KEYINPUT20), .A3(new_n583), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n637), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n629), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n472), .A2(new_n679), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT35), .B(G107), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G9));
  NAND2_X1  g502(.A1(new_n226), .A2(KEYINPUT99), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n232), .A2(KEYINPUT36), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT99), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n691), .B(new_n211), .C1(new_n216), .C2(new_n225), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n690), .B1(new_n689), .B2(new_n692), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n240), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n248), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n472), .A2(new_n649), .A3(new_n657), .A4(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT37), .B(G110), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G12));
  INV_X1    g513(.A(KEYINPUT32), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n653), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n371), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n473), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n672), .B2(new_n673), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n696), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT100), .B(G900), .Z(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n644), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n641), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n683), .A2(new_n629), .A3(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n472), .A2(new_n703), .A3(new_n707), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G128), .ZN(G30));
  XNOR2_X1  g527(.A(new_n710), .B(KEYINPUT39), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n472), .A2(new_n714), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n715), .A2(KEYINPUT40), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(KEYINPUT40), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n674), .B(KEYINPUT38), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n362), .A2(new_n363), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n238), .B1(new_n719), .B2(new_n342), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n256), .B1(new_n345), .B2(new_n328), .ZN(new_n721));
  OAI21_X1  g535(.A(G472), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n701), .A2(new_n702), .A3(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT93), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n581), .A2(new_n576), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n586), .A2(new_n579), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n727), .A2(new_n590), .B1(new_n582), .B2(new_n583), .ZN(new_n728));
  INV_X1    g542(.A(new_n591), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n637), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n629), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n731), .A2(new_n696), .A3(new_n704), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n723), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n716), .A2(new_n717), .A3(new_n718), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT101), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G143), .ZN(G45));
  NAND2_X1  g550(.A1(new_n669), .A2(new_n710), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n472), .A2(new_n703), .A3(new_n707), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  INV_X1    g554(.A(KEYINPUT102), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n701), .A2(new_n702), .ZN(new_n742));
  INV_X1    g556(.A(new_n370), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n354), .A2(new_n356), .A3(new_n360), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n655), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n658), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n666), .A2(new_n667), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n730), .A2(new_n647), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n530), .A2(new_n748), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n455), .A2(new_n456), .A3(new_n238), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n456), .B1(new_n455), .B2(new_n238), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(new_n752), .A3(new_n471), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n741), .B1(new_n746), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n455), .A2(new_n238), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(G469), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n471), .A3(new_n457), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n675), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n372), .A2(new_n758), .A3(KEYINPUT102), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT41), .B(G113), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G15));
  NOR3_X1   g576(.A1(new_n750), .A2(new_n751), .A3(new_n470), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n703), .A2(new_n763), .A3(new_n658), .A4(new_n685), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G116), .ZN(G18));
  INV_X1    g579(.A(new_n696), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n648), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n703), .A2(new_n763), .A3(new_n705), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G119), .ZN(G21));
  NOR2_X1   g583(.A1(new_n530), .A2(new_n731), .ZN(new_n770));
  INV_X1    g584(.A(new_n349), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n344), .A2(new_n347), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n256), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n771), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n656), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n770), .A2(new_n776), .A3(new_n658), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n752), .A2(new_n471), .A3(new_n647), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT103), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n750), .A2(new_n751), .A3(new_n470), .A4(new_n646), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT103), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n775), .A2(new_n656), .A3(new_n250), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .A4(new_n770), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G122), .ZN(G24));
  NOR3_X1   g599(.A1(new_n775), .A2(new_n656), .A3(new_n766), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n763), .A3(new_n738), .A4(new_n705), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G125), .ZN(G27));
  INV_X1    g602(.A(KEYINPUT104), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n701), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n351), .A2(KEYINPUT104), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n790), .A2(new_n371), .A3(new_n702), .A4(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(G469), .B1(new_n466), .B2(G902), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n457), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n528), .A2(new_n529), .A3(new_n704), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n794), .A2(new_n471), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n792), .A2(new_n658), .A3(new_n738), .A4(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n796), .A2(new_n703), .A3(new_n658), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n799));
  AOI22_X1  g613(.A1(KEYINPUT42), .A2(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G131), .ZN(G33));
  NAND4_X1  g615(.A1(new_n796), .A2(new_n703), .A3(new_n658), .A4(new_n711), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT105), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT105), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n372), .A2(new_n804), .A3(new_n711), .A4(new_n796), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G134), .ZN(G36));
  OAI21_X1  g621(.A(new_n696), .B1(new_n654), .B2(new_n656), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT107), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n592), .A2(new_n637), .A3(new_n747), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT106), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT43), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT44), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n795), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n460), .A2(new_n462), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT45), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n456), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n818), .B2(new_n817), .ZN(new_n820));
  NAND2_X1  g634(.A1(G469), .A2(G902), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT46), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n750), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(KEYINPUT46), .A3(new_n821), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n470), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n825), .A2(new_n714), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n814), .B2(KEYINPUT44), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n816), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(new_n260), .ZN(G39));
  XNOR2_X1  g643(.A(new_n825), .B(KEYINPUT47), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n672), .A2(new_n473), .A3(new_n673), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n703), .A2(new_n658), .A3(new_n737), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G140), .ZN(G42));
  NOR4_X1   g648(.A1(new_n810), .A2(new_n250), .A3(new_n470), .A4(new_n704), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT108), .Z(new_n836));
  XOR2_X1   g650(.A(new_n752), .B(KEYINPUT49), .Z(new_n837));
  OR4_X1    g651(.A1(new_n718), .A2(new_n836), .A3(new_n723), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n764), .A2(new_n768), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n760), .A2(new_n784), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n797), .A2(KEYINPUT42), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n798), .A2(new_n799), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n649), .A2(new_n471), .A3(new_n468), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n657), .A2(new_n696), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n847), .B1(new_n746), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n680), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n730), .A2(new_n747), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n851), .B1(new_n730), .B2(new_n630), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n659), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT109), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n472), .A2(new_n679), .A3(new_n850), .A4(new_n852), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT109), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n650), .A2(new_n697), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT110), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n683), .A2(new_n630), .A3(new_n696), .A4(new_n710), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n831), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n703), .A2(new_n862), .A3(new_n471), .A4(new_n468), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n470), .B1(new_n457), .B2(new_n793), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n786), .A2(new_n738), .A3(new_n864), .A4(new_n795), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n860), .B1(new_n806), .B2(new_n867), .ZN(new_n868));
  AOI211_X1 g682(.A(KEYINPUT110), .B(new_n866), .C1(new_n805), .C2(new_n803), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n846), .B(new_n859), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n710), .B(KEYINPUT111), .Z(new_n871));
  NAND3_X1  g685(.A1(new_n248), .A2(new_n695), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT112), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n723), .A2(new_n873), .A3(new_n770), .A4(new_n864), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n712), .A2(new_n739), .A3(new_n787), .A4(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT52), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n840), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n869), .A2(new_n868), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n764), .A2(new_n768), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n754), .B2(new_n759), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n859), .A2(new_n784), .A3(new_n800), .A4(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n876), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n878), .A2(new_n882), .A3(KEYINPUT53), .A4(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n877), .A2(KEYINPUT54), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT54), .B1(new_n877), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n839), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n869), .A2(new_n868), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n881), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT53), .B1(new_n890), .B2(new_n883), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n889), .A2(new_n881), .A3(new_n876), .A4(new_n840), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n877), .A2(KEYINPUT54), .A3(new_n884), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(KEYINPUT113), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n757), .A2(new_n831), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n813), .A2(new_n642), .A3(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n792), .A2(new_n658), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT48), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n723), .A2(new_n250), .A3(new_n641), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n897), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n639), .B1(new_n903), .B2(new_n851), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n757), .A2(new_n530), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n813), .A2(new_n642), .A3(new_n782), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n904), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  OR3_X1    g722(.A1(new_n718), .A2(new_n473), .A3(new_n757), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT115), .B1(new_n909), .B2(new_n906), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT50), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n898), .A2(new_n786), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT116), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n903), .A2(new_n730), .A3(new_n747), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n830), .ZN(new_n916));
  INV_X1    g730(.A(new_n752), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(KEYINPUT114), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(KEYINPUT114), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n470), .A3(new_n919), .ZN(new_n920));
  AOI211_X1 g734(.A(new_n831), .B(new_n906), .C1(new_n916), .C2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n901), .B(new_n908), .C1(new_n922), .C2(KEYINPUT51), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(KEYINPUT51), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT117), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT117), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n926), .A3(KEYINPUT51), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n923), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n896), .A2(KEYINPUT118), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n638), .A2(new_n495), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT118), .B1(new_n896), .B2(new_n928), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n838), .B1(new_n931), .B2(new_n932), .ZN(G75));
  NAND2_X1  g747(.A1(new_n520), .A2(new_n525), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n523), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT55), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n877), .A2(new_n884), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(G210), .A3(G902), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n936), .B1(new_n939), .B2(KEYINPUT56), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n495), .A2(G952), .ZN(new_n941));
  XOR2_X1   g755(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n942));
  NOR2_X1   g756(.A1(new_n936), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT120), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G51));
  NAND2_X1  g761(.A1(new_n893), .A2(new_n894), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n821), .B(KEYINPUT57), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n455), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n937), .A2(G902), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n951), .A2(new_n820), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n941), .B1(new_n950), .B2(new_n952), .ZN(G54));
  NAND4_X1  g767(.A1(new_n937), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n954));
  INV_X1    g768(.A(new_n582), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n941), .ZN(G60));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT59), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n887), .A2(new_n895), .A3(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT122), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n664), .B(KEYINPUT121), .Z(new_n964));
  AND3_X1   g778(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n963), .B1(new_n962), .B2(new_n964), .ZN(new_n966));
  INV_X1    g780(.A(new_n941), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n964), .A2(new_n960), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n948), .B2(new_n968), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n965), .A2(new_n966), .A3(new_n969), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT60), .Z(new_n972));
  NOR2_X1   g786(.A1(new_n693), .A2(new_n694), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT123), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n937), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n937), .A2(new_n972), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n967), .B(new_n975), .C1(new_n976), .C2(new_n235), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT61), .Z(G66));
  INV_X1    g792(.A(G224), .ZN(new_n979));
  OAI21_X1  g793(.A(G953), .B1(new_n645), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n842), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n859), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n980), .B1(new_n983), .B2(G953), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n934), .B1(G898), .B2(new_n495), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT124), .Z(new_n986));
  XNOR2_X1  g800(.A(new_n984), .B(new_n986), .ZN(G69));
  NAND2_X1  g801(.A1(new_n334), .A2(new_n339), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n338), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n532), .B1(new_n535), .B2(new_n187), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(G900), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(G953), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT126), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n833), .B1(new_n816), .B2(new_n827), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n826), .A2(new_n770), .A3(new_n899), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n712), .A2(new_n739), .A3(new_n787), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n996), .A2(new_n997), .A3(new_n800), .A4(new_n806), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n991), .B(new_n994), .C1(new_n999), .C2(G953), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n735), .A2(new_n997), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(KEYINPUT62), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT62), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n735), .A2(new_n1003), .A3(new_n997), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n372), .A2(new_n795), .A3(new_n852), .ZN(new_n1005));
  OAI221_X1 g819(.A(new_n833), .B1(new_n715), .B2(new_n1005), .C1(new_n816), .C2(new_n827), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1002), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n495), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT125), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1000), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n991), .B1(new_n1009), .B2(KEYINPUT125), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(G953), .B1(new_n374), .B2(new_n992), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1012), .A2(new_n1014), .A3(KEYINPUT127), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(KEYINPUT127), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n1015), .A2(KEYINPUT127), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1017), .B(new_n1018), .C1(new_n1013), .C2(new_n1011), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n1016), .A2(new_n1019), .ZN(G72));
  INV_X1    g834(.A(new_n721), .ZN(new_n1021));
  OR2_X1    g835(.A1(new_n1008), .A2(new_n982), .ZN(new_n1022));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  AOI21_X1  g838(.A(new_n1021), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n345), .A2(new_n328), .A3(new_n256), .ZN(new_n1026));
  AND4_X1   g840(.A1(new_n1021), .A2(new_n937), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1024), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(new_n999), .B2(new_n983), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n967), .B1(new_n1029), .B2(new_n1026), .ZN(new_n1030));
  NOR3_X1   g844(.A1(new_n1025), .A2(new_n1027), .A3(new_n1030), .ZN(G57));
endmodule


