//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G116), .A2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n202), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n216), .C1(G97), .C2(G257), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G1), .B2(G20), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  INV_X1    g0019(.A(KEYINPUT64), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(KEYINPUT64), .A2(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G1), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n228), .A2(new_n221), .A3(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT0), .Z(new_n231));
  NOR3_X1   g0031(.A1(new_n219), .A2(new_n227), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND2_X1  g0047(.A1(new_n203), .A2(G20), .ZN(new_n248));
  INV_X1    g0048(.A(G150), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n224), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT70), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(KEYINPUT8), .B(G58), .Z(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n248), .B1(new_n249), .B2(new_n251), .C1(new_n254), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n225), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n228), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n202), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n259), .B1(new_n228), .B2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G50), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n260), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT9), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G222), .A3(new_n271), .ZN(new_n272));
  XOR2_X1   g0072(.A(new_n272), .B(KEYINPUT68), .Z(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n277), .A3(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT69), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n270), .A2(new_n280), .A3(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n281), .A3(G223), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(new_n207), .B2(new_n270), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n269), .B1(new_n273), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n228), .B(G274), .C1(G41), .C2(G45), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT66), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT65), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT65), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(G33), .A3(G41), .ZN(new_n290));
  INV_X1    g0090(.A(new_n225), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT67), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G41), .A2(G45), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(G1), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n228), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n292), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G226), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n284), .A2(new_n286), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(G200), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n260), .A2(KEYINPUT9), .A3(new_n263), .A4(new_n265), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n268), .A2(new_n301), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n266), .B1(new_n299), .B2(G179), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(new_n299), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n292), .A2(G238), .A3(new_n295), .A4(new_n296), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n286), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n269), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n213), .A2(new_n271), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n270), .B(new_n317), .C1(G232), .C2(new_n271), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT73), .ZN(new_n319));
  INV_X1    g0119(.A(G97), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n274), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n316), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n313), .B1(new_n315), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT74), .B1(new_n315), .B2(new_n324), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n315), .A2(new_n324), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT13), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n325), .B(new_n326), .C1(new_n328), .C2(KEYINPUT74), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G179), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT76), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n328), .A2(new_n325), .A3(G169), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n333), .A2(KEYINPUT14), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n329), .A2(KEYINPUT76), .A3(G179), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(KEYINPUT14), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n332), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n221), .A2(G68), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(new_n228), .A3(G13), .ZN(new_n339));
  XOR2_X1   g0139(.A(new_n339), .B(KEYINPUT12), .Z(new_n340));
  INV_X1    g0140(.A(new_n338), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n251), .A2(new_n202), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n341), .B(new_n343), .C1(new_n254), .C2(new_n207), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n259), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT11), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT11), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(new_n347), .A3(new_n259), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n340), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n264), .A2(G68), .ZN(new_n350));
  XOR2_X1   g0150(.A(new_n350), .B(KEYINPUT75), .Z(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n337), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n328), .A2(G200), .A3(new_n325), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n329), .A2(G190), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n349), .A2(new_n351), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n255), .A2(new_n262), .ZN(new_n358));
  INV_X1    g0158(.A(new_n264), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(new_n255), .ZN(new_n360));
  INV_X1    g0160(.A(new_n259), .ZN(new_n361));
  AND2_X1   g0161(.A1(G58), .A2(G68), .ZN(new_n362));
  OAI21_X1  g0162(.A(G20), .B1(new_n362), .B2(new_n201), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT78), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n250), .A2(G159), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n364), .B1(new_n363), .B2(new_n365), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n275), .A2(new_n277), .B1(new_n222), .B2(new_n223), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT77), .B1(new_n369), .B2(KEYINPUT7), .ZN(new_n370));
  INV_X1    g0170(.A(new_n270), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT77), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT7), .ZN(new_n374));
  AND2_X1   g0174(.A1(KEYINPUT64), .A2(G20), .ZN(new_n375));
  NOR2_X1   g0175(.A1(KEYINPUT64), .A2(G20), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n373), .B(new_n374), .C1(new_n377), .C2(new_n270), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n370), .A2(new_n372), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n368), .B1(new_n379), .B2(G68), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n361), .B1(new_n380), .B2(KEYINPUT16), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT79), .B1(new_n276), .B2(G33), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT79), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(new_n274), .A3(KEYINPUT3), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n385), .A3(new_n277), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n374), .B1(new_n270), .B2(G20), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n214), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n363), .A2(new_n365), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n382), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n360), .B1(new_n381), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n213), .A2(G1698), .ZN(new_n393));
  OR2_X1    g0193(.A1(G223), .A2(G1698), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n270), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n316), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n292), .A2(G232), .A3(new_n295), .A4(new_n296), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n398), .A2(G179), .A3(new_n286), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n286), .A2(new_n399), .ZN(new_n401));
  OAI21_X1  g0201(.A(G169), .B1(new_n401), .B2(new_n397), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT18), .B1(new_n392), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n379), .A2(G68), .ZN(new_n406));
  INV_X1    g0206(.A(new_n368), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(KEYINPUT16), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(new_n259), .A3(new_n391), .ZN(new_n409));
  INV_X1    g0209(.A(new_n360), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(new_n403), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT80), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(KEYINPUT17), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n398), .A2(new_n286), .A3(new_n399), .ZN(new_n416));
  INV_X1    g0216(.A(G200), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n416), .B2(G190), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n392), .B2(new_n419), .ZN(new_n420));
  XOR2_X1   g0220(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n421));
  AND4_X1   g0221(.A1(new_n410), .A2(new_n409), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n405), .B(new_n413), .C1(new_n420), .C2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT72), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n279), .A2(new_n281), .A3(G238), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n371), .A2(G107), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n270), .A2(G232), .A3(new_n271), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT71), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n270), .A2(KEYINPUT71), .A3(G232), .A4(new_n271), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n425), .A2(new_n426), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n269), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n297), .A2(G244), .ZN(new_n433));
  AND4_X1   g0233(.A1(new_n424), .A2(new_n432), .A3(new_n286), .A4(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n286), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n431), .B2(new_n269), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n424), .B1(new_n436), .B2(new_n433), .ZN(new_n437));
  OAI21_X1  g0237(.A(G179), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n432), .A2(new_n286), .A3(new_n433), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT72), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n436), .A2(new_n424), .A3(new_n433), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(G169), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n261), .A2(G77), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n359), .A2(new_n207), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n255), .A2(new_n250), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT15), .B(G87), .ZN(new_n447));
  OAI221_X1 g0247(.A(new_n446), .B1(new_n207), .B2(new_n224), .C1(new_n252), .C2(new_n447), .ZN(new_n448));
  AOI211_X1 g0248(.A(new_n444), .B(new_n445), .C1(new_n448), .C2(new_n259), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(G190), .B1(new_n434), .B2(new_n437), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n440), .A2(G200), .A3(new_n441), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(new_n449), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n312), .A2(new_n357), .A3(new_n423), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT81), .ZN(new_n457));
  INV_X1    g0257(.A(G41), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n228), .A2(G45), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(KEYINPUT5), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT5), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G41), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(KEYINPUT81), .A3(new_n228), .A4(G45), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n461), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n292), .A2(G274), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n461), .A2(new_n462), .A3(new_n465), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(G270), .A3(new_n292), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n271), .A2(G257), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G264), .A2(G1698), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n275), .A2(new_n277), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(new_n269), .C1(G303), .C2(new_n270), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n469), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n262), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n228), .A2(G33), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n361), .A2(G116), .A3(new_n261), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  OAI221_X1 g0282(.A(new_n482), .B1(G33), .B2(new_n320), .C1(new_n375), .C2(new_n376), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n258), .A2(new_n225), .B1(G20), .B2(new_n478), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n483), .A2(KEYINPUT20), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT20), .B1(new_n483), .B2(new_n484), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n479), .B(new_n481), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n477), .A2(G179), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n476), .A2(G200), .ZN(new_n489));
  INV_X1    g0289(.A(new_n487), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n489), .B(new_n490), .C1(new_n300), .C2(new_n476), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT21), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n475), .B1(new_n470), .B2(new_n467), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n309), .B1(new_n494), .B2(new_n471), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n492), .B1(new_n495), .B2(new_n487), .ZN(new_n496));
  AND4_X1   g0296(.A1(new_n492), .A2(new_n476), .A3(new_n487), .A4(G169), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n488), .B(new_n491), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT89), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n476), .A2(G169), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT21), .B1(new_n500), .B2(new_n490), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n495), .A2(new_n492), .A3(new_n487), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT89), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(new_n488), .A4(new_n491), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n275), .B(new_n277), .C1(G250), .C2(G1698), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n271), .A2(G257), .ZN(new_n508));
  INV_X1    g0308(.A(G294), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n507), .A2(new_n508), .B1(new_n274), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n269), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n470), .A2(G264), .A3(new_n292), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n469), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n417), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(G190), .B2(new_n513), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n361), .A2(new_n261), .A3(new_n480), .ZN(new_n516));
  INV_X1    g0316(.A(G107), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT92), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT25), .ZN(new_n520));
  AOI211_X1 g0320(.A(G107), .B(new_n261), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n275), .B(new_n277), .C1(new_n375), .C2(new_n376), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(new_n209), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NOR4_X1   g0331(.A1(new_n527), .A2(new_n209), .A3(new_n526), .A4(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT24), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n221), .A2(G33), .A3(G116), .ZN(new_n535));
  XOR2_X1   g0335(.A(KEYINPUT91), .B(KEYINPUT23), .Z(new_n536));
  NAND2_X1  g0336(.A1(new_n517), .A2(G20), .ZN(new_n537));
  NOR2_X1   g0337(.A1(KEYINPUT23), .A2(G107), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n536), .A2(new_n537), .B1(new_n377), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n533), .A2(new_n534), .A3(new_n535), .A4(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n527), .ZN(new_n541));
  INV_X1    g0341(.A(new_n526), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n541), .A2(G87), .A3(new_n542), .A4(new_n530), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n543), .A2(new_n535), .A3(new_n528), .A4(new_n539), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT24), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n515), .B(new_n525), .C1(new_n546), .C2(new_n361), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n513), .A2(new_n309), .ZN(new_n548));
  INV_X1    g0348(.A(G179), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n469), .A2(new_n511), .A3(new_n512), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n361), .B1(new_n540), .B2(new_n545), .ZN(new_n553));
  INV_X1    g0353(.A(new_n525), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G33), .B(G97), .C1(new_n375), .C2(new_n376), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n224), .A2(new_n270), .A3(G68), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR3_X1   g0360(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n321), .A2(KEYINPUT19), .A3(new_n322), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(new_n224), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n259), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n447), .A2(new_n262), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT86), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n564), .A2(KEYINPUT86), .A3(new_n565), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n460), .A2(G274), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n460), .A2(new_n210), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n292), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n215), .A2(new_n271), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n208), .A2(G1698), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(new_n270), .B1(G33), .B2(G116), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n573), .B1(new_n577), .B2(new_n316), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G200), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n516), .A2(new_n209), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G190), .B(new_n573), .C1(new_n577), .C2(new_n316), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT88), .ZN(new_n583));
  XNOR2_X1  g0383(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n570), .A2(new_n579), .A3(new_n581), .A4(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n564), .A2(KEYINPUT86), .A3(new_n565), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT86), .B1(new_n564), .B2(new_n565), .ZN(new_n587));
  XOR2_X1   g0387(.A(new_n447), .B(KEYINPUT87), .Z(new_n588));
  OAI22_X1  g0388(.A1(new_n586), .A2(new_n587), .B1(new_n516), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n573), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n270), .A2(new_n574), .A3(new_n575), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G116), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n316), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(G169), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT85), .ZN(new_n595));
  OAI211_X1 g0395(.A(G179), .B(new_n573), .C1(new_n577), .C2(new_n316), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n595), .B1(new_n594), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n589), .A2(new_n599), .ZN(new_n600));
  AND4_X1   g0400(.A1(new_n547), .A2(new_n555), .A3(new_n585), .A4(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n470), .A2(G257), .A3(new_n292), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT82), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT82), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n470), .A2(new_n604), .A3(G257), .A4(new_n292), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n275), .A2(new_n277), .A3(G244), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT4), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n607), .A2(new_n608), .B1(G33), .B2(G283), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n608), .B1(new_n270), .B2(G250), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n609), .B(new_n610), .C1(new_n271), .C2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(new_n269), .B1(new_n466), .B2(new_n468), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n606), .A2(G190), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n607), .A2(new_n608), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n610), .A2(new_n615), .A3(new_n482), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n270), .A2(G250), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n271), .B1(new_n617), .B2(KEYINPUT4), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n269), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n619), .A2(new_n603), .A3(new_n469), .A4(new_n605), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G200), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n262), .A2(new_n320), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n516), .B2(new_n320), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n387), .A2(new_n388), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G107), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n250), .A2(G77), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n517), .A2(KEYINPUT6), .A3(G97), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n320), .A2(new_n517), .ZN(new_n628));
  NOR2_X1   g0428(.A1(G97), .A2(G107), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n627), .B1(new_n630), .B2(KEYINPUT6), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n377), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n625), .A2(new_n626), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n623), .B1(new_n633), .B2(new_n259), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n614), .A2(new_n621), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT84), .B1(new_n620), .B2(G179), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT84), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n606), .A2(new_n637), .A3(new_n549), .A4(new_n613), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n620), .A2(new_n309), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n624), .A2(G107), .B1(new_n377), .B2(new_n631), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n361), .B1(new_n641), .B2(new_n626), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT83), .B1(new_n642), .B2(new_n623), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n633), .A2(new_n259), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT83), .ZN(new_n645));
  INV_X1    g0445(.A(new_n623), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n635), .B1(new_n640), .B2(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n456), .A2(new_n506), .A3(new_n601), .A4(new_n649), .ZN(G372));
  NAND2_X1  g0450(.A1(new_n405), .A2(new_n413), .ZN(new_n651));
  INV_X1    g0451(.A(new_n356), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n353), .B1(new_n652), .B2(new_n451), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n392), .A2(new_n419), .A3(new_n421), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n409), .A2(new_n410), .A3(new_n419), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n656), .B2(new_n415), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n651), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n307), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n311), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n640), .A2(new_n585), .A3(new_n600), .A4(new_n648), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT26), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n570), .A2(new_n579), .A3(new_n581), .A4(new_n582), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n594), .A2(new_n596), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n589), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n634), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n662), .A2(new_n670), .A3(new_n665), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n555), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n503), .A2(new_n488), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT93), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n490), .A2(new_n549), .A3(new_n476), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n501), .B2(new_n502), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT93), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n673), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n614), .A2(new_n621), .A3(new_n634), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n645), .B1(new_n644), .B2(new_n646), .ZN(new_n683));
  AOI211_X1 g0483(.A(KEYINPUT83), .B(new_n623), .C1(new_n633), .C2(new_n259), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n682), .B1(new_n685), .B2(new_n668), .ZN(new_n686));
  INV_X1    g0486(.A(new_n547), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n663), .A2(new_n665), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n681), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n672), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n660), .B1(new_n456), .B2(new_n691), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT94), .Z(G369));
  INV_X1    g0493(.A(G13), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n377), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  OR3_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .A3(G1), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT27), .B1(new_n696), .B2(G1), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G213), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n487), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT95), .B1(new_n506), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n676), .A2(new_n679), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n702), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n704), .A2(KEYINPUT95), .A3(new_n702), .ZN(new_n707));
  OR3_X1    g0507(.A1(new_n706), .A2(KEYINPUT96), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT96), .B1(new_n706), .B2(new_n707), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n701), .B1(new_n553), .B2(new_n554), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n547), .A2(new_n555), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n701), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n711), .B1(new_n555), .B2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n708), .A2(G330), .A3(new_n709), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n674), .A2(new_n712), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n711), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n673), .B2(new_n712), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n229), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G1), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n561), .A2(new_n478), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n722), .A2(new_n723), .B1(new_n226), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n649), .A2(new_n547), .A3(new_n666), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n680), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n726), .B(new_n712), .C1(new_n728), .C2(new_n671), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT100), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n678), .A2(new_n555), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n730), .B1(new_n678), .B2(new_n555), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n689), .A2(new_n733), .B1(new_n589), .B2(new_n664), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n666), .A2(KEYINPUT99), .A3(new_n669), .A4(KEYINPUT26), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT99), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n661), .B2(new_n667), .ZN(new_n737));
  NOR4_X1   g0537(.A1(new_n688), .A2(new_n667), .A3(new_n668), .A4(new_n634), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n701), .B1(new_n734), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n729), .B1(new_n740), .B2(new_n726), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n606), .A2(new_n477), .A3(new_n613), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n511), .A2(new_n512), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n745), .A2(new_n596), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n743), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n476), .A2(new_n549), .A3(new_n578), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT97), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT97), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n476), .A2(new_n750), .A3(new_n549), .A4(new_n578), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n749), .A2(new_n513), .A3(new_n620), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n747), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OR3_X1    g0554(.A1(new_n744), .A2(new_n743), .A3(new_n746), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n712), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n506), .A2(new_n601), .A3(new_n649), .A4(new_n712), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(new_n757), .B2(KEYINPUT31), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n753), .A2(KEYINPUT98), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT98), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n747), .A2(new_n752), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n759), .A2(new_n755), .A3(new_n761), .ZN(new_n762));
  AND3_X1   g0562(.A1(new_n762), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n763));
  OAI21_X1  g0563(.A(G330), .B1(new_n758), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n742), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n725), .B1(new_n766), .B2(G1), .ZN(G364));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n706), .A2(new_n707), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n722), .B1(G45), .B2(new_n695), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n224), .A2(new_n549), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(new_n300), .A3(new_n417), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n300), .A2(new_n417), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n776), .A2(G311), .B1(new_n779), .B2(G326), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n300), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n549), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n377), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n780), .B1(new_n509), .B2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT104), .Z(new_n786));
  NAND2_X1  g0586(.A1(new_n774), .A2(new_n781), .ZN(new_n787));
  INV_X1    g0587(.A(G322), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n371), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n377), .A2(new_n549), .A3(new_n300), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G329), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n790), .A2(new_n417), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G283), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n774), .A2(new_n300), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n417), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT105), .B(KEYINPUT33), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(G317), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n789), .B(new_n796), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G303), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n777), .A2(G20), .A3(new_n549), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n786), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n794), .A2(new_n517), .B1(new_n778), .B2(new_n202), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n803), .A2(new_n209), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n371), .B(new_n806), .C1(G97), .C2(new_n783), .ZN(new_n807));
  INV_X1    g0607(.A(new_n798), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n214), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT101), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n787), .B(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n805), .B(new_n809), .C1(G58), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n776), .A2(KEYINPUT102), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT102), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n775), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n813), .B1(new_n207), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n791), .A2(G159), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT103), .Z(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT32), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n804), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n225), .B1(G20), .B2(new_n309), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n770), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n719), .A2(new_n270), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n226), .A2(G45), .ZN(new_n826));
  INV_X1    g0626(.A(G45), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n825), .B(new_n826), .C1(new_n243), .C2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n270), .A2(new_n229), .A3(G355), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(G116), .C2(new_n229), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n822), .A2(new_n823), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n772), .A2(new_n773), .A3(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n708), .A2(new_n709), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(G330), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n708), .A2(G330), .A3(new_n709), .ZN(new_n835));
  INV_X1    g0635(.A(new_n773), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n832), .B1(new_n834), .B2(new_n837), .ZN(G396));
  OAI21_X1  g0638(.A(KEYINPUT109), .B1(new_n451), .B2(new_n712), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n449), .B1(new_n438), .B2(new_n442), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT109), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n840), .A2(new_n841), .A3(new_n701), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT108), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n452), .A2(new_n449), .A3(new_n453), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(new_n840), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n450), .A2(new_n701), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AND4_X1   g0648(.A1(new_n844), .A2(new_n451), .A3(new_n454), .A4(new_n847), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n843), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n712), .B1(new_n728), .B2(new_n671), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n850), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(new_n764), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n836), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n817), .A2(new_n478), .B1(new_n795), .B2(new_n808), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT106), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n794), .A2(new_n209), .ZN(new_n857));
  INV_X1    g0657(.A(new_n803), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n270), .B1(new_n858), .B2(G107), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n859), .B1(new_n320), .B2(new_n784), .C1(new_n802), .C2(new_n778), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n857), .B(new_n860), .C1(G311), .C2(new_n791), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n856), .B(new_n861), .C1(new_n509), .C2(new_n787), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n812), .A2(G143), .B1(G150), .B2(new_n798), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n779), .A2(G137), .ZN(new_n864));
  INV_X1    g0664(.A(G159), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n863), .B(new_n864), .C1(new_n865), .C2(new_n817), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT34), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  INV_X1    g0669(.A(G58), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n270), .B1(new_n784), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n794), .A2(new_n214), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n871), .B(new_n872), .C1(G132), .C2(new_n791), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n202), .B2(new_n803), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT107), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n868), .A2(new_n869), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n874), .A2(new_n875), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n862), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n823), .A2(new_n768), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n879), .A2(new_n823), .B1(new_n207), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n881), .B(new_n773), .C1(new_n850), .C2(new_n769), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n854), .A2(new_n882), .ZN(G384));
  NAND2_X1  g0683(.A1(new_n352), .A2(new_n701), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n353), .A2(new_n884), .A3(new_n356), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n352), .B(new_n701), .C1(new_n652), .C2(new_n337), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n756), .A2(KEYINPUT31), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n850), .B(new_n887), .C1(new_n758), .C2(new_n889), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n655), .A2(KEYINPUT112), .ZN(new_n891));
  INV_X1    g0691(.A(new_n699), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n403), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n655), .B(KEYINPUT112), .C1(new_n392), .C2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n891), .A2(new_n894), .A3(KEYINPUT37), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n655), .B(new_n896), .C1(new_n392), .C2(new_n893), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT111), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n404), .A2(new_n699), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT37), .B1(new_n411), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT111), .B1(new_n901), .B2(new_n655), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n895), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n423), .A2(new_n411), .A3(new_n892), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n897), .A2(new_n898), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n901), .A2(KEYINPUT111), .A3(new_n655), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n408), .A2(new_n259), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n380), .A2(KEYINPUT16), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n410), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT110), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(KEYINPUT110), .B(new_n410), .C1(new_n909), .C2(new_n910), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(new_n900), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n655), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT37), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n412), .B1(new_n411), .B2(new_n403), .ZN(new_n918));
  AOI211_X1 g0718(.A(KEYINPUT18), .B(new_n404), .C1(new_n409), .C2(new_n410), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n699), .B1(new_n920), .B2(new_n657), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n406), .A2(new_n407), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n382), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n360), .B1(new_n923), .B2(new_n381), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(new_n912), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n908), .A2(new_n917), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n905), .B1(KEYINPUT38), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT40), .B1(new_n890), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n885), .A2(new_n886), .ZN(new_n929));
  INV_X1    g0729(.A(new_n758), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n929), .B1(new_n930), .B2(new_n888), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT38), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n916), .A2(KEYINPUT37), .B1(new_n906), .B2(new_n907), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n423), .A2(new_n892), .A3(new_n925), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n420), .A2(new_n422), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n892), .B(new_n925), .C1(new_n936), .C2(new_n651), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n899), .A2(new_n902), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n896), .B1(new_n915), .B2(new_n655), .ZN(new_n939));
  OAI211_X1 g0739(.A(KEYINPUT38), .B(new_n937), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT40), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n931), .A2(new_n941), .A3(new_n942), .A4(new_n850), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n928), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n930), .A2(new_n888), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n456), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(G330), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  INV_X1    g0749(.A(new_n940), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n905), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n353), .A2(new_n701), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n935), .A2(KEYINPUT39), .A3(new_n940), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n651), .A2(new_n699), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n451), .A2(new_n701), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n846), .A2(new_n844), .A3(new_n847), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n451), .A2(new_n454), .A3(new_n847), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT108), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n958), .A2(new_n960), .B1(new_n839), .B2(new_n842), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n957), .B1(new_n961), .B2(new_n851), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(new_n941), .A3(new_n887), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n954), .A2(new_n955), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n660), .B1(new_n741), .B2(new_n456), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n948), .B(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n228), .B2(new_n695), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n291), .B(new_n377), .C1(new_n631), .C2(KEYINPUT35), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n478), .B(new_n969), .C1(KEYINPUT35), .C2(new_n631), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT36), .Z(new_n971));
  OAI21_X1  g0771(.A(G77), .B1(new_n870), .B2(new_n214), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n972), .A2(new_n226), .B1(G50), .B2(new_n214), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(G1), .A3(new_n694), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n968), .A2(new_n971), .A3(new_n974), .ZN(G367));
  OAI21_X1  g0775(.A(new_n649), .B1(new_n634), .B2(new_n712), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n669), .A2(new_n701), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n714), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n570), .A2(new_n581), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n701), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n980), .A2(new_n665), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n666), .B2(new_n980), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n976), .A2(new_n977), .ZN(new_n985));
  AND3_X1   g0785(.A1(new_n985), .A2(KEYINPUT42), .A3(new_n716), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT42), .B1(new_n985), .B2(new_n716), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n555), .B1(new_n976), .B2(new_n977), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n640), .A2(new_n648), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n712), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n984), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT43), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n994), .B2(new_n982), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n992), .B(new_n984), .C1(new_n986), .C2(new_n987), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT113), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n978), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT114), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n995), .A2(new_n998), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(new_n978), .ZN(new_n1003));
  OAI21_X1  g0803(.A(G1), .B1(new_n696), .B2(new_n827), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(KEYINPUT115), .B(KEYINPUT41), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n720), .B(new_n1005), .Z(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n716), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n715), .B(new_n711), .C1(new_n555), .C2(new_n712), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n833), .A2(G330), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n835), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n717), .A2(new_n985), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT45), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n717), .A2(new_n985), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT44), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n714), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n714), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1016), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1013), .A2(new_n766), .A3(new_n1019), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1007), .B1(new_n1023), .B2(new_n766), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1001), .B(new_n1003), .C1(new_n1004), .C2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n784), .A2(new_n214), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n270), .B1(new_n870), .B2(new_n803), .C1(new_n808), .C2(new_n865), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(G137), .C2(new_n791), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n779), .A2(G143), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n817), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(G50), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n787), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1032), .A2(G150), .B1(new_n793), .B2(G77), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n858), .A2(G116), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT46), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n270), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n517), .B2(new_n784), .C1(new_n808), .C2(new_n509), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n794), .A2(new_n320), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n791), .ZN(new_n1040));
  INV_X1    g0840(.A(G317), .ZN(new_n1041));
  INV_X1    g0841(.A(G311), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1040), .A2(new_n1041), .B1(new_n778), .B2(new_n1042), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1038), .A2(new_n1039), .A3(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n795), .B2(new_n817), .C1(new_n802), .C2(new_n811), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1034), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT116), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT47), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n836), .B1(new_n1049), .B2(new_n823), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n825), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n824), .B1(new_n229), .B2(new_n447), .C1(new_n239), .C2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(new_n771), .C2(new_n983), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1025), .A2(new_n1053), .ZN(G387));
  OAI22_X1  g0854(.A1(new_n817), .A2(new_n802), .B1(new_n811), .B2(new_n1041), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT118), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1055), .A2(new_n1056), .B1(new_n1042), .B2(new_n808), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n788), .B2(new_n778), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT48), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n783), .A2(G283), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n858), .A2(G294), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT49), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n791), .A2(G326), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n270), .B1(new_n793), .B2(G116), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n588), .A2(new_n784), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n865), .B2(new_n778), .C1(new_n249), .C2(new_n1040), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G50), .B2(new_n1032), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n775), .A2(new_n214), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1073), .B(new_n1039), .C1(new_n255), .C2(new_n798), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1072), .B(new_n1074), .C1(new_n207), .C2(new_n803), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1069), .B1(new_n371), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n823), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n713), .A2(new_n771), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n255), .A2(new_n202), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n723), .B1(new_n1079), .B2(KEYINPUT50), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1080), .B(new_n827), .C1(KEYINPUT50), .C2(new_n1079), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G68), .B2(G77), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n825), .B1(new_n236), .B2(new_n827), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n723), .A2(new_n229), .A3(new_n270), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n229), .A2(G107), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n824), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1077), .A2(new_n773), .A3(new_n1078), .A4(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1013), .A2(new_n766), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1011), .A2(new_n765), .A3(new_n1012), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n720), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1013), .A2(new_n1004), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT117), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT117), .B1(new_n1013), .B2(new_n1004), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(KEYINPUT119), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1093), .B(new_n1094), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT119), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1099), .A2(new_n1100), .A3(new_n1091), .A4(new_n1088), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(G393));
  NAND2_X1  g0902(.A1(new_n1022), .A2(new_n1019), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1089), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n720), .A3(new_n1023), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1022), .A2(new_n1004), .A3(new_n1019), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n371), .B1(new_n803), .B2(new_n795), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n794), .A2(new_n517), .B1(new_n478), .B2(new_n784), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(G322), .C2(new_n791), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n776), .A2(G294), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1042), .A2(new_n787), .B1(new_n778), .B2(new_n1041), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT52), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n798), .A2(G303), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n371), .B1(new_n858), .B2(G68), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n207), .B2(new_n784), .C1(new_n808), .C2(new_n202), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n857), .B(new_n1116), .C1(G143), .C2(new_n791), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n256), .B2(new_n817), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n249), .A2(new_n778), .B1(new_n787), .B2(new_n865), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT51), .Z(new_n1120));
  OAI21_X1  g0920(.A(new_n1114), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n836), .B1(new_n1121), .B2(new_n823), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n824), .B1(new_n320), .B2(new_n229), .C1(new_n246), .C2(new_n1051), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(new_n771), .C2(new_n985), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1105), .A2(new_n1106), .A3(new_n1124), .ZN(G390));
  INV_X1    g0925(.A(new_n905), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n952), .B1(new_n1126), .B2(new_n940), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n956), .B1(new_n740), .B2(new_n850), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n929), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n764), .A2(new_n961), .A3(new_n929), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n935), .A2(KEYINPUT39), .A3(new_n940), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT39), .B1(new_n1126), .B2(new_n940), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n952), .B1(new_n962), .B2(new_n887), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1129), .B(new_n1131), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT120), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(G330), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n890), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n962), .A2(new_n887), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n952), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1141), .A2(new_n1142), .B1(new_n951), .B2(new_n953), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1129), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1140), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n701), .B1(new_n672), .B2(new_n690), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n956), .B1(new_n1146), .B2(new_n850), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1142), .B1(new_n1147), .B2(new_n929), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n951), .A2(new_n953), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1150), .A2(KEYINPUT120), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1138), .A2(new_n1145), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(G330), .B1(new_n758), .B2(new_n889), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(KEYINPUT121), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT121), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(G330), .C1(new_n758), .C2(new_n889), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n850), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n929), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1128), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(new_n1130), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n764), .A2(new_n961), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1162), .A2(new_n887), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n962), .B1(new_n1163), .B2(new_n1140), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n945), .A2(new_n456), .A3(G330), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n965), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1152), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1167), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1171), .A2(new_n1145), .A3(new_n1138), .A4(new_n1151), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n720), .A3(new_n1172), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1138), .A2(new_n1145), .A3(new_n1151), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1040), .A2(new_n509), .B1(new_n778), .B2(new_n795), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n872), .B(new_n1175), .C1(G116), .C2(new_n1032), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n371), .B1(new_n784), .B2(new_n207), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n806), .B(new_n1177), .C1(new_n798), .C2(G107), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1176), .B(new_n1178), .C1(new_n320), .C2(new_n817), .ZN(new_n1179));
  INV_X1    g0979(.A(G132), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n787), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(G125), .ZN(new_n1182));
  INV_X1    g0982(.A(G128), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1040), .A2(new_n1182), .B1(new_n778), .B2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1181), .B(new_n1184), .C1(G50), .C2(new_n793), .ZN(new_n1185));
  XOR2_X1   g0985(.A(KEYINPUT54), .B(G143), .Z(new_n1186));
  NAND2_X1  g0986(.A1(new_n1030), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n784), .A2(new_n865), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n858), .A2(G150), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n270), .B1(new_n1189), .B2(KEYINPUT53), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1188), .B(new_n1190), .C1(G137), .C2(new_n798), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(KEYINPUT53), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1185), .A2(new_n1187), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1179), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n823), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n880), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1195), .B1(new_n255), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1149), .B2(new_n768), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1174), .A2(new_n1004), .B1(new_n773), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1173), .A2(new_n1199), .ZN(G378));
  AND3_X1   g1000(.A1(new_n964), .A2(G330), .A3(new_n944), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1139), .B1(new_n928), .B2(new_n943), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1202), .A2(new_n964), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n312), .B(KEYINPUT55), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n266), .A2(new_n892), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT56), .Z(new_n1206));
  XNOR2_X1  g1006(.A(new_n1204), .B(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1201), .A2(new_n1203), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n944), .A2(G330), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n964), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1202), .A2(new_n964), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1207), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1004), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1032), .A2(G128), .B1(new_n858), .B2(new_n1186), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT122), .Z(new_n1217));
  OAI22_X1  g1017(.A1(new_n808), .A2(new_n1180), .B1(new_n249), .B2(new_n784), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G137), .B2(new_n776), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1217), .B(new_n1219), .C1(new_n1182), .C2(new_n778), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1220), .B(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(G33), .B1(new_n793), .B2(G159), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G41), .B1(new_n791), .B2(G124), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G41), .B1(new_n858), .B2(G77), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n478), .B2(new_n778), .C1(new_n808), .C2(new_n320), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1032), .A2(G107), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1026), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n793), .A2(G58), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n791), .A2(G283), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n588), .A2(new_n775), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1227), .A2(new_n1232), .A3(new_n270), .A4(new_n1233), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT58), .Z(new_n1235));
  AOI21_X1  g1035(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1225), .B(new_n1235), .C1(G50), .C2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n836), .B1(new_n1237), .B2(new_n823), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(G50), .B2(new_n1196), .C1(new_n1208), .C2(new_n769), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1215), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1168), .B1(new_n1152), .B2(new_n1169), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1208), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1212), .A2(new_n1207), .A3(new_n1213), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1242), .A2(new_n1245), .A3(KEYINPUT57), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n720), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT57), .B1(new_n1242), .B2(new_n1245), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1241), .B1(new_n1247), .B2(new_n1248), .ZN(G375));
  NAND3_X1  g1049(.A1(new_n1161), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1169), .A2(new_n1006), .A3(new_n1250), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n817), .A2(new_n517), .B1(new_n478), .B2(new_n808), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT124), .Z(new_n1253));
  OAI221_X1 g1053(.A(new_n371), .B1(new_n320), .B2(new_n803), .C1(new_n794), .C2(new_n207), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1070), .B1(new_n509), .B2(new_n778), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1254), .B(new_n1255), .C1(G303), .C2(new_n791), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1253), .B(new_n1256), .C1(new_n795), .C2(new_n787), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1230), .B1(new_n1180), .B2(new_n778), .C1(new_n1040), .C2(new_n1183), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G137), .B2(new_n812), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n270), .B1(new_n803), .B2(new_n865), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n798), .B2(new_n1186), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n775), .A2(new_n249), .B1(new_n202), .B2(new_n784), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT125), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1259), .A2(new_n1261), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1257), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n823), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(G68), .B2(new_n1196), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n836), .B(new_n1267), .C1(new_n768), .C2(new_n929), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1165), .B2(new_n1004), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1251), .A2(new_n1269), .ZN(G381));
  NAND2_X1  g1070(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT57), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n720), .A3(new_n1246), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(G378), .A2(new_n1240), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(G390), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1025), .A3(new_n1053), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1278), .A2(G384), .A3(G381), .ZN(new_n1279));
  INV_X1    g1079(.A(G396), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1098), .A2(new_n1101), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1276), .A2(new_n1279), .A3(new_n1281), .ZN(G407));
  INV_X1    g1082(.A(G213), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(new_n1276), .B2(new_n700), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(G407), .ZN(G409));
  INV_X1    g1085(.A(G378), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1172), .A2(new_n1168), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1006), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1286), .A2(new_n1241), .A3(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1283), .A2(G343), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n721), .B1(new_n1287), .B2(KEYINPUT57), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1240), .B1(new_n1292), .B2(new_n1273), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1289), .B(new_n1291), .C1(new_n1293), .C2(new_n1286), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT60), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1250), .A2(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1161), .A2(new_n1167), .A3(new_n1164), .A4(KEYINPUT60), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1296), .A2(new_n1169), .A3(new_n720), .A4(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(G384), .A3(new_n1269), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT126), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1269), .ZN(new_n1301));
  INV_X1    g1101(.A(G384), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1298), .A2(new_n1304), .A3(G384), .A4(new_n1269), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1300), .A2(new_n1303), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1290), .A2(G2897), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1307), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1300), .A2(new_n1303), .A3(new_n1305), .A4(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT61), .B1(new_n1294), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(G375), .A2(G378), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1290), .B1(new_n1275), .B2(new_n1288), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1306), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT62), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1313), .A2(new_n1314), .A3(new_n1318), .A4(new_n1315), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1312), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1278), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1277), .B1(new_n1025), .B2(new_n1053), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1280), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1323));
  OAI22_X1  g1123(.A1(new_n1321), .A2(new_n1322), .B1(new_n1281), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G393), .A2(G396), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(G387), .A2(G390), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1098), .A2(new_n1101), .A3(new_n1280), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1325), .A2(new_n1326), .A3(new_n1278), .A4(new_n1327), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1324), .A2(new_n1328), .A3(KEYINPUT127), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT127), .B1(new_n1324), .B2(new_n1328), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1320), .A2(new_n1331), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1313), .A2(new_n1314), .A3(KEYINPUT63), .A4(new_n1315), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT61), .B1(new_n1324), .B2(new_n1328), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1335), .B1(new_n1294), .B2(new_n1311), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1316), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1333), .B(new_n1334), .C1(new_n1336), .C2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1332), .A2(new_n1338), .ZN(G405));
  NAND2_X1  g1139(.A1(new_n1324), .A2(new_n1328), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1286), .B1(new_n1274), .B2(new_n1241), .ZN(new_n1341));
  OR2_X1    g1141(.A1(new_n1276), .A2(new_n1341), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1342), .A2(new_n1315), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1276), .A2(new_n1341), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1344), .A2(new_n1306), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1340), .B1(new_n1343), .B2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1342), .A2(new_n1315), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1344), .A2(new_n1306), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1347), .A2(new_n1328), .A3(new_n1324), .A4(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1346), .A2(new_n1349), .ZN(G402));
endmodule


