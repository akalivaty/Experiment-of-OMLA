

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743;

  INV_X1 U371 ( .A(G953), .ZN(n470) );
  NOR2_X2 U372 ( .A1(n551), .A2(n550), .ZN(n572) );
  XNOR2_X2 U373 ( .A(n361), .B(n359), .ZN(n691) );
  NOR2_X2 U374 ( .A1(n675), .A2(n679), .ZN(n361) );
  XNOR2_X2 U375 ( .A(n494), .B(KEYINPUT0), .ZN(n525) );
  NOR2_X2 U376 ( .A1(n568), .A2(n493), .ZN(n494) );
  XNOR2_X2 U377 ( .A(n400), .B(G143), .ZN(n456) );
  NOR2_X1 U378 ( .A1(n740), .A2(n639), .ZN(n532) );
  NOR2_X2 U379 ( .A1(n673), .A2(n528), .ZN(n512) );
  AND2_X2 U380 ( .A1(n375), .A2(n352), .ZN(n708) );
  XNOR2_X1 U381 ( .A(n496), .B(KEYINPUT22), .ZN(n508) );
  XNOR2_X1 U382 ( .A(n401), .B(KEYINPUT110), .ZN(n675) );
  NAND2_X1 U383 ( .A1(n523), .A2(n521), .ZN(n679) );
  INV_X1 U384 ( .A(G128), .ZN(n400) );
  XNOR2_X1 U385 ( .A(G902), .B(KEYINPUT15), .ZN(n606) );
  BUF_X1 U386 ( .A(n708), .Z(n712) );
  INV_X1 U387 ( .A(n508), .ZN(n392) );
  NAND2_X1 U388 ( .A1(n570), .A2(n569), .ZN(n644) );
  NOR2_X1 U389 ( .A1(n656), .A2(n554), .ZN(n555) );
  XNOR2_X1 U390 ( .A(n724), .B(n427), .ZN(n476) );
  XNOR2_X1 U391 ( .A(n456), .B(KEYINPUT4), .ZN(n404) );
  XNOR2_X1 U392 ( .A(n398), .B(G125), .ZN(n478) );
  XNOR2_X1 U393 ( .A(n351), .B(n426), .ZN(n724) );
  XOR2_X1 U394 ( .A(G101), .B(KEYINPUT64), .Z(n477) );
  XOR2_X1 U395 ( .A(G104), .B(G107), .Z(n351) );
  XNOR2_X1 U396 ( .A(G110), .B(KEYINPUT74), .ZN(n426) );
  NOR2_X1 U397 ( .A1(n620), .A2(n716), .ZN(n621) );
  NOR2_X1 U398 ( .A1(n630), .A2(n716), .ZN(n632) );
  NOR2_X1 U399 ( .A1(n613), .A2(n716), .ZN(n614) );
  XNOR2_X2 U400 ( .A(n539), .B(n538), .ZN(n717) );
  NOR2_X2 U401 ( .A1(n537), .A2(n536), .ZN(n539) );
  XNOR2_X1 U402 ( .A(n404), .B(n432), .ZN(n732) );
  XNOR2_X1 U403 ( .A(KEYINPUT67), .B(G137), .ZN(n430) );
  XOR2_X1 U404 ( .A(G131), .B(G134), .Z(n431) );
  NAND2_X1 U405 ( .A1(n369), .A2(n368), .ZN(n378) );
  XNOR2_X1 U406 ( .A(n436), .B(n435), .ZN(n560) );
  XNOR2_X1 U407 ( .A(n434), .B(G469), .ZN(n435) );
  INV_X1 U408 ( .A(KEYINPUT81), .ZN(n364) );
  AND2_X1 U409 ( .A1(n509), .A2(n532), .ZN(n516) );
  INV_X1 U410 ( .A(G146), .ZN(n398) );
  XNOR2_X1 U411 ( .A(n574), .B(KEYINPUT38), .ZN(n678) );
  XNOR2_X1 U412 ( .A(n506), .B(KEYINPUT104), .ZN(n507) );
  INV_X1 U413 ( .A(KEYINPUT6), .ZN(n506) );
  NOR2_X1 U414 ( .A1(G953), .A2(G237), .ZN(n497) );
  XNOR2_X1 U415 ( .A(n442), .B(n441), .ZN(n443) );
  INV_X1 U416 ( .A(G104), .ZN(n441) );
  XNOR2_X1 U417 ( .A(n478), .B(n397), .ZN(n731) );
  XNOR2_X1 U418 ( .A(KEYINPUT10), .B(G140), .ZN(n397) );
  XNOR2_X1 U419 ( .A(n503), .B(n402), .ZN(n703) );
  XNOR2_X1 U420 ( .A(n476), .B(n403), .ZN(n402) );
  XNOR2_X1 U421 ( .A(n429), .B(n428), .ZN(n403) );
  NAND2_X1 U422 ( .A1(n379), .A2(n376), .ZN(n375) );
  NAND2_X1 U423 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U424 ( .A1(n381), .A2(n380), .ZN(n379) );
  XNOR2_X1 U425 ( .A(n455), .B(n454), .ZN(n523) );
  BUF_X1 U426 ( .A(n557), .Z(n365) );
  AND2_X1 U427 ( .A1(n612), .A2(G953), .ZN(n716) );
  XNOR2_X1 U428 ( .A(n388), .B(n387), .ZN(n740) );
  INV_X1 U429 ( .A(KEYINPUT32), .ZN(n387) );
  NAND2_X1 U430 ( .A1(n392), .A2(n356), .ZN(n388) );
  XNOR2_X1 U431 ( .A(n363), .B(n362), .ZN(n588) );
  INV_X1 U432 ( .A(KEYINPUT80), .ZN(n362) );
  XNOR2_X1 U433 ( .A(KEYINPUT78), .B(n547), .ZN(n554) );
  XNOR2_X1 U434 ( .A(n366), .B(KEYINPUT107), .ZN(n544) );
  XOR2_X1 U435 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n417) );
  XOR2_X1 U436 ( .A(KEYINPUT100), .B(KEYINPUT98), .Z(n440) );
  XNOR2_X1 U437 ( .A(G143), .B(G131), .ZN(n442) );
  XNOR2_X1 U438 ( .A(n732), .B(n433), .ZN(n503) );
  XNOR2_X1 U439 ( .A(KEYINPUT18), .B(KEYINPUT90), .ZN(n472) );
  XNOR2_X1 U440 ( .A(KEYINPUT17), .B(KEYINPUT77), .ZN(n473) );
  XNOR2_X1 U441 ( .A(n370), .B(n482), .ZN(n383) );
  INV_X1 U442 ( .A(n404), .ZN(n370) );
  INV_X1 U443 ( .A(KEYINPUT82), .ZN(n377) );
  NAND2_X1 U444 ( .A1(G234), .A2(G237), .ZN(n488) );
  INV_X1 U445 ( .A(G237), .ZN(n483) );
  INV_X1 U446 ( .A(G902), .ZN(n484) );
  AND2_X1 U447 ( .A1(n542), .A2(n396), .ZN(n549) );
  INV_X1 U448 ( .A(n554), .ZN(n396) );
  INV_X1 U449 ( .A(KEYINPUT76), .ZN(n548) );
  INV_X1 U450 ( .A(KEYINPUT88), .ZN(n390) );
  XOR2_X1 U451 ( .A(G110), .B(G137), .Z(n412) );
  XNOR2_X1 U452 ( .A(G119), .B(G128), .ZN(n411) );
  XNOR2_X1 U453 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n414) );
  XNOR2_X1 U454 ( .A(n395), .B(n552), .ZN(n598) );
  AND2_X1 U455 ( .A1(n572), .A2(n678), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n371), .B(n405), .ZN(n673) );
  INV_X1 U457 ( .A(KEYINPUT33), .ZN(n405) );
  AND2_X1 U458 ( .A1(n562), .A2(n561), .ZN(n570) );
  NOR2_X1 U459 ( .A1(n560), .A2(n661), .ZN(n542) );
  XNOR2_X1 U460 ( .A(n451), .B(n450), .ZN(n609) );
  XNOR2_X1 U461 ( .A(n394), .B(n393), .ZN(n742) );
  INV_X1 U462 ( .A(KEYINPUT40), .ZN(n393) );
  NOR2_X1 U463 ( .A1(n598), .A2(n645), .ZN(n394) );
  OR2_X1 U464 ( .A1(n523), .A2(n522), .ZN(n645) );
  NAND2_X1 U465 ( .A1(n662), .A2(n386), .ZN(n385) );
  NOR2_X1 U466 ( .A1(n518), .A2(n365), .ZN(n386) );
  XNOR2_X1 U467 ( .A(n374), .B(n373), .ZN(n372) );
  XNOR2_X1 U468 ( .A(n704), .B(n707), .ZN(n373) );
  NAND2_X1 U469 ( .A1(n712), .A2(G469), .ZN(n374) );
  INV_X1 U470 ( .A(G143), .ZN(n624) );
  AND2_X1 U471 ( .A1(n391), .A2(n358), .ZN(n350) );
  XNOR2_X1 U472 ( .A(n557), .B(n507), .ZN(n578) );
  OR2_X1 U473 ( .A1(n697), .A2(n696), .ZN(n352) );
  AND2_X1 U474 ( .A1(n540), .A2(KEYINPUT82), .ZN(n353) );
  AND2_X1 U475 ( .A1(n586), .A2(n582), .ZN(n354) );
  AND2_X1 U476 ( .A1(n485), .A2(G210), .ZN(n355) );
  AND2_X1 U477 ( .A1(n354), .A2(n657), .ZN(n356) );
  AND2_X1 U478 ( .A1(n582), .A2(n390), .ZN(n357) );
  OR2_X1 U479 ( .A1(n582), .A2(n390), .ZN(n358) );
  XOR2_X1 U480 ( .A(n553), .B(KEYINPUT41), .Z(n359) );
  XOR2_X1 U481 ( .A(G122), .B(KEYINPUT126), .Z(n360) );
  NAND2_X1 U482 ( .A1(n576), .A2(n577), .ZN(n363) );
  NOR2_X1 U483 ( .A1(n713), .A2(G902), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n420), .B(n421), .ZN(n713) );
  XNOR2_X1 U485 ( .A(n571), .B(n364), .ZN(n577) );
  NOR2_X1 U486 ( .A1(n543), .A2(n470), .ZN(n366) );
  NAND2_X1 U487 ( .A1(n678), .A2(n677), .ZN(n401) );
  NAND2_X1 U488 ( .A1(n367), .A2(n696), .ZN(n381) );
  NAND2_X1 U489 ( .A1(n353), .A2(n369), .ZN(n367) );
  XNOR2_X1 U490 ( .A(n383), .B(n475), .ZN(n382) );
  XNOR2_X2 U491 ( .A(n519), .B(KEYINPUT106), .ZN(n743) );
  NOR2_X1 U492 ( .A1(n717), .A2(n606), .ZN(n368) );
  INV_X1 U493 ( .A(n607), .ZN(n369) );
  XNOR2_X1 U494 ( .A(n733), .B(KEYINPUT75), .ZN(n607) );
  NAND2_X1 U495 ( .A1(n527), .A2(n578), .ZN(n371) );
  AND2_X1 U496 ( .A1(n438), .A2(n406), .ZN(n527) );
  NOR2_X1 U497 ( .A1(n372), .A2(n716), .ZN(G54) );
  INV_X1 U498 ( .A(n606), .ZN(n380) );
  NAND2_X1 U499 ( .A1(n615), .A2(n606), .ZN(n399) );
  XNOR2_X1 U500 ( .A(n382), .B(n384), .ZN(n615) );
  XNOR2_X1 U501 ( .A(n476), .B(n725), .ZN(n384) );
  XNOR2_X1 U502 ( .A(n498), .B(n481), .ZN(n725) );
  NOR2_X1 U503 ( .A1(n508), .A2(n385), .ZN(n639) );
  NOR2_X1 U504 ( .A1(n579), .A2(n558), .ZN(n559) );
  NAND2_X1 U505 ( .A1(n350), .A2(n389), .ZN(n409) );
  NAND2_X1 U506 ( .A1(n392), .A2(n357), .ZN(n389) );
  NAND2_X1 U507 ( .A1(n508), .A2(KEYINPUT88), .ZN(n391) );
  NAND2_X1 U508 ( .A1(n510), .A2(n511), .ZN(n661) );
  XNOR2_X2 U509 ( .A(n399), .B(n355), .ZN(n583) );
  XNOR2_X1 U510 ( .A(n531), .B(n360), .ZN(G24) );
  XNOR2_X1 U511 ( .A(n531), .B(KEYINPUT65), .ZN(n515) );
  INV_X1 U512 ( .A(n438), .ZN(n662) );
  INV_X1 U513 ( .A(n661), .ZN(n406) );
  AND2_X1 U514 ( .A1(n676), .A2(KEYINPUT47), .ZN(n407) );
  XNOR2_X1 U515 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n408) );
  OR2_X1 U516 ( .A1(n676), .A2(n530), .ZN(n410) );
  NOR2_X1 U517 ( .A1(n623), .A2(n407), .ZN(n576) );
  INV_X1 U518 ( .A(KEYINPUT69), .ZN(n434) );
  INV_X1 U519 ( .A(KEYINPUT5), .ZN(n500) );
  XNOR2_X1 U520 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U521 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U522 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U523 ( .A(n423), .B(KEYINPUT25), .ZN(n424) );
  BUF_X1 U524 ( .A(n574), .Z(n602) );
  INV_X1 U525 ( .A(KEYINPUT44), .ZN(n509) );
  XNOR2_X1 U526 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U527 ( .A(n731), .B(n413), .ZN(n421) );
  XNOR2_X1 U528 ( .A(n414), .B(KEYINPUT94), .ZN(n415) );
  XOR2_X1 U529 ( .A(KEYINPUT23), .B(n415), .Z(n419) );
  NAND2_X1 U530 ( .A1(G234), .A2(n470), .ZN(n416) );
  XNOR2_X1 U531 ( .A(n417), .B(n416), .ZN(n460) );
  NAND2_X1 U532 ( .A1(G221), .A2(n460), .ZN(n418) );
  XNOR2_X1 U533 ( .A(n419), .B(n418), .ZN(n420) );
  NAND2_X1 U534 ( .A1(n606), .A2(G234), .ZN(n422) );
  XNOR2_X1 U535 ( .A(n422), .B(KEYINPUT20), .ZN(n466) );
  NAND2_X1 U536 ( .A1(n466), .A2(G217), .ZN(n423) );
  XNOR2_X1 U537 ( .A(n425), .B(n424), .ZN(n510) );
  INV_X1 U538 ( .A(n510), .ZN(n657) );
  INV_X1 U539 ( .A(n657), .ZN(n518) );
  INV_X1 U540 ( .A(G140), .ZN(n428) );
  INV_X1 U541 ( .A(KEYINPUT70), .ZN(n427) );
  NAND2_X1 U542 ( .A1(G227), .A2(n470), .ZN(n429) );
  XNOR2_X1 U543 ( .A(G146), .B(n477), .ZN(n433) );
  XNOR2_X1 U544 ( .A(n431), .B(n430), .ZN(n432) );
  NOR2_X1 U545 ( .A1(n703), .A2(G902), .ZN(n436) );
  INV_X1 U546 ( .A(KEYINPUT1), .ZN(n437) );
  XNOR2_X1 U547 ( .A(n560), .B(n437), .ZN(n438) );
  XNOR2_X1 U548 ( .A(KEYINPUT11), .B(KEYINPUT99), .ZN(n439) );
  XNOR2_X1 U549 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U550 ( .A(n731), .B(n445), .Z(n451) );
  XOR2_X1 U551 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n447) );
  XNOR2_X1 U552 ( .A(G113), .B(G122), .ZN(n446) );
  XNOR2_X1 U553 ( .A(n447), .B(n446), .ZN(n449) );
  NAND2_X1 U554 ( .A1(G214), .A2(n497), .ZN(n448) );
  NOR2_X1 U555 ( .A1(n609), .A2(G902), .ZN(n455) );
  XOR2_X1 U556 ( .A(KEYINPUT13), .B(KEYINPUT101), .Z(n453) );
  XNOR2_X1 U557 ( .A(KEYINPUT102), .B(G475), .ZN(n452) );
  XOR2_X1 U558 ( .A(n453), .B(n452), .Z(n454) );
  XNOR2_X1 U559 ( .A(G134), .B(KEYINPUT9), .ZN(n459) );
  XNOR2_X1 U560 ( .A(n456), .B(G116), .ZN(n457) );
  XNOR2_X1 U561 ( .A(n457), .B(G107), .ZN(n458) );
  XNOR2_X1 U562 ( .A(n459), .B(n458), .ZN(n464) );
  XOR2_X1 U563 ( .A(G122), .B(KEYINPUT7), .Z(n462) );
  NAND2_X1 U564 ( .A1(G217), .A2(n460), .ZN(n461) );
  XNOR2_X1 U565 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U566 ( .A(n464), .B(n463), .ZN(n709) );
  NOR2_X1 U567 ( .A1(G902), .A2(n709), .ZN(n465) );
  XNOR2_X1 U568 ( .A(G478), .B(n465), .ZN(n521) );
  INV_X1 U569 ( .A(n679), .ZN(n468) );
  NAND2_X1 U570 ( .A1(G221), .A2(n466), .ZN(n467) );
  XNOR2_X1 U571 ( .A(KEYINPUT21), .B(n467), .ZN(n656) );
  XOR2_X1 U572 ( .A(KEYINPUT96), .B(n656), .Z(n511) );
  NAND2_X1 U573 ( .A1(n468), .A2(n511), .ZN(n469) );
  XNOR2_X1 U574 ( .A(n469), .B(KEYINPUT105), .ZN(n495) );
  NAND2_X1 U575 ( .A1(n470), .A2(G224), .ZN(n471) );
  XNOR2_X1 U576 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U577 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U578 ( .A(n478), .B(n477), .ZN(n482) );
  XNOR2_X1 U579 ( .A(G116), .B(G113), .ZN(n480) );
  XNOR2_X1 U580 ( .A(KEYINPUT3), .B(G119), .ZN(n479) );
  XNOR2_X1 U581 ( .A(n480), .B(n479), .ZN(n498) );
  XNOR2_X1 U582 ( .A(KEYINPUT16), .B(G122), .ZN(n481) );
  NAND2_X1 U583 ( .A1(n484), .A2(n483), .ZN(n485) );
  NAND2_X1 U584 ( .A1(n485), .A2(G214), .ZN(n677) );
  NAND2_X1 U585 ( .A1(n583), .A2(n677), .ZN(n487) );
  INV_X1 U586 ( .A(KEYINPUT19), .ZN(n486) );
  XNOR2_X1 U587 ( .A(n487), .B(n486), .ZN(n568) );
  XNOR2_X1 U588 ( .A(n488), .B(KEYINPUT14), .ZN(n490) );
  NAND2_X1 U589 ( .A1(G952), .A2(n490), .ZN(n688) );
  NOR2_X1 U590 ( .A1(n688), .A2(G953), .ZN(n489) );
  XNOR2_X1 U591 ( .A(n489), .B(KEYINPUT92), .ZN(n545) );
  NAND2_X1 U592 ( .A1(G902), .A2(n490), .ZN(n543) );
  NOR2_X1 U593 ( .A1(G898), .A2(n470), .ZN(n491) );
  XNOR2_X1 U594 ( .A(KEYINPUT93), .B(n491), .ZN(n728) );
  NOR2_X1 U595 ( .A1(n543), .A2(n728), .ZN(n492) );
  NOR2_X1 U596 ( .A1(n545), .A2(n492), .ZN(n493) );
  NAND2_X1 U597 ( .A1(n495), .A2(n525), .ZN(n496) );
  NAND2_X1 U598 ( .A1(n497), .A2(G210), .ZN(n499) );
  XOR2_X1 U599 ( .A(n499), .B(n498), .Z(n501) );
  XNOR2_X1 U600 ( .A(n503), .B(n502), .ZN(n627) );
  NOR2_X1 U601 ( .A1(n627), .A2(G902), .ZN(n505) );
  XNOR2_X1 U602 ( .A(G472), .B(KEYINPUT71), .ZN(n504) );
  XNOR2_X1 U603 ( .A(n505), .B(n504), .ZN(n557) );
  INV_X1 U604 ( .A(n662), .ZN(n586) );
  INV_X1 U605 ( .A(n525), .ZN(n528) );
  XNOR2_X1 U606 ( .A(n512), .B(KEYINPUT34), .ZN(n513) );
  NOR2_X1 U607 ( .A1(n523), .A2(n521), .ZN(n573) );
  NAND2_X1 U608 ( .A1(n513), .A2(n573), .ZN(n514) );
  XNOR2_X2 U609 ( .A(n514), .B(KEYINPUT35), .ZN(n531) );
  NAND2_X1 U610 ( .A1(n516), .A2(n515), .ZN(n520) );
  NOR2_X1 U611 ( .A1(n586), .A2(n409), .ZN(n517) );
  NAND2_X1 U612 ( .A1(n518), .A2(n517), .ZN(n519) );
  NAND2_X1 U613 ( .A1(n520), .A2(n743), .ZN(n537) );
  INV_X1 U614 ( .A(n521), .ZN(n522) );
  AND2_X1 U615 ( .A1(n523), .A2(n522), .ZN(n650) );
  INV_X1 U616 ( .A(n650), .ZN(n640) );
  NAND2_X1 U617 ( .A1(n640), .A2(n645), .ZN(n524) );
  XNOR2_X1 U618 ( .A(n524), .B(KEYINPUT103), .ZN(n676) );
  NAND2_X1 U619 ( .A1(n542), .A2(n525), .ZN(n526) );
  NOR2_X1 U620 ( .A1(n365), .A2(n526), .ZN(n635) );
  NAND2_X1 U621 ( .A1(n365), .A2(n527), .ZN(n667) );
  NOR2_X1 U622 ( .A1(n528), .A2(n667), .ZN(n529) );
  XOR2_X1 U623 ( .A(KEYINPUT31), .B(n529), .Z(n651) );
  NOR2_X1 U624 ( .A1(n635), .A2(n651), .ZN(n530) );
  NOR2_X1 U625 ( .A1(n531), .A2(KEYINPUT65), .ZN(n533) );
  NAND2_X1 U626 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U627 ( .A1(n534), .A2(KEYINPUT44), .ZN(n535) );
  NAND2_X1 U628 ( .A1(n410), .A2(n535), .ZN(n536) );
  XNOR2_X1 U629 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n538) );
  INV_X1 U630 ( .A(n717), .ZN(n540) );
  NAND2_X1 U631 ( .A1(n557), .A2(n677), .ZN(n541) );
  XNOR2_X1 U632 ( .A(KEYINPUT30), .B(n541), .ZN(n551) );
  NOR2_X1 U633 ( .A1(G900), .A2(n544), .ZN(n546) );
  NOR2_X1 U634 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U635 ( .A(n549), .B(n548), .ZN(n550) );
  INV_X1 U636 ( .A(n583), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT87), .B(KEYINPUT39), .Z(n552) );
  INV_X1 U638 ( .A(KEYINPUT111), .ZN(n553) );
  NAND2_X1 U639 ( .A1(n555), .A2(n657), .ZN(n556) );
  XNOR2_X1 U640 ( .A(n556), .B(KEYINPUT68), .ZN(n579) );
  INV_X1 U641 ( .A(n557), .ZN(n558) );
  XNOR2_X1 U642 ( .A(n559), .B(KEYINPUT28), .ZN(n562) );
  XNOR2_X1 U643 ( .A(n560), .B(KEYINPUT109), .ZN(n561) );
  NAND2_X1 U644 ( .A1(n691), .A2(n570), .ZN(n564) );
  XNOR2_X1 U645 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n563) );
  XNOR2_X1 U646 ( .A(n564), .B(n563), .ZN(n625) );
  NAND2_X1 U647 ( .A1(n742), .A2(n625), .ZN(n567) );
  INV_X1 U648 ( .A(KEYINPUT86), .ZN(n565) );
  XNOR2_X1 U649 ( .A(n565), .B(KEYINPUT46), .ZN(n566) );
  XNOR2_X1 U650 ( .A(n567), .B(n566), .ZN(n595) );
  INV_X1 U651 ( .A(n568), .ZN(n569) );
  NAND2_X1 U652 ( .A1(n644), .A2(KEYINPUT47), .ZN(n571) );
  NAND2_X1 U653 ( .A1(n573), .A2(n572), .ZN(n575) );
  NOR2_X1 U654 ( .A1(n575), .A2(n602), .ZN(n623) );
  INV_X1 U655 ( .A(n578), .ZN(n582) );
  NOR2_X1 U656 ( .A1(n579), .A2(n645), .ZN(n580) );
  NAND2_X1 U657 ( .A1(n580), .A2(n677), .ZN(n581) );
  NOR2_X1 U658 ( .A1(n582), .A2(n581), .ZN(n599) );
  NAND2_X1 U659 ( .A1(n599), .A2(n583), .ZN(n585) );
  INV_X1 U660 ( .A(KEYINPUT36), .ZN(n584) );
  XNOR2_X1 U661 ( .A(n585), .B(n584), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n587), .A2(n586), .ZN(n654) );
  NAND2_X1 U663 ( .A1(n588), .A2(n654), .ZN(n593) );
  NOR2_X1 U664 ( .A1(n676), .A2(KEYINPUT47), .ZN(n589) );
  XNOR2_X1 U665 ( .A(n589), .B(KEYINPUT73), .ZN(n590) );
  NOR2_X1 U666 ( .A1(n590), .A2(n644), .ZN(n591) );
  XNOR2_X1 U667 ( .A(n591), .B(KEYINPUT72), .ZN(n592) );
  NOR2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n597) );
  XNOR2_X1 U670 ( .A(KEYINPUT85), .B(KEYINPUT48), .ZN(n596) );
  XNOR2_X1 U671 ( .A(n597), .B(n596), .ZN(n605) );
  OR2_X1 U672 ( .A1(n598), .A2(n640), .ZN(n655) );
  NAND2_X1 U673 ( .A1(n599), .A2(n662), .ZN(n601) );
  XNOR2_X1 U674 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n600) );
  XNOR2_X1 U675 ( .A(n601), .B(n600), .ZN(n603) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n622) );
  AND2_X1 U677 ( .A1(n655), .A2(n622), .ZN(n604) );
  AND2_X2 U678 ( .A1(n605), .A2(n604), .ZN(n733) );
  INV_X1 U679 ( .A(n733), .ZN(n608) );
  OR2_X1 U680 ( .A1(n717), .A2(n608), .ZN(n697) );
  INV_X1 U681 ( .A(KEYINPUT2), .ZN(n696) );
  NAND2_X1 U682 ( .A1(n708), .A2(G475), .ZN(n611) );
  XNOR2_X1 U683 ( .A(n609), .B(n408), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n611), .B(n610), .ZN(n613) );
  INV_X1 U685 ( .A(G952), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U687 ( .A1(n708), .A2(G210), .ZN(n619) );
  XNOR2_X1 U688 ( .A(KEYINPUT55), .B(KEYINPUT79), .ZN(n616) );
  XOR2_X1 U689 ( .A(n616), .B(KEYINPUT54), .Z(n617) );
  XNOR2_X1 U690 ( .A(n615), .B(n617), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U692 ( .A(n621), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U693 ( .A(n622), .B(G140), .ZN(G42) );
  XNOR2_X1 U694 ( .A(n624), .B(n623), .ZN(G45) );
  XNOR2_X1 U695 ( .A(n625), .B(G137), .ZN(G39) );
  NAND2_X1 U696 ( .A1(n708), .A2(G472), .ZN(n629) );
  XOR2_X1 U697 ( .A(KEYINPUT91), .B(KEYINPUT62), .Z(n626) );
  XNOR2_X1 U698 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U700 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(G57) );
  XOR2_X1 U702 ( .A(G104), .B(KEYINPUT113), .Z(n634) );
  INV_X1 U703 ( .A(n645), .ZN(n647) );
  NAND2_X1 U704 ( .A1(n635), .A2(n647), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n634), .B(n633), .ZN(G6) );
  XOR2_X1 U706 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n637) );
  NAND2_X1 U707 ( .A1(n635), .A2(n650), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U709 ( .A(G107), .B(n638), .ZN(G9) );
  XOR2_X1 U710 ( .A(G110), .B(n639), .Z(G12) );
  NOR2_X1 U711 ( .A1(n640), .A2(n644), .ZN(n642) );
  XNOR2_X1 U712 ( .A(KEYINPUT114), .B(KEYINPUT29), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U714 ( .A(G128), .B(n643), .ZN(G30) );
  NOR2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U716 ( .A(G146), .B(n646), .Z(G48) );
  XOR2_X1 U717 ( .A(G113), .B(KEYINPUT115), .Z(n649) );
  NAND2_X1 U718 ( .A1(n651), .A2(n647), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n649), .B(n648), .ZN(G15) );
  NAND2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U721 ( .A(n652), .B(G116), .ZN(G18) );
  XOR2_X1 U722 ( .A(G125), .B(KEYINPUT37), .Z(n653) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(G27) );
  XNOR2_X1 U724 ( .A(G134), .B(n655), .ZN(G36) );
  AND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U726 ( .A(KEYINPUT49), .B(n658), .Z(n659) );
  NOR2_X1 U727 ( .A1(n365), .A2(n659), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n660), .B(KEYINPUT116), .ZN(n666) );
  XOR2_X1 U729 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n664) );
  NAND2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n668) );
  NAND2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U734 ( .A(KEYINPUT51), .B(n669), .ZN(n670) );
  XNOR2_X1 U735 ( .A(n670), .B(KEYINPUT118), .ZN(n672) );
  INV_X1 U736 ( .A(n691), .ZN(n671) );
  NOR2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n685) );
  BUF_X1 U738 ( .A(n673), .Z(n674) );
  NOR2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n682) );
  NOR2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n680) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U743 ( .A1(n674), .A2(n683), .ZN(n684) );
  NOR2_X1 U744 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U745 ( .A(n686), .B(KEYINPUT52), .ZN(n687) );
  NOR2_X1 U746 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U747 ( .A(KEYINPUT119), .B(n689), .Z(n690) );
  NOR2_X1 U748 ( .A1(G953), .A2(n690), .ZN(n695) );
  INV_X1 U749 ( .A(n674), .ZN(n692) );
  NAND2_X1 U750 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U751 ( .A(n693), .B(KEYINPUT120), .ZN(n694) );
  NAND2_X1 U752 ( .A1(n695), .A2(n694), .ZN(n701) );
  NAND2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U754 ( .A1(n352), .A2(n698), .ZN(n699) );
  XNOR2_X1 U755 ( .A(KEYINPUT83), .B(n699), .ZN(n700) );
  NOR2_X1 U756 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U757 ( .A(KEYINPUT53), .B(n702), .ZN(G75) );
  INV_X1 U758 ( .A(n703), .ZN(n704) );
  XOR2_X1 U759 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n706) );
  XNOR2_X1 U760 ( .A(KEYINPUT122), .B(KEYINPUT121), .ZN(n705) );
  XNOR2_X1 U761 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U762 ( .A1(n712), .A2(G478), .ZN(n710) );
  XNOR2_X1 U763 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n716), .A2(n711), .ZN(G63) );
  NAND2_X1 U765 ( .A1(n712), .A2(G217), .ZN(n714) );
  XNOR2_X1 U766 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U767 ( .A1(n716), .A2(n715), .ZN(G66) );
  OR2_X1 U768 ( .A1(n717), .A2(G953), .ZN(n723) );
  XOR2_X1 U769 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n719) );
  NAND2_X1 U770 ( .A1(G224), .A2(G953), .ZN(n718) );
  XNOR2_X1 U771 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U772 ( .A(KEYINPUT124), .B(n720), .ZN(n721) );
  NAND2_X1 U773 ( .A1(G898), .A2(n721), .ZN(n722) );
  NAND2_X1 U774 ( .A1(n723), .A2(n722), .ZN(n730) );
  XNOR2_X1 U775 ( .A(n724), .B(G101), .ZN(n726) );
  XNOR2_X1 U776 ( .A(n726), .B(n725), .ZN(n727) );
  NAND2_X1 U777 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U778 ( .A(n730), .B(n729), .Z(G69) );
  XOR2_X1 U779 ( .A(n732), .B(n731), .Z(n735) );
  XOR2_X1 U780 ( .A(n735), .B(n733), .Z(n734) );
  NAND2_X1 U781 ( .A1(n734), .A2(n470), .ZN(n739) );
  XNOR2_X1 U782 ( .A(G227), .B(n735), .ZN(n736) );
  NAND2_X1 U783 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n737), .A2(G953), .ZN(n738) );
  NAND2_X1 U785 ( .A1(n739), .A2(n738), .ZN(G72) );
  XNOR2_X1 U786 ( .A(G119), .B(KEYINPUT127), .ZN(n741) );
  XNOR2_X1 U787 ( .A(n741), .B(n740), .ZN(G21) );
  XNOR2_X1 U788 ( .A(n742), .B(G131), .ZN(G33) );
  XNOR2_X1 U789 ( .A(n743), .B(G101), .ZN(G3) );
endmodule

