//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G50), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(KEYINPUT65), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n207), .B1(new_n208), .B2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G13), .ZN(new_n210));
  NAND4_X1  g0010(.A1(new_n210), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G116), .A2(G270), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G50), .A2(G226), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT67), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  AOI211_X1 g0021(.A(new_n220), .B(new_n221), .C1(G107), .C2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G97), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G87), .ZN(new_n228));
  INV_X1    g0028(.A(G250), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n208), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g0035(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n237));
  NAND3_X1  g0037(.A1(new_n236), .A2(G50), .A3(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(new_n239));
  AOI211_X1 g0039(.A(new_n214), .B(new_n232), .C1(new_n235), .C2(new_n239), .ZN(G361));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT68), .B(G264), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G358));
  XNOR2_X1  g0049(.A(G68), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT69), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n203), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(new_n223), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  NOR2_X1   g0057(.A1(new_n210), .A2(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n203), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n233), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(G20), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n260), .B1(new_n264), .B2(new_n203), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT73), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n261), .A2(new_n233), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n223), .A2(KEYINPUT8), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT71), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT8), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G58), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT72), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT71), .B1(new_n273), .B2(new_n223), .ZN(new_n274));
  OAI221_X1 g0074(.A(new_n270), .B1(new_n272), .B2(new_n273), .C1(new_n274), .C2(new_n271), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n234), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n275), .A2(new_n277), .B1(G150), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n204), .A2(G20), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n267), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n266), .A2(new_n281), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n282), .A2(KEYINPUT9), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n233), .ZN(new_n290));
  NAND3_X1  g0090(.A1(KEYINPUT70), .A2(G33), .A3(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n284), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n286), .B1(new_n294), .B2(G226), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n290), .A2(new_n287), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT3), .B(G33), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G222), .ZN(new_n299));
  INV_X1    g0099(.A(G223), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n297), .B(new_n299), .C1(new_n300), .C2(new_n298), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(G77), .B2(new_n297), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n295), .B1(new_n296), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G200), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n282), .B2(KEYINPUT9), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n283), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(G179), .B2(new_n303), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(new_n282), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n268), .A2(new_n272), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(new_n278), .B1(G20), .B2(G77), .ZN(new_n320));
  XOR2_X1   g0120(.A(KEYINPUT15), .B(G87), .Z(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n320), .B1(new_n276), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G77), .ZN(new_n324));
  INV_X1    g0124(.A(new_n259), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n323), .A2(new_n262), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n264), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n326), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n286), .ZN(new_n329));
  INV_X1    g0129(.A(G244), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n293), .B2(new_n330), .ZN(new_n331));
  XOR2_X1   g0131(.A(new_n331), .B(KEYINPUT74), .Z(new_n332));
  NAND2_X1  g0132(.A1(G238), .A2(G1698), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n297), .B(new_n333), .C1(new_n224), .C2(G1698), .ZN(new_n334));
  INV_X1    g0134(.A(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT3), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G33), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G107), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n296), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n332), .B1(new_n334), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n328), .B1(new_n342), .B2(G190), .ZN(new_n343));
  INV_X1    g0143(.A(G200), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n344), .B2(new_n342), .ZN(new_n345));
  INV_X1    g0145(.A(G179), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n328), .C1(G169), .C2(new_n342), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n317), .B1(KEYINPUT75), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n296), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n297), .A2(G232), .A3(G1698), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT76), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT76), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n297), .A2(new_n355), .A3(G232), .A4(G1698), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n297), .A2(G226), .A3(new_n298), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n352), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT77), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n286), .B1(new_n294), .B2(G238), .ZN(new_n364));
  OAI211_X1 g0164(.A(KEYINPUT77), .B(new_n352), .C1(new_n357), .C2(new_n360), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT13), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n363), .A2(KEYINPUT13), .A3(new_n364), .A4(new_n365), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(G169), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT14), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n366), .A2(new_n372), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(G179), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT14), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n368), .A2(new_n376), .A3(G169), .A4(new_n369), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n371), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n277), .A2(G77), .ZN(new_n379));
  INV_X1    g0179(.A(G68), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n278), .A2(G50), .B1(G20), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n267), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT11), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n327), .A2(new_n380), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n258), .A2(G20), .A3(new_n380), .ZN(new_n385));
  XOR2_X1   g0185(.A(new_n385), .B(KEYINPUT12), .Z(new_n386));
  NOR3_X1   g0186(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n378), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT75), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(new_n349), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT7), .B1(new_n339), .B2(new_n234), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  AOI211_X1 g0194(.A(new_n394), .B(G20), .C1(new_n336), .C2(new_n338), .ZN(new_n395));
  OAI21_X1  g0195(.A(G68), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n223), .A2(new_n380), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n202), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n278), .A2(G159), .ZN(new_n399));
  XOR2_X1   g0199(.A(new_n399), .B(KEYINPUT79), .Z(new_n400));
  NAND3_X1  g0200(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n398), .A4(new_n400), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n262), .A3(new_n404), .ZN(new_n405));
  OR2_X1    g0205(.A1(new_n275), .A2(new_n259), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n275), .A2(new_n264), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n294), .A2(G232), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n329), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n300), .A2(new_n298), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n297), .B(new_n411), .C1(G226), .C2(new_n298), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n296), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n344), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(G190), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n408), .A2(KEYINPUT17), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT17), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n405), .A2(new_n418), .A3(new_n406), .A4(new_n407), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n416), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n412), .A2(new_n413), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n329), .B(new_n409), .C1(new_n424), .C2(new_n296), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(G179), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n312), .B2(new_n425), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n423), .A2(new_n427), .A3(KEYINPUT18), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT18), .B1(new_n423), .B2(new_n427), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n419), .B(new_n422), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n373), .A2(G190), .A3(new_n374), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n368), .A2(G200), .A3(new_n369), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n387), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n351), .A2(new_n392), .A3(new_n431), .A4(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n297), .A2(new_n234), .A3(G87), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT22), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT22), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n297), .A2(new_n438), .A3(new_n234), .A4(G87), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n340), .A2(G20), .ZN(new_n441));
  XOR2_X1   g0241(.A(new_n441), .B(KEYINPUT23), .Z(new_n442));
  NAND3_X1  g0242(.A1(new_n234), .A2(G33), .A3(G116), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT24), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n440), .A2(KEYINPUT24), .A3(new_n442), .A4(new_n443), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n262), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n263), .A2(G33), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n267), .A2(new_n259), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G107), .ZN(new_n451));
  INV_X1    g0251(.A(new_n258), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(new_n441), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT25), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n448), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G1), .ZN(new_n457));
  AND2_X1   g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  NOR2_X1   g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n292), .A2(new_n460), .A3(G264), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT87), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n292), .A2(new_n460), .A3(KEYINPUT87), .A4(G264), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n229), .A2(new_n298), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n226), .A2(G1698), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n297), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G294), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n352), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n457), .B(G274), .C1(new_n459), .C2(new_n458), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n465), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT88), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n463), .A2(new_n464), .B1(new_n352), .B2(new_n470), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT88), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n472), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n474), .A2(G169), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n473), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G179), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n478), .A2(KEYINPUT89), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT89), .B1(new_n478), .B2(new_n480), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n455), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT90), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(KEYINPUT90), .B(new_n455), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n474), .A2(new_n477), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n305), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n473), .A2(new_n344), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n455), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n278), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT80), .B1(new_n494), .B2(new_n324), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT80), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n278), .A2(new_n496), .A3(G77), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n340), .A2(KEYINPUT6), .A3(G97), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  XNOR2_X1  g0300(.A(G97), .B(G107), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n495), .B(new_n497), .C1(new_n502), .C2(new_n234), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT81), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(G107), .B1(new_n393), .B2(new_n395), .ZN(new_n506));
  AND2_X1   g0306(.A1(G97), .A2(G107), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n500), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n498), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G20), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n511), .A2(KEYINPUT81), .A3(new_n495), .A4(new_n497), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n505), .A2(new_n506), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n262), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n325), .A2(new_n225), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n450), .A2(G97), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n297), .A2(KEYINPUT4), .A3(G244), .A4(new_n298), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n336), .A2(new_n338), .A3(G244), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT4), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n518), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n297), .A2(G250), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n298), .B1(new_n524), .B2(KEYINPUT4), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n352), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n292), .A2(new_n460), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G257), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n472), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT83), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT83), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n526), .A2(new_n531), .A3(new_n472), .A4(new_n528), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n312), .A3(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n519), .A2(new_n520), .B1(G33), .B2(G283), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n520), .B1(new_n297), .B2(G250), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n534), .B(new_n518), .C1(new_n298), .C2(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(new_n352), .B1(G257), .B2(new_n527), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(new_n346), .A3(new_n472), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n517), .A2(new_n533), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n305), .B1(new_n530), .B2(new_n532), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n540), .B(KEYINPUT84), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n529), .A2(G200), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n517), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n513), .A2(new_n262), .B1(new_n225), .B2(new_n325), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(KEYINPUT82), .A3(new_n516), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n539), .B1(new_n541), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G116), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n325), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n267), .A2(new_n259), .A3(new_n449), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n522), .B(new_n234), .C1(G33), .C2(new_n225), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n553), .B(new_n262), .C1(new_n234), .C2(G116), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT20), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  OAI221_X1 g0357(.A(new_n551), .B1(new_n550), .B2(new_n552), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G264), .A2(G1698), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n297), .B(new_n559), .C1(new_n226), .C2(G1698), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n560), .B(new_n352), .C1(G303), .C2(new_n297), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n527), .A2(G270), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n472), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n558), .A2(G169), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT86), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT21), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n565), .B1(new_n564), .B2(new_n566), .ZN(new_n568));
  INV_X1    g0368(.A(new_n558), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n561), .A2(new_n562), .A3(new_n472), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G179), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n563), .A2(KEYINPUT21), .A3(G169), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n567), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n563), .A2(G200), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n569), .B(new_n575), .C1(new_n305), .C2(new_n563), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(G238), .A2(G1698), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n330), .B2(G1698), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n580), .A2(new_n297), .B1(G33), .B2(G116), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n581), .A2(new_n296), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n263), .A2(G45), .A3(G274), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n457), .B2(new_n229), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n292), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(G200), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n508), .A2(new_n228), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n359), .A2(new_n234), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(KEYINPUT19), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n336), .A2(new_n338), .A3(new_n234), .A4(G68), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT19), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n359), .B2(G20), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(new_n262), .B1(new_n325), .B2(new_n322), .ZN(new_n596));
  OAI211_X1 g0396(.A(G190), .B(new_n585), .C1(new_n581), .C2(new_n296), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n450), .A2(G87), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n588), .A2(new_n599), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n581), .A2(new_n296), .ZN(new_n601));
  AOI21_X1  g0401(.A(G169), .B1(new_n601), .B2(new_n585), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n595), .A2(new_n262), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n450), .A2(new_n321), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n322), .A2(new_n325), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT85), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n596), .A2(KEYINPUT85), .A3(new_n604), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n602), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n582), .A2(new_n586), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n346), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n600), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n549), .A2(new_n578), .A3(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n435), .A2(new_n493), .A3(new_n614), .ZN(G372));
  INV_X1    g0415(.A(new_n435), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n587), .B(KEYINPUT91), .ZN(new_n617));
  INV_X1    g0417(.A(new_n599), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n610), .A2(new_n612), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n478), .A2(new_n480), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n455), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n574), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n549), .A2(new_n492), .A3(new_n621), .A4(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(KEYINPUT82), .A2(new_n514), .A3(new_n515), .A4(new_n516), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT82), .B1(new_n546), .B2(new_n516), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n533), .A2(new_n538), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .A4(new_n621), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT92), .ZN(new_n632));
  INV_X1    g0432(.A(new_n620), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n613), .A2(new_n533), .A3(new_n538), .A4(new_n517), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n633), .B1(new_n634), .B2(KEYINPUT26), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n631), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n632), .B1(new_n631), .B2(new_n635), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n625), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n616), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n428), .A2(new_n429), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n348), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n390), .B1(new_n642), .B2(new_n434), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n419), .A2(new_n422), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n315), .B1(new_n645), .B2(new_n311), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n639), .A2(new_n646), .ZN(G369));
  OR3_X1    g0447(.A1(new_n452), .A2(KEYINPUT27), .A3(G20), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT27), .B1(new_n452), .B2(G20), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n493), .B1(new_n455), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n483), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(new_n652), .ZN(new_n655));
  INV_X1    g0455(.A(new_n652), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n569), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n577), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n574), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n657), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n493), .A2(new_n623), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n624), .A3(new_n656), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(G399));
  INV_X1    g0467(.A(new_n212), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n508), .A2(new_n228), .A3(new_n550), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(G1), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n238), .B2(new_n670), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT28), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n638), .A2(new_n656), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n634), .A2(new_n629), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT95), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n628), .A2(KEYINPUT26), .A3(new_n630), .A4(new_n621), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n634), .A2(KEYINPUT95), .A3(new_n629), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n539), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n542), .B1(new_n626), .B2(new_n627), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n531), .B1(new_n537), .B2(new_n472), .ZN(new_n686));
  INV_X1    g0486(.A(new_n532), .ZN(new_n687));
  OAI21_X1  g0487(.A(G190), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT84), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT84), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n540), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n492), .B(new_n684), .C1(new_n685), .C2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(new_n487), .B2(new_n574), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n683), .B1(new_n694), .B2(new_n619), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n652), .B1(new_n695), .B2(new_n620), .ZN(new_n696));
  MUX2_X1   g0496(.A(new_n676), .B(new_n696), .S(KEYINPUT29), .Z(new_n697));
  NOR2_X1   g0497(.A1(new_n479), .A2(new_n570), .ZN(new_n698));
  INV_X1    g0498(.A(new_n611), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n698), .A2(new_n346), .A3(new_n699), .A4(new_n529), .ZN(new_n700));
  INV_X1    g0500(.A(new_n571), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n475), .A2(new_n611), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n701), .B(new_n702), .C1(new_n686), .C2(new_n687), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(KEYINPUT30), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n571), .B1(new_n530), .B2(new_n532), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n706), .B2(new_n702), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n700), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT93), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n613), .B(new_n684), .C1(new_n685), .C2(new_n692), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n577), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n491), .B1(new_n485), .B2(new_n486), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n712), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n708), .A2(KEYINPUT94), .ZN(new_n717));
  INV_X1    g0517(.A(new_n700), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n703), .A2(KEYINPUT30), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n706), .A2(new_n705), .A3(new_n702), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT94), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n656), .B1(new_n724), .B2(new_n712), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n711), .B1(new_n716), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n697), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n675), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n210), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n263), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n669), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n661), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT97), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n734), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n312), .A2(KEYINPUT98), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n234), .B1(KEYINPUT98), .B2(new_n312), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n233), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n234), .A2(new_n305), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n344), .A2(G179), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G303), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n234), .A2(G190), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G283), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n346), .A2(new_n344), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n749), .ZN(new_n754));
  INV_X1    g0554(.A(G317), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n749), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n752), .B(new_n758), .C1(G329), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n346), .A2(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n749), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G311), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n234), .B1(new_n759), .B2(G190), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G294), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n744), .A2(new_n753), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n297), .B1(new_n772), .B2(G326), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n762), .A2(new_n767), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n744), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n764), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n748), .B(new_n774), .C1(G322), .C2(new_n776), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n769), .A2(KEYINPUT99), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n769), .A2(KEYINPUT99), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G97), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n766), .A2(G77), .B1(new_n772), .B2(G50), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n760), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT32), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n785), .A2(new_n786), .B1(new_n380), .B2(new_n754), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n786), .B2(new_n785), .ZN(new_n788));
  INV_X1    g0588(.A(new_n746), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G87), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n782), .A2(new_n783), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n750), .A2(new_n340), .ZN(new_n792));
  INV_X1    g0592(.A(new_n776), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n223), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n791), .A2(new_n339), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n743), .B1(new_n777), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n253), .A2(G45), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n668), .A2(new_n297), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n797), .B(new_n798), .C1(G45), .C2(new_n238), .ZN(new_n799));
  INV_X1    g0599(.A(G355), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n212), .A2(new_n297), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT96), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n799), .B1(G116), .B2(new_n212), .C1(new_n800), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n738), .A2(new_n743), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n739), .A2(new_n796), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G330), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n735), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n808), .A2(new_n662), .A3(new_n734), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT100), .ZN(G396));
  NAND2_X1  g0611(.A1(new_n328), .A2(new_n652), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n345), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n348), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n642), .A2(new_n656), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n676), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n816), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n638), .A2(new_n656), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n717), .A2(new_n723), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n652), .B1(new_n821), .B2(KEYINPUT31), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT31), .B1(new_n493), .B2(new_n614), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n807), .B1(new_n824), .B2(new_n711), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n820), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n734), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n782), .B1(new_n751), .B2(new_n754), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n750), .A2(new_n228), .B1(new_n760), .B2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT102), .Z(new_n831));
  INV_X1    g0631(.A(new_n766), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n832), .A2(new_n550), .B1(new_n747), .B2(new_n771), .ZN(new_n833));
  NOR4_X1   g0633(.A1(new_n828), .A2(new_n297), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G294), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n340), .B2(new_n746), .C1(new_n835), .C2(new_n793), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n766), .A2(G159), .B1(new_n776), .B2(G143), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  INV_X1    g0638(.A(G150), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n838), .B2(new_n771), .C1(new_n839), .C2(new_n754), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT34), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n339), .B1(new_n761), .B2(G132), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n746), .A2(new_n203), .B1(new_n750), .B2(new_n380), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G58), .B2(new_n769), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n836), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT103), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n734), .B1(new_n847), .B2(new_n743), .ZN(new_n848));
  INV_X1    g0648(.A(new_n737), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(new_n743), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT101), .Z(new_n851));
  OAI221_X1 g0651(.A(new_n848), .B1(G77), .B2(new_n851), .C1(new_n818), .C2(new_n737), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT104), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n827), .A2(new_n853), .ZN(G384));
  OR2_X1    g0654(.A1(new_n697), .A2(new_n435), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n646), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT108), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n821), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n716), .B2(new_n725), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n388), .A2(new_n652), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n434), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT105), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n378), .A2(new_n863), .A3(new_n388), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(new_n378), .B2(new_n388), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n389), .A2(new_n656), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n816), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n859), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT40), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT106), .ZN(new_n872));
  INV_X1    g0672(.A(new_n650), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n423), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n872), .B1(new_n423), .B2(new_n873), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n430), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n423), .A2(new_n873), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT106), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n874), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n423), .A2(new_n427), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n421), .A2(new_n416), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n879), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n423), .A2(new_n427), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n887), .B(new_n880), .C1(new_n416), .C2(new_n421), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n878), .B(KEYINPUT38), .C1(new_n886), .C2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT107), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n887), .B1(new_n416), .B2(new_n421), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT37), .B1(new_n877), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n885), .A2(new_n879), .A3(new_n880), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n896), .A2(KEYINPUT107), .A3(KEYINPUT38), .A4(new_n878), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n431), .A2(new_n880), .B1(new_n899), .B2(new_n889), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n871), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n878), .B1(new_n886), .B2(new_n889), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n901), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n890), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n859), .A2(new_n906), .A3(new_n869), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n870), .A2(new_n903), .B1(new_n907), .B2(new_n871), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n616), .A2(new_n859), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(G330), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n857), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n898), .A2(new_n902), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n864), .A2(new_n865), .A3(new_n652), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n890), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n866), .A2(new_n868), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n819), .B2(new_n815), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n906), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n641), .A2(new_n873), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n918), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n912), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n263), .B2(new_n730), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n550), .B1(new_n510), .B2(KEYINPUT35), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n927), .B(new_n235), .C1(KEYINPUT35), .C2(new_n510), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT36), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n238), .A2(new_n324), .A3(new_n397), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n380), .A2(G50), .ZN(new_n931));
  OAI211_X1 g0731(.A(G1), .B(new_n210), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n926), .A2(new_n929), .A3(new_n932), .ZN(G367));
  NAND2_X1  g0733(.A1(new_n628), .A2(new_n652), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n549), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n628), .A2(new_n630), .A3(new_n652), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n664), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n574), .A2(new_n652), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n653), .A2(new_n549), .A3(new_n934), .A4(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT42), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n684), .B1(new_n938), .B2(new_n487), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n656), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT109), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n596), .A2(new_n598), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n652), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n621), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n620), .A2(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n948), .A2(new_n949), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n954), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n943), .A2(new_n944), .B1(new_n656), .B2(new_n946), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n956), .B1(new_n957), .B2(KEYINPUT109), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n955), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT43), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n955), .B2(new_n958), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n939), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n939), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n955), .A2(new_n958), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n965), .B(new_n960), .C1(new_n966), .C2(new_n962), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n669), .B(KEYINPUT41), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n655), .B(new_n662), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(new_n940), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n666), .A2(new_n937), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT45), .Z(new_n973));
  NOR2_X1   g0773(.A1(new_n666), .A2(new_n549), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n663), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n973), .A2(new_n664), .A3(new_n975), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n971), .A2(new_n977), .A3(new_n728), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n969), .B1(new_n979), .B2(new_n728), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n964), .B(new_n967), .C1(new_n980), .C2(new_n732), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n297), .B1(new_n750), .B2(new_n324), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n746), .A2(new_n223), .B1(new_n760), .B2(new_n838), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT111), .ZN(new_n984));
  INV_X1    g0784(.A(new_n754), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G143), .A2(new_n772), .B1(new_n985), .B2(G159), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n984), .B(new_n986), .C1(new_n380), .C2(new_n780), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n982), .B(new_n987), .C1(G150), .C2(new_n776), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n766), .A2(G50), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n761), .A2(G317), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n793), .A2(new_n747), .B1(new_n829), .B2(new_n771), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT110), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n746), .A2(new_n550), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n993), .A2(KEYINPUT46), .B1(G107), .B2(new_n769), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n994), .B(new_n339), .C1(new_n835), .C2(new_n754), .ZN(new_n995));
  INV_X1    g0795(.A(new_n750), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(G97), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n993), .B2(KEYINPUT46), .C1(new_n832), .C2(new_n751), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n992), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n988), .A2(new_n989), .B1(new_n990), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT47), .Z(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n743), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n956), .A2(new_n738), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n798), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n804), .B1(new_n212), .B2(new_n322), .C1(new_n248), .C2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n733), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n981), .A2(new_n1006), .ZN(G387));
  OR2_X1    g0807(.A1(new_n971), .A2(new_n728), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n971), .A2(new_n728), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n669), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n655), .A2(new_n738), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n318), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(new_n671), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(G68), .A2(G77), .ZN(new_n1014));
  OAI21_X1  g0814(.A(KEYINPUT50), .B1(new_n318), .B2(G50), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1013), .A2(new_n456), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n798), .B(new_n1016), .C1(new_n244), .C2(new_n456), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(G107), .B2(new_n212), .C1(new_n672), .C2(new_n802), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n734), .B1(new_n1018), .B2(new_n804), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1011), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n339), .B1(new_n275), .B2(new_n985), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n324), .B2(new_n746), .C1(new_n784), .C2(new_n771), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n781), .A2(new_n321), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n839), .B2(new_n760), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1022), .B(new_n1024), .C1(G50), .C2(new_n776), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1025), .B(new_n997), .C1(new_n380), .C2(new_n832), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT112), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n766), .A2(G303), .B1(new_n776), .B2(G317), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT113), .Z(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n829), .B2(new_n754), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G322), .B2(new_n772), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT48), .Z(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n751), .B2(new_n768), .C1(new_n835), .C2(new_n746), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT49), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n996), .A2(G116), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n761), .A2(G326), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1035), .A2(new_n339), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1027), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1020), .B1(new_n1040), .B2(new_n743), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n971), .B2(new_n732), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1010), .A2(new_n1042), .ZN(G393));
  NAND3_X1  g0843(.A1(new_n977), .A2(new_n732), .A3(new_n978), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n938), .A2(new_n738), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n776), .A2(G311), .B1(new_n772), .B2(G317), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT52), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n832), .A2(new_n835), .B1(new_n768), .B2(new_n550), .ZN(new_n1048));
  INV_X1    g0848(.A(G322), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n339), .B1(new_n760), .B2(new_n1049), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1047), .A2(new_n792), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n751), .B2(new_n746), .C1(new_n747), .C2(new_n754), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n339), .B1(new_n761), .B2(G143), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n380), .B2(new_n746), .C1(new_n228), .C2(new_n750), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT114), .Z(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n319), .B2(new_n766), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n780), .A2(new_n324), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1056), .B(new_n1058), .C1(new_n203), .C2(new_n754), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n776), .A2(G159), .B1(new_n772), .B2(G150), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT51), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1052), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n743), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n798), .A2(new_n256), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1064), .B(new_n804), .C1(new_n225), .C2(new_n212), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1045), .A2(new_n733), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1044), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n977), .A2(new_n978), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n670), .B1(new_n1009), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1067), .B1(new_n1069), .B2(new_n979), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(G390));
  INV_X1    g0871(.A(KEYINPUT115), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n866), .A2(new_n868), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n825), .A2(new_n1072), .A3(new_n818), .A4(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n726), .A2(G330), .A3(new_n818), .A4(new_n1073), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(KEYINPUT115), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n807), .B1(new_n824), .B2(new_n858), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n818), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1074), .A2(new_n1076), .B1(new_n1078), .B2(new_n919), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n815), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n696), .B2(new_n814), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n819), .A2(new_n815), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n919), .B1(new_n727), .B2(new_n816), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1077), .A2(new_n869), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1079), .A2(new_n1081), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n616), .A2(G330), .A3(new_n859), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n646), .B(new_n1087), .C1(new_n697), .C2(new_n435), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n916), .B1(new_n898), .B2(new_n902), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1081), .B2(new_n919), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT39), .B1(new_n898), .B2(new_n902), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n917), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n920), .A2(new_n916), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1091), .A2(new_n1074), .A3(new_n1076), .A4(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1093), .B1(new_n913), .B2(new_n914), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n916), .B1(new_n1082), .B2(new_n1073), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT89), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n622), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n478), .A2(KEYINPUT89), .A3(new_n480), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT90), .B1(new_n1101), .B2(new_n455), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n486), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n574), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n693), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n619), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(new_n620), .A3(new_n682), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1107), .A2(new_n656), .A3(new_n814), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n919), .B1(new_n1108), .B2(new_n815), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n916), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n913), .A2(new_n1110), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1096), .A2(new_n1097), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n1084), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1095), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1089), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1078), .A2(new_n919), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1081), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1085), .A2(new_n1082), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1088), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1095), .A2(new_n1113), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1115), .A2(new_n669), .A3(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1096), .A2(new_n737), .ZN(new_n1126));
  INV_X1    g0926(.A(G125), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n297), .B1(new_n760), .B2(new_n1127), .C1(new_n838), .C2(new_n754), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n789), .A2(G150), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1129), .A2(KEYINPUT53), .B1(new_n996), .B2(G50), .ZN(new_n1130));
  INV_X1    g0930(.A(G132), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1130), .B1(KEYINPUT53), .B2(new_n1129), .C1(new_n1131), .C2(new_n793), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT54), .B(G143), .Z(new_n1133));
  AOI211_X1 g0933(.A(new_n1128), .B(new_n1132), .C1(new_n766), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(G128), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n771), .C1(new_n784), .C2(new_n780), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT116), .Z(new_n1137));
  OAI22_X1  g0937(.A1(new_n832), .A2(new_n225), .B1(new_n751), .B2(new_n771), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G107), .B2(new_n985), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT117), .Z(new_n1140));
  NAND2_X1  g0940(.A1(new_n790), .A2(new_n339), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1141), .A2(KEYINPUT118), .B1(G68), .B2(new_n996), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(new_n835), .C2(new_n760), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1058), .B1(KEYINPUT118), .B2(new_n1141), .C1(new_n550), .C2(new_n793), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n743), .B1(new_n1137), .B2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1146), .B(new_n733), .C1(new_n275), .C2(new_n851), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1126), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n1114), .B2(new_n732), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT119), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1125), .B1(new_n1151), .B2(new_n1152), .ZN(G378));
  NAND2_X1  g0953(.A1(new_n317), .A2(KEYINPUT123), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT123), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n311), .A2(new_n1155), .A3(new_n316), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n282), .A2(new_n650), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1154), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1155), .B1(new_n311), .B2(new_n316), .ZN(new_n1160));
  AOI211_X1 g0960(.A(KEYINPUT123), .B(new_n315), .C1(new_n309), .C2(new_n310), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1157), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1159), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n908), .B2(G330), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n913), .A2(KEYINPUT40), .A3(new_n859), .A4(new_n869), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n907), .A2(new_n871), .ZN(new_n1169));
  AND4_X1   g0969(.A1(G330), .A2(new_n1168), .A3(new_n1169), .A4(new_n1166), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n924), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1168), .A2(new_n1169), .A3(G330), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1166), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n918), .A2(new_n921), .A3(new_n923), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1168), .A2(new_n1169), .A3(new_n1166), .A4(G330), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT124), .B1(new_n1171), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1175), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT124), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n732), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1166), .A2(new_n849), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n780), .A2(new_n380), .B1(new_n340), .B2(new_n793), .ZN(new_n1184));
  AOI211_X1 g0984(.A(G41), .B(new_n297), .C1(new_n761), .C2(G283), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n223), .B2(new_n750), .C1(new_n324), .C2(new_n746), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT121), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1184), .B(new_n1187), .C1(G97), .C2(new_n985), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n550), .B2(new_n771), .C1(new_n322), .C2(new_n832), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT58), .Z(new_n1190));
  NOR2_X1   g0990(.A1(G33), .A2(G41), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT120), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n203), .C1(G41), .C2(new_n297), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n771), .A2(new_n1127), .B1(new_n754), .B2(new_n1131), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n780), .A2(new_n839), .B1(new_n838), .B2(new_n832), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(new_n789), .C2(new_n1133), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n1135), .B2(new_n793), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT59), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(KEYINPUT122), .A2(G124), .ZN(new_n1199));
  AND2_X1   g0999(.A1(KEYINPUT122), .A2(G124), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n761), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n996), .A2(G159), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1192), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1193), .B1(new_n1198), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n743), .B1(new_n1190), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n850), .A2(new_n203), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1183), .A2(new_n733), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1182), .A2(KEYINPUT125), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT125), .B1(new_n1182), .B2(new_n1208), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1121), .B1(new_n1123), .B2(new_n1086), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1171), .A2(new_n1177), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(KEYINPUT57), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1088), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1180), .B1(new_n1216), .B2(new_n1179), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1171), .A2(KEYINPUT124), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1215), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n669), .B(new_n1214), .C1(new_n1219), .C2(KEYINPUT57), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1211), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(G375));
  OAI221_X1 g1022(.A(new_n297), .B1(new_n1131), .B2(new_n771), .C1(new_n793), .C2(new_n838), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G159), .B2(new_n789), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n766), .A2(G150), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n781), .A2(G50), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G58), .A2(new_n996), .B1(new_n761), .B2(G128), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n985), .B2(new_n1133), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n985), .A2(G116), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n761), .A2(G303), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n297), .B1(new_n776), .B2(G283), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1023), .A2(new_n1230), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n832), .A2(new_n340), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n746), .A2(new_n225), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n771), .A2(new_n835), .B1(new_n750), .B2(new_n324), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n743), .B1(new_n1229), .B2(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1238), .B(new_n733), .C1(G68), .C2(new_n851), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n919), .B2(new_n849), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n1120), .B2(new_n732), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1118), .A2(new_n1088), .A3(new_n1119), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n968), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1241), .B1(new_n1243), .B2(new_n1089), .ZN(G381));
  NAND2_X1  g1044(.A1(new_n1125), .A2(new_n1149), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n981), .A2(new_n1006), .A3(new_n1070), .ZN(new_n1247));
  OR2_X1    g1047(.A1(G381), .A2(G384), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1247), .A2(G396), .A3(G393), .A4(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1221), .A2(new_n1246), .A3(new_n1249), .ZN(G407));
  OAI211_X1 g1050(.A(new_n1221), .B(new_n1246), .C1(new_n1249), .C2(new_n651), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(G213), .ZN(G409));
  INV_X1    g1052(.A(KEYINPUT62), .ZN(new_n1253));
  INV_X1    g1053(.A(G213), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(G343), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1086), .A2(KEYINPUT60), .A3(new_n1088), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT60), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1242), .A2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1256), .A2(new_n1258), .A3(new_n669), .A4(new_n1122), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G384), .B1(new_n1259), .B2(new_n1241), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(G384), .A3(new_n1241), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1220), .B(G378), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1213), .A2(new_n732), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1212), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1208), .B(new_n1265), .C1(new_n1266), .C2(new_n969), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1246), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1255), .B(new_n1263), .C1(new_n1264), .C2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1253), .B1(new_n1269), .B2(KEYINPUT127), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1264), .A2(new_n1268), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1255), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1262), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G2897), .B(new_n1255), .C1(new_n1274), .C2(new_n1260), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1255), .A2(G2897), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1261), .A2(new_n1262), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT61), .B1(new_n1273), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1263), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1271), .A2(new_n1272), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n1283), .A3(KEYINPUT62), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1270), .A2(new_n1280), .A3(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G387), .A2(G390), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(new_n1287), .B2(new_n1247), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(G393), .B(G396), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1247), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT126), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1287), .A2(new_n1286), .A3(new_n1247), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1290), .B1(new_n1294), .B2(new_n1289), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1285), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1278), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1282), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  OR2_X1    g1099(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1247), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1070), .B1(new_n981), .B2(new_n1006), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1301), .A2(KEYINPUT126), .A3(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1289), .B1(new_n1303), .B2(new_n1288), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT61), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1269), .A2(KEYINPUT63), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1299), .A2(new_n1305), .A3(new_n1306), .A4(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1296), .A2(new_n1308), .ZN(G405));
  OAI211_X1 g1109(.A(new_n1264), .B(new_n1263), .C1(new_n1221), .C2(new_n1245), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1245), .B1(new_n1211), .B2(new_n1220), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1264), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1281), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1314), .B(new_n1295), .ZN(G402));
endmodule


