//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  AOI21_X1  g002(.A(KEYINPUT23), .B1(new_n188), .B2(G119), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(G119), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n194), .A3(G119), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n191), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G110), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n199), .A2(KEYINPUT16), .A3(G140), .ZN(new_n200));
  XNOR2_X1  g014(.A(G125), .B(G140), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(KEYINPUT16), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  AOI211_X1 g018(.A(new_n204), .B(new_n200), .C1(KEYINPUT16), .C2(new_n201), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n198), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n190), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n195), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT70), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n195), .A2(new_n211), .A3(new_n208), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g027(.A(KEYINPUT24), .B(G110), .Z(new_n214));
  AOI21_X1  g028(.A(KEYINPUT71), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n195), .A2(new_n211), .A3(new_n208), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n211), .B1(new_n195), .B2(new_n208), .ZN(new_n217));
  OAI211_X1 g031(.A(KEYINPUT71), .B(new_n214), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n207), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  OR3_X1    g034(.A1(new_n216), .A2(new_n217), .A3(new_n214), .ZN(new_n221));
  OR2_X1    g035(.A1(new_n197), .A2(G110), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n202), .A2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n201), .A2(new_n204), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT22), .B(G137), .ZN(new_n229));
  INV_X1    g043(.A(G953), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n230), .A2(G221), .A3(G234), .ZN(new_n231));
  XOR2_X1   g045(.A(new_n229), .B(new_n231), .Z(new_n232));
  NAND3_X1  g046(.A1(new_n220), .A2(new_n228), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n232), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n206), .B1(new_n237), .B2(new_n218), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n226), .B1(new_n221), .B2(new_n222), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n234), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G902), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n233), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n233), .A2(new_n240), .A3(KEYINPUT25), .A4(new_n241), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n244), .A2(KEYINPUT72), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n242), .A2(new_n247), .A3(new_n243), .ZN(new_n248));
  INV_X1    g062(.A(G217), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(G234), .B2(new_n241), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n187), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n244), .A2(KEYINPUT72), .A3(new_n245), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n253), .A2(KEYINPUT73), .A3(new_n250), .A4(new_n248), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n233), .A2(new_n240), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n250), .A2(G902), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n252), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n252), .A2(KEYINPUT74), .A3(new_n254), .A4(new_n258), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n204), .A2(G143), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  OR2_X1    g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(G143), .B(G146), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT0), .A3(G128), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT11), .ZN(new_n274));
  INV_X1    g088(.A(G134), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(G137), .ZN(new_n276));
  INV_X1    g090(.A(G137), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT11), .A3(G134), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(G137), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G131), .ZN(new_n281));
  INV_X1    g095(.A(G131), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n276), .A2(new_n278), .A3(new_n282), .A4(new_n279), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n281), .A2(KEYINPUT67), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT67), .B1(new_n281), .B2(new_n283), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n273), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT64), .B(G128), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(G143), .B2(new_n204), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n267), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n271), .A2(new_n288), .A3(G128), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n279), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n275), .A2(G137), .ZN(new_n294));
  OAI21_X1  g108(.A(G131), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(new_n283), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n286), .A2(KEYINPUT30), .A3(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n281), .A2(new_n283), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n270), .A2(new_n272), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT30), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n303));
  INV_X1    g117(.A(G113), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT65), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT65), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT2), .A3(G113), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G116), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(G119), .ZN(new_n310));
  INV_X1    g124(.A(G119), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(G116), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n303), .A2(new_n304), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n308), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT66), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n310), .B2(new_n312), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n311), .A2(G116), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n309), .A2(G119), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT66), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n305), .A2(new_n307), .B1(new_n303), .B2(new_n304), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n297), .A2(new_n302), .A3(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(G237), .A2(G953), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G210), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT27), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT26), .B(G101), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n323), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n286), .A2(new_n330), .A3(new_n296), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n324), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT31), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n300), .A2(new_n323), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n286), .A2(new_n330), .A3(KEYINPUT28), .A4(new_n296), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n329), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT31), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n324), .A2(new_n341), .A3(new_n329), .A4(new_n331), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n333), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT68), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(G472), .A2(G902), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n333), .A2(new_n340), .A3(KEYINPUT68), .A4(new_n342), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT32), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT32), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n345), .A2(new_n350), .A3(new_n346), .A4(new_n347), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n335), .A2(new_n337), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n286), .A2(new_n296), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n323), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n339), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(G902), .B1(new_n357), .B2(KEYINPUT69), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n338), .A2(new_n329), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n324), .A2(new_n339), .A3(new_n331), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI221_X1 g175(.A(new_n358), .B1(KEYINPUT69), .B2(new_n357), .C1(new_n361), .C2(KEYINPUT29), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n349), .A2(new_n351), .B1(new_n362), .B2(G472), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n263), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G221), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT9), .B(G234), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n365), .B1(new_n367), .B2(new_n241), .ZN(new_n368));
  INV_X1    g182(.A(G469), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n284), .A2(new_n285), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n290), .A2(new_n291), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n372));
  INV_X1    g186(.A(G104), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT3), .B1(new_n373), .B2(G107), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n375));
  INV_X1    g189(.A(G107), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(G104), .ZN(new_n377));
  INV_X1    g191(.A(G101), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n373), .A2(G107), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n374), .A2(new_n377), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n373), .A2(G107), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n376), .A2(G104), .ZN(new_n382));
  OAI21_X1  g196(.A(G101), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n371), .A2(new_n372), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n374), .A2(new_n377), .A3(new_n379), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(G101), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n388), .A2(new_n272), .A3(new_n270), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(G101), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT4), .A3(new_n380), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT75), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n389), .A2(KEYINPUT75), .A3(new_n391), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n385), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT78), .ZN(new_n397));
  AND4_X1   g211(.A1(new_n288), .A2(new_n264), .A3(new_n266), .A4(G128), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT1), .B1(new_n265), .B2(G146), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT76), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT76), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n401), .B(KEYINPUT1), .C1(new_n265), .C2(G146), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(G128), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n398), .B1(new_n403), .B2(new_n267), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT77), .B1(new_n404), .B2(new_n384), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(G128), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n401), .B1(new_n264), .B2(KEYINPUT1), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n267), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n291), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT77), .ZN(new_n410));
  INV_X1    g224(.A(new_n384), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n405), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n397), .B1(new_n413), .B2(new_n372), .ZN(new_n414));
  AOI211_X1 g228(.A(KEYINPUT78), .B(KEYINPUT10), .C1(new_n405), .C2(new_n412), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n370), .B(new_n396), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G110), .B(G140), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n230), .A2(G227), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n417), .B(new_n418), .Z(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n416), .A2(KEYINPUT79), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT79), .B1(new_n416), .B2(new_n420), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT12), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n405), .A2(new_n412), .B1(new_n371), .B2(new_n384), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n423), .B1(new_n424), .B2(new_n370), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n404), .A2(KEYINPUT77), .A3(new_n384), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n410), .B1(new_n409), .B2(new_n411), .ZN(new_n427));
  OAI22_X1  g241(.A1(new_n426), .A2(new_n427), .B1(new_n292), .B2(new_n411), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n298), .A2(new_n423), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n421), .A2(new_n422), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n396), .B1(new_n414), .B2(new_n415), .ZN(new_n434));
  INV_X1    g248(.A(new_n370), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n420), .B1(new_n436), .B2(new_n416), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n369), .B(new_n241), .C1(new_n433), .C2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n369), .A2(new_n241), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n416), .A2(new_n431), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n419), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n436), .A2(new_n416), .A3(new_n420), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n439), .B1(new_n443), .B2(G469), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n368), .B1(new_n438), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G210), .B1(G237), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n371), .A2(new_n199), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n299), .A2(G125), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G224), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(G953), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n450), .B(new_n452), .Z(new_n453));
  NAND3_X1  g267(.A1(new_n323), .A2(new_n391), .A3(new_n388), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT5), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n317), .B2(new_n320), .ZN(new_n456));
  OAI21_X1  g270(.A(G113), .B1(new_n318), .B2(KEYINPUT5), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n411), .B(new_n315), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G110), .B(G122), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AND4_X1   g275(.A1(KEYINPUT81), .A2(new_n459), .A3(KEYINPUT6), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n454), .B2(new_n458), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT6), .B1(new_n463), .B2(KEYINPUT81), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n454), .A2(new_n458), .A3(new_n460), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT80), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n459), .A2(new_n461), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n454), .A2(new_n458), .A3(KEYINPUT80), .A4(new_n460), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n453), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT7), .B1(new_n451), .B2(G953), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n450), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n474), .ZN(new_n476));
  AOI211_X1 g290(.A(KEYINPUT82), .B(new_n476), .C1(new_n448), .C2(new_n449), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n315), .B(new_n384), .C1(new_n456), .C2(new_n457), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n460), .B(KEYINPUT8), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n457), .B1(new_n313), .B2(KEYINPUT5), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n322), .B2(new_n313), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n479), .B(new_n480), .C1(new_n482), .C2(new_n384), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n448), .A2(new_n449), .A3(new_n476), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n468), .A2(new_n470), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n241), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n447), .B1(new_n472), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n459), .A2(KEYINPUT81), .A3(new_n461), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n463), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n471), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n453), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n485), .A2(new_n475), .A3(new_n477), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n468), .A2(new_n470), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n446), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n490), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(G234), .A2(G237), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(G952), .A3(new_n230), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(G902), .A3(G953), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT21), .B(G898), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G214), .B1(G237), .B2(G902), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n502), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  NOR2_X1   g328(.A1(G475), .A2(G902), .ZN(new_n515));
  XNOR2_X1  g329(.A(G113), .B(G122), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(new_n373), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n325), .A2(G143), .A3(G214), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(G143), .B1(new_n325), .B2(G214), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(KEYINPUT18), .A2(G131), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(KEYINPUT18), .B(G131), .C1(new_n519), .C2(new_n520), .ZN(new_n524));
  INV_X1    g338(.A(G140), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G125), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n199), .A2(G140), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G146), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n225), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n523), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT16), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n204), .B1(new_n533), .B2(new_n200), .ZN(new_n534));
  OAI211_X1 g348(.A(KEYINPUT17), .B(G131), .C1(new_n519), .C2(new_n520), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n224), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G131), .B1(new_n519), .B2(new_n520), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n325), .A2(G214), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n265), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n282), .A3(new_n518), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n537), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n517), .B(new_n531), .C1(new_n536), .C2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n537), .A2(new_n540), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n201), .A2(KEYINPUT19), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n201), .A2(KEYINPUT19), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n545), .B(new_n224), .C1(G146), .C2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n517), .B1(new_n549), .B2(new_n531), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n514), .B(new_n515), .C1(new_n544), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT84), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n544), .A2(new_n550), .ZN(new_n555));
  INV_X1    g369(.A(new_n515), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n549), .A2(new_n531), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n543), .B1(new_n558), .B2(new_n517), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT84), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n514), .A4(new_n515), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n552), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n531), .B1(new_n536), .B2(new_n542), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(new_n517), .ZN(new_n564));
  OAI21_X1  g378(.A(G475), .B1(new_n564), .B2(G902), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT89), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n192), .A2(new_n194), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n571), .A2(KEYINPUT86), .A3(new_n265), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT86), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n287), .B2(G143), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT85), .B1(new_n188), .B2(G143), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT85), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n265), .A3(G128), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI22_X1  g392(.A1(new_n572), .A2(new_n574), .B1(KEYINPUT13), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n577), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT87), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT87), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n575), .A2(new_n577), .A3(new_n583), .A4(KEYINPUT13), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G134), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(G116), .B(G122), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G107), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT86), .B1(new_n571), .B2(new_n265), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n287), .A2(new_n573), .A3(G143), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n578), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n588), .B1(new_n591), .B2(new_n275), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n309), .A2(G122), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n376), .B1(new_n594), .B2(KEYINPUT14), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(new_n587), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n591), .A2(new_n275), .ZN(new_n597));
  AOI211_X1 g411(.A(G134), .B(new_n578), .C1(new_n589), .C2(new_n590), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n366), .A2(new_n249), .A3(G953), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n593), .A2(new_n599), .A3(new_n601), .ZN(new_n604));
  AOI21_X1  g418(.A(G902), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n570), .B1(new_n605), .B2(KEYINPUT88), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n593), .A2(new_n599), .A3(new_n601), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n601), .B1(new_n593), .B2(new_n599), .ZN(new_n608));
  OAI211_X1 g422(.A(KEYINPUT88), .B(new_n241), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n569), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n567), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n605), .A2(KEYINPUT88), .A3(new_n570), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n569), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n613), .A3(KEYINPUT89), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n513), .A2(new_n566), .A3(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n445), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n364), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  AND3_X1   g433(.A1(new_n445), .A2(new_n261), .A3(new_n262), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n345), .A2(new_n241), .A3(new_n347), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT90), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n345), .A2(KEYINPUT90), .A3(new_n241), .A4(new_n347), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(G472), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n348), .A2(KEYINPUT91), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT91), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n623), .A2(new_n628), .A3(G472), .A4(new_n624), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n620), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n497), .A2(new_n446), .A3(new_n500), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n511), .B1(new_n632), .B2(KEYINPUT92), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT92), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n490), .A2(new_n634), .A3(new_n501), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n568), .A2(new_n241), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n605), .B2(new_n568), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n603), .A2(new_n604), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n602), .B2(KEYINPUT93), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n603), .A2(new_n604), .A3(new_n642), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n568), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n566), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n636), .A2(new_n509), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n631), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT94), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT34), .B(G104), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  INV_X1    g467(.A(new_n615), .ZN(new_n654));
  INV_X1    g468(.A(new_n509), .ZN(new_n655));
  INV_X1    g469(.A(new_n557), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n555), .A2(new_n556), .A3(new_n554), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n565), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n636), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n631), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NAND2_X1  g476(.A1(new_n220), .A2(new_n228), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n234), .A2(KEYINPUT36), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n257), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT95), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n252), .A2(new_n254), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT96), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n252), .A2(KEYINPUT96), .A3(new_n668), .A4(new_n254), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n630), .A2(new_n617), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  INV_X1    g490(.A(new_n636), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n671), .A2(new_n677), .A3(new_n672), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n349), .A2(new_n351), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n362), .A2(G472), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n506), .A2(G900), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n504), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n565), .B(new_n683), .C1(new_n656), .C2(new_n657), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n615), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT97), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n678), .A2(new_n681), .A3(new_n445), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  AND3_X1   g503(.A1(new_n252), .A2(new_n254), .A3(new_n668), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n490), .A2(new_n501), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n691), .B1(new_n490), .B2(new_n501), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n511), .B1(new_n562), .B2(new_n565), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n615), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n690), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(G472), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n324), .A2(new_n331), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n329), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n331), .A2(new_n339), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(G902), .B1(new_n702), .B2(new_n354), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n698), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n349), .B2(new_n351), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT99), .B1(new_n697), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n691), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n446), .B1(new_n497), .B2(new_n500), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n707), .B1(new_n632), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n490), .A2(new_n501), .A3(new_n691), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n615), .A3(new_n695), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n669), .ZN(new_n712));
  INV_X1    g526(.A(new_n704), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n679), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT99), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT40), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n683), .B(KEYINPUT39), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n445), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n438), .A2(new_n444), .ZN(new_n720));
  INV_X1    g534(.A(new_n368), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n721), .A3(new_n718), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n706), .A2(new_n716), .A3(new_n719), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G143), .ZN(G45));
  INV_X1    g539(.A(new_n645), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n642), .B1(new_n603), .B2(new_n604), .ZN(new_n727));
  OAI21_X1  g541(.A(G478), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n566), .A2(new_n728), .A3(new_n638), .A4(new_n683), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n678), .A2(new_n681), .A3(new_n445), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G146), .ZN(G48));
  INV_X1    g546(.A(KEYINPUT101), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n416), .A2(new_n420), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT79), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n432), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n416), .A2(KEYINPUT79), .A3(new_n420), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n437), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(G469), .B1(new_n738), .B2(G902), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n438), .A3(new_n721), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT100), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT100), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n739), .A2(new_n438), .A3(new_n742), .A4(new_n721), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n681), .A2(new_n261), .A3(new_n262), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n733), .B1(new_n746), .B2(new_n649), .ZN(new_n747));
  INV_X1    g561(.A(new_n649), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n744), .A2(new_n745), .A3(new_n748), .A4(KEYINPUT101), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT41), .B(G113), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G15));
  NAND2_X1  g566(.A1(new_n746), .A2(new_n659), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G116), .ZN(G18));
  AND3_X1   g568(.A1(new_n739), .A2(new_n721), .A3(new_n438), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT102), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n756), .A3(new_n677), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT102), .B1(new_n740), .B2(new_n636), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n615), .A2(new_n566), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n681), .A2(new_n671), .A3(new_n672), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n759), .A2(new_n760), .A3(new_n655), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G119), .ZN(G21));
  AND2_X1   g577(.A1(new_n621), .A2(G472), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n352), .A2(new_n354), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n333), .B(new_n342), .C1(new_n765), .C2(new_n329), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n346), .B(KEYINPUT103), .Z(new_n767));
  AND2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n764), .A2(new_n259), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n633), .A2(new_n615), .A3(new_n566), .A4(new_n635), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n509), .ZN(new_n771));
  AND4_X1   g585(.A1(new_n741), .A2(new_n769), .A3(new_n743), .A4(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(G122), .Z(G24));
  NAND4_X1  g587(.A1(new_n647), .A2(KEYINPUT104), .A3(new_n566), .A4(new_n683), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT104), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n729), .A2(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n768), .B1(G472), .B2(new_n621), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n777), .A2(new_n669), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n756), .B1(new_n755), .B2(new_n677), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n740), .A2(KEYINPUT102), .A3(new_n636), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G125), .ZN(G27));
  NOR2_X1   g597(.A1(new_n502), .A2(new_n511), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n720), .A2(new_n784), .A3(new_n721), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT42), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n777), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n364), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n259), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n681), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n777), .A2(new_n445), .A3(new_n784), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT42), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G131), .ZN(G33));
  NAND3_X1  g608(.A1(new_n364), .A2(new_n687), .A3(new_n785), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G134), .ZN(G36));
  INV_X1    g610(.A(new_n385), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT75), .B1(new_n389), .B2(new_n391), .ZN(new_n798));
  AND4_X1   g612(.A1(KEYINPUT75), .A2(new_n391), .A3(new_n273), .A4(new_n388), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n372), .B1(new_n426), .B2(new_n427), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT78), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n413), .A2(new_n397), .A3(new_n372), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n804), .A2(new_n370), .B1(new_n425), .B2(new_n430), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n803), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n370), .B1(new_n806), .B2(new_n396), .ZN(new_n807));
  OAI22_X1  g621(.A1(new_n805), .A2(new_n420), .B1(new_n734), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT45), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n369), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT45), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT105), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT105), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n441), .A2(new_n442), .A3(new_n813), .A4(KEYINPUT45), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n810), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT106), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT106), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n810), .A2(new_n812), .A3(new_n817), .A4(new_n814), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n439), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT46), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n738), .A2(G469), .A3(G902), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n439), .A2(new_n822), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n824), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n368), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n566), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT107), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n647), .B(new_n828), .C1(new_n829), .C2(KEYINPUT43), .ZN(new_n830));
  XNOR2_X1  g644(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n728), .A2(new_n638), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n833), .B2(new_n566), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n690), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n627), .A3(new_n629), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT44), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n784), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n837), .B2(new_n838), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n827), .A2(new_n839), .A3(new_n718), .A4(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G137), .ZN(G39));
  NAND2_X1  g657(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n819), .A2(new_n825), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n438), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT46), .B1(new_n819), .B2(new_n820), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n721), .B(new_n844), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n363), .A2(new_n263), .A3(new_n730), .A4(new_n784), .ZN(new_n849));
  INV_X1    g663(.A(new_n844), .ZN(new_n850));
  NOR2_X1   g664(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n848), .B(new_n849), .C1(new_n827), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(G140), .ZN(G42));
  INV_X1    g668(.A(G952), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n230), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n740), .A2(new_n840), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n504), .B1(new_n830), .B2(new_n834), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n681), .A3(new_n789), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT48), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n858), .A2(new_n789), .A3(new_n778), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n759), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n857), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n705), .A2(new_n261), .A3(new_n262), .A4(new_n505), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n864), .A2(new_n865), .A3(new_n648), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n866), .A2(new_n855), .A3(G953), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n861), .A2(new_n863), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n865), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n647), .A2(new_n566), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n857), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n871), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n864), .A2(new_n865), .A3(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n690), .A2(new_n764), .A3(new_n768), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n876), .A2(KEYINPUT116), .B1(new_n877), .B2(new_n859), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n740), .A2(new_n510), .A3(new_n694), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n862), .A2(new_n879), .A3(KEYINPUT50), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT50), .ZN(new_n881));
  INV_X1    g695(.A(new_n694), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n755), .A2(new_n511), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n858), .A2(new_n789), .A3(new_n778), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT115), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n886), .B1(new_n880), .B2(new_n885), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n874), .B(new_n878), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n848), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n823), .A2(new_n826), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n852), .B1(new_n891), .B2(new_n721), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n739), .A2(new_n438), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n890), .A2(new_n892), .B1(new_n721), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n862), .A2(new_n784), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT114), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n889), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n869), .B1(new_n897), .B2(KEYINPUT51), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n876), .A2(KEYINPUT116), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n859), .A2(new_n877), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n874), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT117), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT117), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n878), .A2(new_n903), .A3(new_n874), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n880), .A2(new_n885), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n902), .A2(KEYINPUT51), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n896), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n894), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n721), .B1(new_n846), .B2(new_n847), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n851), .B2(new_n850), .ZN(new_n911));
  INV_X1    g725(.A(new_n893), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n911), .A2(new_n848), .B1(new_n368), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT118), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n906), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT119), .B1(new_n898), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n889), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n913), .B2(new_n907), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT51), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n868), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n906), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n896), .B1(new_n913), .B2(KEYINPUT118), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n894), .A2(new_n908), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n920), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n916), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT110), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n445), .A2(new_n616), .A3(new_n671), .A4(new_n672), .ZN(new_n929));
  AOI22_X1  g743(.A1(new_n929), .A2(new_n630), .B1(new_n364), .B2(new_n617), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n612), .A2(new_n613), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n648), .B1(new_n566), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n933), .A2(new_n502), .A3(new_n512), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n620), .A2(new_n630), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n928), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n928), .A2(new_n935), .A3(new_n618), .A4(new_n674), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n772), .B1(new_n746), .B2(new_n659), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n939), .B(new_n762), .C1(new_n747), .C2(new_n749), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT111), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n778), .A2(new_n669), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n941), .B1(new_n791), .B2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n785), .A2(new_n877), .A3(KEYINPUT111), .A4(new_n777), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n761), .A2(new_n932), .A3(new_n685), .A4(new_n785), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n793), .A2(new_n795), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n938), .A2(new_n940), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n683), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n770), .A2(new_n669), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n445), .A3(new_n714), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n782), .A2(new_n688), .A3(new_n731), .A4(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT52), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT112), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n952), .A2(new_n955), .A3(new_n953), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n952), .B2(new_n953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT53), .B1(new_n948), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n618), .A2(new_n674), .ZN(new_n960));
  INV_X1    g774(.A(new_n935), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT110), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n930), .A2(new_n928), .A3(new_n935), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n945), .A2(new_n946), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n788), .A2(new_n795), .A3(new_n792), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n772), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n762), .A2(new_n753), .A3(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n964), .A2(new_n750), .A3(new_n967), .A4(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n952), .B(KEYINPUT52), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT53), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(KEYINPUT54), .B1(new_n959), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n948), .A2(KEYINPUT53), .A3(new_n958), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n972), .B1(new_n970), .B2(new_n971), .ZN(new_n976));
  XOR2_X1   g790(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n856), .B1(new_n927), .B2(new_n979), .ZN(new_n980));
  NOR4_X1   g794(.A1(new_n833), .A2(new_n566), .A3(new_n368), .A4(new_n511), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT49), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n789), .B(new_n981), .C1(new_n912), .C2(new_n982), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT109), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n912), .A2(new_n982), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n984), .A2(new_n705), .A3(new_n882), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n980), .A2(new_n986), .ZN(G75));
  XNOR2_X1  g801(.A(new_n495), .B(new_n453), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT55), .Z(new_n989));
  INV_X1    g803(.A(G210), .ZN(new_n990));
  AOI211_X1 g804(.A(new_n990), .B(new_n241), .C1(new_n975), .C2(new_n976), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n989), .B1(new_n991), .B2(KEYINPUT56), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n241), .B1(new_n975), .B2(new_n976), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(G210), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT56), .ZN(new_n995));
  INV_X1    g809(.A(new_n989), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n230), .A2(G952), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n992), .A2(new_n997), .A3(new_n999), .ZN(G51));
  XNOR2_X1  g814(.A(new_n439), .B(KEYINPUT120), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT57), .Z(new_n1002));
  AND3_X1   g816(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n977), .B1(new_n975), .B2(new_n976), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n738), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n993), .A2(new_n818), .A3(new_n816), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n998), .B1(new_n1007), .B2(new_n1008), .ZN(G54));
  AND2_X1   g823(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n993), .A2(new_n559), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n559), .B1(new_n993), .B2(new_n1010), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1011), .A2(new_n1012), .A3(new_n998), .ZN(G60));
  NOR2_X1   g827(.A1(new_n726), .A2(new_n727), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n637), .B(KEYINPUT59), .Z(new_n1015));
  OAI211_X1 g829(.A(new_n1014), .B(new_n1015), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n999), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1014), .B1(new_n979), .B2(new_n1015), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1017), .A2(new_n1018), .ZN(G63));
  INV_X1    g833(.A(KEYINPUT61), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G217), .A2(G902), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT60), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1022), .B1(new_n975), .B2(new_n976), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n665), .A2(new_n666), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n999), .B1(new_n1023), .B2(new_n256), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1020), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n975), .A2(new_n976), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n255), .B1(new_n1029), .B2(new_n1022), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1030), .A2(KEYINPUT61), .A3(new_n999), .A4(new_n1025), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1028), .A2(new_n1031), .ZN(G66));
  INV_X1    g846(.A(new_n508), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n230), .B1(new_n1033), .B2(G224), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n938), .A2(new_n940), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1034), .B1(new_n1036), .B2(new_n230), .ZN(new_n1037));
  OAI211_X1 g851(.A(new_n465), .B(new_n471), .C1(G898), .C2(new_n230), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(KEYINPUT121), .Z(new_n1039));
  XNOR2_X1  g853(.A(new_n1037), .B(new_n1039), .ZN(G69));
  NAND2_X1  g854(.A1(new_n297), .A2(new_n302), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT122), .Z(new_n1042));
  XNOR2_X1  g856(.A(new_n1042), .B(new_n548), .ZN(new_n1043));
  NAND2_X1  g857(.A1(G900), .A2(G953), .ZN(new_n1044));
  AND2_X1   g858(.A1(new_n853), .A2(new_n842), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n671), .A2(new_n677), .A3(new_n672), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n720), .A2(new_n721), .ZN(new_n1047));
  NOR3_X1   g861(.A1(new_n1046), .A2(new_n363), .A3(new_n1047), .ZN(new_n1048));
  AOI22_X1  g862(.A1(new_n759), .A2(new_n779), .B1(new_n1048), .B2(new_n687), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1049), .A2(new_n731), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n1050), .A2(new_n966), .ZN(new_n1051));
  NOR2_X1   g865(.A1(new_n790), .A2(new_n770), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n827), .A2(new_n718), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1045), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  OAI211_X1 g868(.A(new_n1043), .B(new_n1044), .C1(new_n1054), .C2(G953), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n724), .A2(new_n782), .A3(new_n688), .A4(new_n731), .ZN(new_n1056));
  INV_X1    g870(.A(KEYINPUT123), .ZN(new_n1057));
  AND3_X1   g871(.A1(new_n1056), .A2(new_n1057), .A3(KEYINPUT62), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n1057), .B1(new_n1056), .B2(KEYINPUT62), .ZN(new_n1059));
  NOR2_X1   g873(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g874(.A(KEYINPUT62), .ZN(new_n1061));
  NAND4_X1  g875(.A1(new_n1049), .A2(new_n1061), .A3(new_n724), .A4(new_n731), .ZN(new_n1062));
  INV_X1    g876(.A(new_n722), .ZN(new_n1063));
  NAND4_X1  g877(.A1(new_n364), .A2(new_n1063), .A3(new_n784), .A4(new_n933), .ZN(new_n1064));
  NAND4_X1  g878(.A1(new_n853), .A2(new_n1062), .A3(new_n842), .A4(new_n1064), .ZN(new_n1065));
  OAI21_X1  g879(.A(KEYINPUT124), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n1056), .A2(KEYINPUT62), .ZN(new_n1067));
  NAND2_X1  g881(.A1(new_n1067), .A2(KEYINPUT123), .ZN(new_n1068));
  NAND3_X1  g882(.A1(new_n1056), .A2(new_n1057), .A3(KEYINPUT62), .ZN(new_n1069));
  NAND2_X1  g883(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g884(.A(KEYINPUT124), .ZN(new_n1071));
  AND2_X1   g885(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1072));
  NAND4_X1  g886(.A1(new_n1070), .A2(new_n1045), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g887(.A(G953), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g888(.A(new_n1055), .B1(new_n1074), .B2(new_n1043), .ZN(new_n1075));
  AOI21_X1  g889(.A(new_n230), .B1(G227), .B2(G900), .ZN(new_n1076));
  INV_X1    g890(.A(KEYINPUT125), .ZN(new_n1077));
  AOI21_X1  g891(.A(new_n1076), .B1(new_n1055), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g892(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g893(.A(new_n1055), .B1(new_n1077), .B2(new_n1076), .C1(new_n1074), .C2(new_n1043), .ZN(new_n1080));
  AND2_X1   g894(.A1(new_n1079), .A2(new_n1080), .ZN(G72));
  NAND2_X1  g895(.A1(G472), .A2(G902), .ZN(new_n1082));
  XOR2_X1   g896(.A(new_n1082), .B(KEYINPUT63), .Z(new_n1083));
  OAI21_X1  g897(.A(new_n1083), .B1(new_n1054), .B2(new_n1036), .ZN(new_n1084));
  XNOR2_X1  g898(.A(new_n360), .B(KEYINPUT127), .ZN(new_n1085));
  AOI21_X1  g899(.A(new_n998), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g900(.A1(new_n959), .A2(new_n973), .ZN(new_n1087));
  NAND3_X1  g901(.A1(new_n700), .A2(new_n360), .A3(new_n1083), .ZN(new_n1088));
  OAI21_X1  g902(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g903(.A1(new_n1066), .A2(new_n1073), .A3(new_n1035), .ZN(new_n1090));
  NAND2_X1  g904(.A1(new_n1090), .A2(new_n1083), .ZN(new_n1091));
  INV_X1    g905(.A(new_n700), .ZN(new_n1092));
  NAND2_X1  g906(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g907(.A(KEYINPUT126), .ZN(new_n1094));
  NAND2_X1  g908(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g909(.A1(new_n1091), .A2(KEYINPUT126), .A3(new_n1092), .ZN(new_n1096));
  AOI21_X1  g910(.A(new_n1089), .B1(new_n1095), .B2(new_n1096), .ZN(G57));
endmodule


