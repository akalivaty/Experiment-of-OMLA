//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  XOR2_X1   g000(.A(G78gat), .B(G106gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT31), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G141gat), .B(G148gat), .Z(new_n207));
  AOI21_X1  g006(.A(KEYINPUT75), .B1(KEYINPUT76), .B2(KEYINPUT2), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(KEYINPUT76), .B2(KEYINPUT2), .ZN(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n207), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  XOR2_X1   g012(.A(new_n213), .B(KEYINPUT75), .Z(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n211), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n215), .B2(KEYINPUT2), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n212), .A2(new_n214), .B1(new_n216), .B2(new_n207), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT29), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G197gat), .B(G204gat), .ZN(new_n220));
  INV_X1    g019(.A(G211gat), .ZN(new_n221));
  INV_X1    g020(.A(G218gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(KEYINPUT22), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G211gat), .B(G218gat), .Z(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT80), .B1(new_n219), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(G228gat), .A3(G233gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT29), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT3), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  OAI22_X1  g029(.A1(new_n230), .A2(new_n217), .B1(new_n219), .B2(new_n226), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n231), .A2(G228gat), .A3(G233gat), .A4(new_n227), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n233), .A2(G22gat), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(G22gat), .B1(new_n233), .B2(new_n234), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n206), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT81), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI211_X1 g038(.A(KEYINPUT81), .B(new_n206), .C1(new_n235), .C2(new_n236), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n205), .B1(new_n236), .B2(KEYINPUT82), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n235), .B1(KEYINPUT82), .B2(new_n236), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT83), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n236), .A2(KEYINPUT82), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n233), .A2(G22gat), .A3(new_n234), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT83), .B1(new_n249), .B2(new_n242), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n241), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n252));
  XNOR2_X1  g051(.A(G1gat), .B(G29gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G57gat), .B(G85gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  XOR2_X1   g055(.A(G113gat), .B(G120gat), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT70), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259));
  XNOR2_X1  g058(.A(G113gat), .B(G120gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT68), .B(G127gat), .ZN(new_n264));
  INV_X1    g063(.A(G134gat), .ZN(new_n265));
  OR3_X1    g064(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(G127gat), .ZN(new_n267));
  OAI211_X1 g066(.A(KEYINPUT69), .B(new_n267), .C1(new_n264), .C2(new_n265), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G127gat), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT1), .B1(new_n270), .B2(G134gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n257), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n217), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT4), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n269), .A2(new_n217), .A3(new_n275), .A4(new_n272), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n212), .A2(new_n214), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n216), .A2(new_n207), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI22_X1  g078(.A1(KEYINPUT3), .A2(new_n279), .B1(new_n269), .B2(new_n272), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n217), .A2(new_n218), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n274), .A2(new_n276), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G225gat), .A2(G233gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n273), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n217), .B1(new_n269), .B2(new_n272), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n282), .A2(new_n283), .B1(new_n287), .B2(KEYINPUT77), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT77), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n292), .B(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n282), .A2(new_n283), .B1(new_n293), .B2(new_n289), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n256), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n294), .ZN(new_n296));
  INV_X1    g095(.A(new_n256), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n296), .B(new_n297), .C1(new_n290), .C2(new_n288), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n295), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n291), .A2(new_n294), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(KEYINPUT6), .A3(new_n297), .ZN(new_n302));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(new_n304), .B2(KEYINPUT23), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT64), .B(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(G169gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(KEYINPUT23), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n305), .B1(new_n308), .B2(KEYINPUT65), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT65), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n306), .A2(new_n311), .A3(KEYINPUT23), .A4(new_n307), .ZN(new_n312));
  NAND2_X1  g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(KEYINPUT24), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n313), .A2(KEYINPUT24), .ZN(new_n315));
  INV_X1    g114(.A(G183gat), .ZN(new_n316));
  INV_X1    g115(.A(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n309), .A2(new_n310), .A3(new_n312), .A4(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT26), .ZN(new_n321));
  OR3_X1    g120(.A1(new_n304), .A2(KEYINPUT67), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT67), .B1(new_n304), .B2(new_n321), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n321), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .A4(new_n303), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT27), .B(G183gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT28), .B1(new_n327), .B2(G190gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n316), .A2(KEYINPUT27), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT28), .B1(new_n329), .B2(KEYINPUT66), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n330), .B(new_n317), .C1(KEYINPUT66), .C2(new_n326), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n325), .A2(new_n328), .A3(new_n331), .A4(new_n313), .ZN(new_n332));
  INV_X1    g131(.A(new_n319), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n304), .A2(KEYINPUT23), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n334), .A2(new_n305), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT25), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(G226gat), .A2(G233gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n337), .B2(new_n229), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n226), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n337), .A2(KEYINPUT73), .A3(new_n338), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n341), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n344), .B1(new_n348), .B2(new_n343), .ZN(new_n349));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT74), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(G64gat), .ZN(new_n352));
  INV_X1    g151(.A(G92gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n344), .B(new_n354), .C1(new_n348), .C2(new_n343), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(KEYINPUT30), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n349), .A2(new_n359), .A3(new_n355), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n300), .A2(new_n302), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n337), .A2(new_n269), .A3(new_n272), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n269), .A2(new_n272), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n363), .A2(new_n332), .A3(new_n320), .A4(new_n336), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n362), .A2(new_n364), .A3(G227gat), .A4(G233gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT32), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT33), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G15gat), .B(G43gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(G71gat), .ZN(new_n370));
  INV_X1    g169(.A(G99gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n366), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(KEYINPUT33), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n365), .A2(KEYINPUT32), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(KEYINPUT71), .A3(new_n375), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n362), .A2(new_n364), .B1(G227gat), .B2(G233gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n377), .B(KEYINPUT34), .Z(new_n378));
  INV_X1    g177(.A(KEYINPUT71), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n366), .A2(new_n368), .A3(new_n379), .A4(new_n372), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n376), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n378), .B1(new_n376), .B2(new_n380), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n251), .A2(new_n361), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT35), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n251), .A2(new_n361), .A3(KEYINPUT35), .A4(new_n383), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT86), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n358), .A2(new_n360), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n282), .B2(new_n283), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n274), .A2(new_n276), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n280), .A2(new_n281), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(KEYINPUT84), .A3(new_n284), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT39), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n285), .A2(new_n286), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n397), .B1(new_n398), .B2(new_n283), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n392), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n282), .A2(new_n391), .A3(new_n283), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT84), .B1(new_n395), .B2(new_n284), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n397), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT85), .B1(new_n403), .B2(new_n256), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT39), .B1(new_n392), .B2(new_n396), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n405), .A2(new_n406), .A3(new_n297), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n400), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT40), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n390), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n400), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n403), .A2(KEYINPUT85), .A3(new_n256), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n406), .B1(new_n405), .B2(new_n297), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n298), .B1(new_n414), .B2(KEYINPUT40), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n389), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n358), .A2(new_n360), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n414), .B2(KEYINPUT40), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n408), .A2(new_n409), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT86), .A4(new_n298), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT37), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n348), .B2(new_n343), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(new_n343), .B2(new_n342), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT87), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT88), .B(KEYINPUT37), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n349), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n355), .A2(KEYINPUT38), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n300), .A2(new_n302), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n426), .B1(new_n421), .B2(new_n349), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT38), .B1(new_n430), .B2(new_n355), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n428), .A2(new_n429), .A3(new_n356), .A4(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n416), .A2(new_n420), .A3(new_n251), .A4(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT72), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT36), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n383), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n438), .B(new_n439), .C1(new_n381), .C2(new_n382), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n436), .B(new_n440), .C1(new_n361), .C2(new_n251), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n388), .B1(new_n433), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G229gat), .A2(G233gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(KEYINPUT13), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT95), .ZN(new_n447));
  XNOR2_X1  g246(.A(G15gat), .B(G22gat), .ZN(new_n448));
  INV_X1    g247(.A(G1gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT16), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n448), .A2(G1gat), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n451), .A2(new_n452), .A3(G8gat), .ZN(new_n453));
  INV_X1    g252(.A(G8gat), .ZN(new_n454));
  XOR2_X1   g253(.A(G15gat), .B(G22gat), .Z(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n449), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(new_n450), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n447), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(G8gat), .B1(new_n451), .B2(new_n452), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n456), .A2(new_n454), .A3(new_n457), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT95), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G29gat), .ZN(new_n464));
  INV_X1    g263(.A(G36gat), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT14), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT14), .ZN(new_n468));
  XOR2_X1   g267(.A(KEYINPUT91), .B(G36gat), .Z(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT90), .B(G29gat), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n467), .B(new_n468), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n204), .A2(KEYINPUT92), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT92), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(G50gat), .ZN(new_n474));
  INV_X1    g273(.A(G43gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT93), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n475), .B2(G50gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT15), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n472), .A2(new_n474), .A3(KEYINPUT93), .A4(new_n475), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n475), .A2(G50gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n204), .A2(G43gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT15), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n471), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n471), .A2(new_n486), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT94), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT94), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n486), .ZN(new_n491));
  INV_X1    g290(.A(new_n486), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n482), .A2(new_n481), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(new_n480), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n490), .B(new_n491), .C1(new_n494), .C2(new_n471), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n463), .A2(new_n489), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n463), .B1(new_n489), .B2(new_n495), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n446), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT97), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(KEYINPUT97), .B(new_n446), .C1(new_n496), .C2(new_n497), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n496), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT96), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT18), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n504), .A2(new_n505), .B1(G229gat), .B2(G233gat), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT17), .B1(new_n489), .B2(new_n495), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n487), .A2(new_n488), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n453), .A2(new_n458), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n503), .B(new_n506), .C1(new_n510), .C2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n504), .A2(new_n505), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT94), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n482), .A2(new_n481), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT92), .B(G50gat), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n478), .B1(new_n519), .B2(new_n475), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n486), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n471), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n490), .B1(new_n523), .B2(new_n491), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n508), .B1(new_n517), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n509), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n511), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n528), .A2(new_n514), .A3(new_n503), .A4(new_n506), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n502), .A2(new_n516), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT89), .B(G197gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT11), .B(G169gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT12), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n502), .A2(new_n516), .A3(new_n529), .A4(new_n536), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G230gat), .ZN(new_n542));
  INV_X1    g341(.A(G233gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT7), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(G85gat), .A3(G92gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  INV_X1    g350(.A(G85gat), .ZN(new_n552));
  AOI22_X1  g351(.A1(KEYINPUT8), .A2(new_n551), .B1(new_n552), .B2(new_n353), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G99gat), .B(G106gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n550), .A2(new_n553), .A3(new_n555), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(KEYINPUT99), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n555), .B1(new_n550), .B2(new_n553), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT99), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n559), .A2(KEYINPUT100), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT100), .B1(new_n559), .B2(new_n562), .ZN(new_n564));
  NAND2_X1  g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  OR2_X1    g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G64gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(G57gat), .ZN(new_n570));
  INV_X1    g369(.A(G57gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(G64gat), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n570), .A2(new_n572), .A3(KEYINPUT98), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT98), .B1(new_n570), .B2(new_n572), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n568), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n570), .A2(new_n572), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n565), .B(new_n566), .C1(new_n576), .C2(new_n567), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n577), .A3(KEYINPUT10), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n563), .A2(new_n564), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(new_n577), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n550), .A2(new_n555), .A3(new_n553), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n581), .A2(new_n560), .A3(new_n561), .ZN(new_n582));
  INV_X1    g381(.A(new_n562), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n575), .B(new_n577), .C1(new_n581), .C2(new_n560), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT10), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n545), .B1(new_n579), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(new_n544), .A3(new_n585), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G120gat), .B(G148gat), .ZN(new_n590));
  INV_X1    g389(.A(G176gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(G204gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n587), .A2(new_n588), .A3(new_n593), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n541), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n443), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G190gat), .B(G218gat), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n563), .A2(new_n564), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(new_n525), .B2(new_n526), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n489), .A2(new_n495), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(new_n582), .B2(new_n583), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n559), .A2(KEYINPUT100), .A3(new_n562), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT41), .ZN(new_n610));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611));
  OAI22_X1  g410(.A1(new_n605), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n602), .B1(new_n604), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n611), .A2(new_n610), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n517), .A2(new_n524), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n614), .B1(new_n615), .B2(new_n603), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n609), .B1(new_n507), .B2(new_n509), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n617), .A3(new_n601), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n611), .A2(new_n610), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  NAND4_X1  g420(.A1(new_n613), .A2(KEYINPUT101), .A3(new_n618), .A4(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n625), .A2(new_n621), .B1(new_n613), .B2(new_n618), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT21), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n580), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G127gat), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n459), .B(new_n462), .C1(new_n629), .C2(new_n580), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g433(.A(G155gat), .B(G183gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n633), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(new_n221), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n638), .A2(new_n642), .A3(new_n639), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n628), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n600), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n429), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(new_n449), .ZN(G1324gat));
  INV_X1    g450(.A(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n390), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(G8gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT102), .B(G8gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  MUX2_X1   g457(.A(new_n655), .B(KEYINPUT42), .S(new_n658), .Z(G1325gat));
  NAND2_X1  g458(.A1(new_n436), .A2(new_n440), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n652), .A2(G15gat), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n600), .A2(new_n647), .A3(new_n383), .ZN(new_n668));
  INV_X1    g467(.A(G15gat), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n668), .A2(KEYINPUT103), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT103), .B1(new_n668), .B2(new_n669), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n667), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1326gat));
  INV_X1    g473(.A(G22gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n251), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n600), .A2(new_n647), .A3(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(KEYINPUT106), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(KEYINPUT106), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n679), .B1(new_n678), .B2(new_n680), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n675), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n678), .A2(new_n680), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT43), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(G22gat), .A3(new_n681), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(G1327gat));
  NAND3_X1  g487(.A1(new_n600), .A2(new_n628), .A3(new_n646), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n429), .A3(new_n470), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT44), .B1(new_n443), .B2(new_n627), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n433), .A2(new_n442), .ZN(new_n696));
  INV_X1    g495(.A(new_n388), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT109), .B1(new_n623), .B2(new_n626), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n613), .A2(new_n618), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n612), .B1(new_n527), .B2(new_n609), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT101), .B1(new_n701), .B2(new_n601), .ZN(new_n702));
  INV_X1    g501(.A(new_n621), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n705), .A3(new_n622), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT44), .B1(new_n699), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n698), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n695), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n646), .B(KEYINPUT108), .Z(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n598), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n694), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  AOI211_X1 g512(.A(KEYINPUT110), .B(new_n711), .C1(new_n695), .C2(new_n708), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n649), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n693), .B1(new_n716), .B2(new_n470), .ZN(G1328gat));
  NAND3_X1  g516(.A1(new_n690), .A2(new_n469), .A3(new_n390), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT46), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n718), .A2(KEYINPUT46), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n715), .A2(new_n417), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n719), .B(new_n720), .C1(new_n721), .C2(new_n469), .ZN(G1329gat));
  INV_X1    g521(.A(new_n383), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n689), .A2(G43gat), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n709), .A2(new_n660), .A3(new_n712), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n725), .B(KEYINPUT47), .C1(new_n475), .C2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n666), .B1(new_n713), .B2(new_n714), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n724), .B1(new_n728), .B2(G43gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n729), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g529(.A1(new_n709), .A2(new_n676), .A3(new_n712), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n709), .A2(KEYINPUT111), .A3(new_n676), .A4(new_n712), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n519), .A3(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n689), .A2(new_n519), .A3(new_n251), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n735), .A2(KEYINPUT48), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n676), .B1(new_n713), .B2(new_n714), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n736), .B1(new_n739), .B2(new_n519), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n740), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g540(.A1(new_n443), .A2(new_n628), .A3(new_n646), .A4(new_n540), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n597), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n649), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(new_n571), .ZN(G1332gat));
  INV_X1    g544(.A(KEYINPUT49), .ZN(new_n746));
  NAND2_X1  g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n417), .B(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n742), .A2(new_n597), .A3(new_n747), .A4(new_n749), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n750), .A2(KEYINPUT113), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(KEYINPUT113), .ZN(new_n752));
  AND4_X1   g551(.A1(new_n746), .A2(new_n751), .A3(new_n569), .A4(new_n752), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n751), .A2(new_n752), .B1(new_n746), .B2(new_n569), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(G1333gat));
  OR3_X1    g554(.A1(new_n743), .A2(G71gat), .A3(new_n723), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n757));
  OAI21_X1  g556(.A(G71gat), .B1(new_n743), .B2(new_n665), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(G1334gat));
  NOR2_X1   g560(.A1(new_n743), .A2(new_n251), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT114), .B(G78gat), .Z(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1335gat));
  INV_X1    g563(.A(new_n646), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n765), .A2(new_n540), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n698), .A2(new_n628), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n767), .B2(new_n768), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n774), .A2(new_n552), .A3(new_n429), .A4(new_n597), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n709), .A2(new_n597), .A3(new_n766), .ZN(new_n776));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n649), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1336gat));
  NOR2_X1   g577(.A1(new_n776), .A2(new_n417), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n353), .ZN(new_n780));
  INV_X1    g579(.A(new_n749), .ZN(new_n781));
  INV_X1    g580(.A(new_n597), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n781), .A2(G92gat), .A3(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n769), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT52), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  OAI21_X1  g585(.A(G92gat), .B1(new_n776), .B2(new_n781), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(new_n788));
  INV_X1    g587(.A(new_n783), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n786), .B(new_n787), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n785), .A2(new_n790), .ZN(G1337gat));
  NAND4_X1  g590(.A1(new_n774), .A2(new_n371), .A3(new_n597), .A4(new_n383), .ZN(new_n792));
  OAI21_X1  g591(.A(G99gat), .B1(new_n776), .B2(new_n665), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(G1338gat));
  NAND2_X1  g593(.A1(KEYINPUT116), .A2(G106gat), .ZN(new_n795));
  OR2_X1    g594(.A1(KEYINPUT116), .A2(G106gat), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n795), .B(new_n796), .C1(new_n776), .C2(new_n251), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n251), .A2(G106gat), .A3(new_n782), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n769), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT53), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  INV_X1    g601(.A(new_n798), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n802), .B(new_n797), .C1(new_n788), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(G1339gat));
  NAND3_X1  g604(.A1(new_n647), .A2(new_n782), .A3(new_n541), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n699), .A2(new_n706), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT10), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n559), .A2(new_n562), .B1(new_n575), .B2(new_n577), .ZN(new_n810));
  INV_X1    g609(.A(new_n585), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n578), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n607), .A2(new_n608), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n814), .A3(new_n544), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n587), .A2(KEYINPUT54), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n544), .B1(new_n812), .B2(new_n814), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n593), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n816), .A2(new_n819), .A3(KEYINPUT55), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n596), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n822), .A2(new_n596), .A3(KEYINPUT117), .A4(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n444), .B1(new_n528), .B2(new_n503), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n496), .A2(new_n497), .A3(new_n446), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n535), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n539), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n808), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n828), .A2(new_n540), .B1(new_n597), .B2(new_n832), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n808), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n807), .B1(new_n835), .B2(new_n710), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n781), .A2(new_n429), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n676), .A2(new_n723), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n540), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n597), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(G120gat), .ZN(G1341gat));
  INV_X1    g644(.A(new_n264), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n840), .A2(new_n846), .A3(new_n710), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n841), .A2(new_n765), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n846), .B2(new_n848), .ZN(G1342gat));
  NOR2_X1   g648(.A1(new_n390), .A2(new_n627), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n429), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI211_X1 g651(.A(new_n852), .B(new_n836), .C1(new_n851), .C2(new_n850), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n265), .A3(new_n839), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n840), .B2(new_n627), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  NAND2_X1  g657(.A1(new_n665), .A2(new_n676), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n838), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(G141gat), .A3(new_n541), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT58), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n816), .A2(new_n819), .A3(KEYINPUT55), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT55), .B1(new_n816), .B2(new_n819), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT117), .B1(new_n867), .B2(new_n596), .ZN(new_n868));
  INV_X1    g667(.A(new_n827), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n540), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n832), .A2(new_n597), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n808), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n808), .A2(new_n828), .A3(new_n832), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n710), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n251), .B1(new_n874), .B2(new_n806), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT119), .B1(new_n875), .B2(KEYINPUT57), .ZN(new_n876));
  INV_X1    g675(.A(new_n824), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n540), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n628), .B1(new_n878), .B2(new_n871), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n806), .B1(new_n880), .B2(new_n765), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(KEYINPUT57), .A3(new_n676), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n883), .B(new_n884), .C1(new_n836), .C2(new_n251), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n876), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n837), .A2(new_n660), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n540), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G141gat), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n864), .B(new_n889), .C1(new_n863), .C2(new_n862), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n888), .A2(new_n891), .A3(G141gat), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n888), .B2(G141gat), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(new_n862), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n890), .B1(new_n894), .B2(new_n895), .ZN(G1344gat));
  OR3_X1    g695(.A1(new_n861), .A2(G148gat), .A3(new_n782), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n628), .A2(new_n877), .A3(new_n832), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n879), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n807), .B1(new_n900), .B2(new_n646), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n884), .B1(new_n901), .B2(new_n251), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n875), .A2(KEYINPUT57), .ZN(new_n905));
  OAI211_X1 g704(.A(KEYINPUT122), .B(new_n884), .C1(new_n901), .C2(new_n251), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n597), .A3(new_n887), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n898), .B1(new_n908), .B2(G148gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n886), .A2(new_n597), .A3(new_n887), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n910), .A2(new_n898), .A3(G148gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n897), .B1(new_n909), .B2(new_n911), .ZN(G1345gat));
  OAI21_X1  g711(.A(new_n210), .B1(new_n861), .B2(new_n646), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n710), .A2(new_n210), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n886), .A2(new_n887), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT123), .ZN(G1346gat));
  NAND3_X1  g716(.A1(new_n853), .A2(new_n211), .A3(new_n860), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n886), .A2(new_n808), .A3(new_n887), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n211), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n836), .A2(new_n429), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n839), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n749), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n540), .A2(new_n307), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n922), .A2(new_n541), .A3(new_n417), .ZN(new_n926));
  OAI22_X1  g725(.A1(new_n924), .A2(new_n925), .B1(new_n926), .B2(new_n307), .ZN(G1348gat));
  NAND3_X1  g726(.A1(new_n923), .A2(new_n597), .A3(new_n749), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n922), .A2(new_n417), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n782), .A2(new_n306), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n928), .A2(new_n591), .B1(new_n929), .B2(new_n930), .ZN(G1349gat));
  NAND2_X1  g730(.A1(new_n765), .A2(new_n326), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n922), .A2(new_n417), .A3(new_n710), .ZN(new_n933));
  OAI22_X1  g732(.A1(new_n924), .A2(new_n932), .B1(new_n933), .B2(new_n316), .ZN(new_n934));
  NAND2_X1  g733(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n934), .B(new_n935), .Z(G1350gat));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n929), .A2(new_n628), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(G190gat), .ZN(new_n939));
  AOI211_X1 g738(.A(KEYINPUT61), .B(new_n317), .C1(new_n929), .C2(new_n628), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n808), .A2(new_n317), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n939), .A2(new_n940), .B1(new_n924), .B2(new_n941), .ZN(G1351gat));
  NAND2_X1  g741(.A1(new_n907), .A2(KEYINPUT125), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n666), .A2(new_n429), .A3(new_n417), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n904), .A2(new_n945), .A3(new_n905), .A4(new_n906), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n541), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n921), .A2(new_n749), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(new_n859), .ZN(new_n950));
  INV_X1    g749(.A(G197gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(new_n951), .A3(new_n540), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n948), .A2(new_n952), .ZN(G1352gat));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n950), .A2(new_n597), .ZN(new_n956));
  XNOR2_X1  g755(.A(KEYINPUT126), .B(G204gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n958), .B(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n947), .B2(new_n782), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1353gat));
  NAND3_X1  g761(.A1(new_n950), .A2(new_n221), .A3(new_n765), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n907), .A2(new_n765), .A3(new_n944), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  NOR3_X1   g766(.A1(new_n947), .A2(new_n222), .A3(new_n627), .ZN(new_n968));
  AOI21_X1  g767(.A(G218gat), .B1(new_n950), .B2(new_n808), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(new_n969), .ZN(G1355gat));
endmodule


