

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592;

  NOR2_X1 U325 ( .A1(n388), .A2(n582), .ZN(n389) );
  XNOR2_X1 U326 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U327 ( .A(n309), .B(n308), .ZN(n310) );
  INV_X1 U328 ( .A(KEYINPUT26), .ZN(n465) );
  NOR2_X1 U329 ( .A1(n468), .A2(n528), .ZN(n466) );
  XNOR2_X1 U330 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U331 ( .A(n376), .B(n295), .ZN(n377) );
  XNOR2_X1 U332 ( .A(KEYINPUT119), .B(n448), .ZN(n550) );
  AND2_X1 U333 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  AND2_X1 U334 ( .A1(G228GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U335 ( .A(n375), .B(n374), .Z(n295) );
  XNOR2_X1 U336 ( .A(n387), .B(KEYINPUT45), .ZN(n388) );
  XOR2_X1 U337 ( .A(G162GAT), .B(G50GAT), .Z(n330) );
  XNOR2_X1 U338 ( .A(n330), .B(n294), .ZN(n302) );
  XNOR2_X1 U339 ( .A(n370), .B(n302), .ZN(n303) );
  XNOR2_X1 U340 ( .A(n335), .B(n293), .ZN(n336) );
  XNOR2_X1 U341 ( .A(n435), .B(G176GAT), .ZN(n436) );
  INV_X1 U342 ( .A(KEYINPUT22), .ZN(n308) );
  XNOR2_X1 U343 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U344 ( .A(n437), .B(n436), .ZN(n440) );
  INV_X1 U345 ( .A(KEYINPUT99), .ZN(n480) );
  NOR2_X1 U346 ( .A1(n522), .A2(n459), .ZN(n576) );
  XNOR2_X1 U347 ( .A(n378), .B(n377), .ZN(n380) );
  XNOR2_X1 U348 ( .A(n481), .B(n480), .ZN(n498) );
  XNOR2_X1 U349 ( .A(n444), .B(n443), .ZN(n445) );
  INV_X1 U350 ( .A(KEYINPUT58), .ZN(n462) );
  XOR2_X1 U351 ( .A(n346), .B(n379), .Z(n495) );
  XOR2_X1 U352 ( .A(n582), .B(KEYINPUT41), .Z(n557) );
  INV_X1 U353 ( .A(G43GAT), .ZN(n491) );
  XNOR2_X1 U354 ( .A(n462), .B(G190GAT), .ZN(n463) );
  XNOR2_X1 U355 ( .A(n453), .B(G134GAT), .ZN(n454) );
  XNOR2_X1 U356 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U357 ( .A(n464), .B(n463), .ZN(G1351GAT) );
  XNOR2_X1 U358 ( .A(n494), .B(n493), .ZN(G1330GAT) );
  XOR2_X1 U359 ( .A(G197GAT), .B(KEYINPUT21), .Z(n297) );
  XNOR2_X1 U360 ( .A(G211GAT), .B(KEYINPUT85), .ZN(n296) );
  XNOR2_X1 U361 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U362 ( .A(n298), .B(KEYINPUT86), .Z(n300) );
  XNOR2_X1 U363 ( .A(G218GAT), .B(G204GAT), .ZN(n299) );
  XNOR2_X1 U364 ( .A(n300), .B(n299), .ZN(n398) );
  XNOR2_X1 U365 ( .A(G148GAT), .B(G106GAT), .ZN(n301) );
  XNOR2_X1 U366 ( .A(n301), .B(G78GAT), .ZN(n370) );
  XOR2_X1 U367 ( .A(n303), .B(KEYINPUT88), .Z(n307) );
  XOR2_X1 U368 ( .A(G141GAT), .B(KEYINPUT87), .Z(n305) );
  XNOR2_X1 U369 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n304) );
  XNOR2_X1 U370 ( .A(n305), .B(n304), .ZN(n424) );
  XNOR2_X1 U371 ( .A(n424), .B(KEYINPUT23), .ZN(n306) );
  XNOR2_X1 U372 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U373 ( .A(G155GAT), .B(G22GAT), .Z(n321) );
  XNOR2_X1 U374 ( .A(n321), .B(KEYINPUT24), .ZN(n309) );
  XOR2_X1 U375 ( .A(n398), .B(n312), .Z(n468) );
  XOR2_X1 U376 ( .A(KEYINPUT28), .B(n468), .Z(n530) );
  XOR2_X1 U377 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n314) );
  XNOR2_X1 U378 ( .A(G71GAT), .B(G64GAT), .ZN(n313) );
  XNOR2_X1 U379 ( .A(n314), .B(n313), .ZN(n329) );
  XOR2_X1 U380 ( .A(G211GAT), .B(G78GAT), .Z(n316) );
  XOR2_X1 U381 ( .A(G183GAT), .B(G8GAT), .Z(n400) );
  XOR2_X1 U382 ( .A(G1GAT), .B(KEYINPUT68), .Z(n358) );
  XNOR2_X1 U383 ( .A(n400), .B(n358), .ZN(n315) );
  XNOR2_X1 U384 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U385 ( .A(G127GAT), .B(G15GAT), .Z(n442) );
  XOR2_X1 U386 ( .A(n317), .B(n442), .Z(n327) );
  XOR2_X1 U387 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n319) );
  XNOR2_X1 U388 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n318) );
  XNOR2_X1 U389 ( .A(n319), .B(n318), .ZN(n325) );
  XNOR2_X1 U390 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n320) );
  XNOR2_X1 U391 ( .A(n320), .B(KEYINPUT71), .ZN(n371) );
  XOR2_X1 U392 ( .A(n371), .B(n321), .Z(n323) );
  NAND2_X1 U393 ( .A1(G231GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U394 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U395 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U396 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U397 ( .A(n329), .B(n328), .ZN(n586) );
  INV_X1 U398 ( .A(n586), .ZN(n573) );
  XOR2_X1 U399 ( .A(KEYINPUT10), .B(G218GAT), .Z(n332) );
  XOR2_X1 U400 ( .A(G190GAT), .B(G36GAT), .Z(n401) );
  XNOR2_X1 U401 ( .A(n330), .B(n401), .ZN(n331) );
  XNOR2_X1 U402 ( .A(n332), .B(n331), .ZN(n337) );
  XOR2_X1 U403 ( .A(KEYINPUT77), .B(KEYINPUT64), .Z(n334) );
  XNOR2_X1 U404 ( .A(G134GAT), .B(G106GAT), .ZN(n333) );
  XNOR2_X1 U405 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U406 ( .A(n338), .B(KEYINPUT9), .Z(n342) );
  XOR2_X1 U407 ( .A(G43GAT), .B(KEYINPUT7), .Z(n340) );
  XNOR2_X1 U408 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n339) );
  XNOR2_X1 U409 ( .A(n340), .B(n339), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n357), .B(KEYINPUT11), .ZN(n341) );
  XNOR2_X1 U411 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U412 ( .A(KEYINPUT73), .B(G99GAT), .Z(n344) );
  XNOR2_X1 U413 ( .A(KEYINPUT74), .B(G92GAT), .ZN(n343) );
  XNOR2_X1 U414 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U415 ( .A(G85GAT), .B(n345), .ZN(n379) );
  INV_X1 U416 ( .A(n495), .ZN(n562) );
  XOR2_X1 U417 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n348) );
  XNOR2_X1 U418 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n347) );
  XNOR2_X1 U419 ( .A(n348), .B(n347), .ZN(n366) );
  XOR2_X1 U420 ( .A(G22GAT), .B(G36GAT), .Z(n350) );
  XNOR2_X1 U421 ( .A(G141GAT), .B(G50GAT), .ZN(n349) );
  XNOR2_X1 U422 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U423 ( .A(G197GAT), .B(G169GAT), .Z(n352) );
  XNOR2_X1 U424 ( .A(G113GAT), .B(G15GAT), .ZN(n351) );
  XNOR2_X1 U425 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U426 ( .A(n354), .B(n353), .Z(n364) );
  XOR2_X1 U427 ( .A(KEYINPUT65), .B(KEYINPUT69), .Z(n356) );
  XNOR2_X1 U428 ( .A(KEYINPUT67), .B(KEYINPUT70), .ZN(n355) );
  XNOR2_X1 U429 ( .A(n356), .B(n355), .ZN(n362) );
  XOR2_X1 U430 ( .A(n358), .B(n357), .Z(n360) );
  NAND2_X1 U431 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U432 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U433 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U434 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n366), .B(n365), .ZN(n555) );
  INV_X1 U436 ( .A(n555), .ZN(n577) );
  XOR2_X1 U437 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n368) );
  NAND2_X1 U438 ( .A1(G230GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U439 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U440 ( .A(n369), .B(KEYINPUT76), .Z(n373) );
  XNOR2_X1 U441 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U442 ( .A(n373), .B(n372), .ZN(n378) );
  XOR2_X1 U443 ( .A(G120GAT), .B(G71GAT), .Z(n433) );
  XOR2_X1 U444 ( .A(G64GAT), .B(G176GAT), .Z(n395) );
  XNOR2_X1 U445 ( .A(n433), .B(n395), .ZN(n376) );
  XOR2_X1 U446 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n375) );
  XNOR2_X1 U447 ( .A(G204GAT), .B(KEYINPUT72), .ZN(n374) );
  XNOR2_X1 U448 ( .A(n380), .B(n379), .ZN(n582) );
  INV_X1 U449 ( .A(n557), .ZN(n567) );
  NOR2_X1 U450 ( .A1(n577), .A2(n567), .ZN(n382) );
  XNOR2_X1 U451 ( .A(KEYINPUT116), .B(KEYINPUT46), .ZN(n381) );
  XNOR2_X1 U452 ( .A(n382), .B(n381), .ZN(n383) );
  NOR2_X1 U453 ( .A1(n562), .A2(n383), .ZN(n384) );
  NAND2_X1 U454 ( .A1(n573), .A2(n384), .ZN(n385) );
  XNOR2_X1 U455 ( .A(KEYINPUT47), .B(n385), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n386), .B(KEYINPUT117), .ZN(n391) );
  XOR2_X1 U457 ( .A(KEYINPUT36), .B(n495), .Z(n590) );
  NAND2_X1 U458 ( .A1(n590), .A2(n586), .ZN(n387) );
  NAND2_X1 U459 ( .A1(n389), .A2(n577), .ZN(n390) );
  NAND2_X1 U460 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X1 U461 ( .A(KEYINPUT48), .B(n392), .ZN(n456) );
  XOR2_X1 U462 ( .A(G169GAT), .B(KEYINPUT19), .Z(n394) );
  XNOR2_X1 U463 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n394), .B(n393), .ZN(n434) );
  XOR2_X1 U465 ( .A(n395), .B(G92GAT), .Z(n397) );
  NAND2_X1 U466 ( .A1(G226GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U467 ( .A(n397), .B(n396), .ZN(n399) );
  XOR2_X1 U468 ( .A(n399), .B(n398), .Z(n403) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U471 ( .A(n434), .B(n404), .ZN(n540) );
  XOR2_X1 U472 ( .A(n540), .B(KEYINPUT27), .Z(n467) );
  XOR2_X1 U473 ( .A(KEYINPUT6), .B(KEYINPUT89), .Z(n406) );
  XNOR2_X1 U474 ( .A(KEYINPUT93), .B(KEYINPUT95), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U476 ( .A(KEYINPUT90), .B(G57GAT), .Z(n408) );
  XNOR2_X1 U477 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n407) );
  XNOR2_X1 U478 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U479 ( .A(n410), .B(n409), .Z(n415) );
  XOR2_X1 U480 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n412) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U482 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U483 ( .A(KEYINPUT91), .B(n413), .ZN(n414) );
  XNOR2_X1 U484 ( .A(n415), .B(n414), .ZN(n428) );
  XOR2_X1 U485 ( .A(G148GAT), .B(G85GAT), .Z(n417) );
  XNOR2_X1 U486 ( .A(G29GAT), .B(G162GAT), .ZN(n416) );
  XNOR2_X1 U487 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U488 ( .A(KEYINPUT94), .B(G127GAT), .Z(n419) );
  XNOR2_X1 U489 ( .A(G155GAT), .B(G120GAT), .ZN(n418) );
  XNOR2_X1 U490 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U491 ( .A(n421), .B(n420), .Z(n426) );
  XOR2_X1 U492 ( .A(G113GAT), .B(KEYINPUT82), .Z(n423) );
  XNOR2_X1 U493 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n422) );
  XNOR2_X1 U494 ( .A(n423), .B(n422), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n424), .B(n438), .ZN(n425) );
  XNOR2_X1 U496 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U497 ( .A(n428), .B(n427), .ZN(n501) );
  XNOR2_X1 U498 ( .A(G1GAT), .B(n501), .ZN(n522) );
  NAND2_X1 U499 ( .A1(n467), .A2(n522), .ZN(n429) );
  XOR2_X1 U500 ( .A(n429), .B(KEYINPUT96), .Z(n476) );
  NAND2_X1 U501 ( .A1(n456), .A2(n476), .ZN(n430) );
  XNOR2_X1 U502 ( .A(KEYINPUT118), .B(n430), .ZN(n553) );
  NOR2_X1 U503 ( .A1(n530), .A2(n553), .ZN(n447) );
  XOR2_X1 U504 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n432) );
  XNOR2_X1 U505 ( .A(G99GAT), .B(KEYINPUT84), .ZN(n431) );
  XNOR2_X1 U506 ( .A(n432), .B(n431), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n434), .B(n433), .ZN(n437) );
  AND2_X1 U508 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XOR2_X1 U509 ( .A(n438), .B(G183GAT), .Z(n439) );
  XNOR2_X1 U510 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U511 ( .A(G43GAT), .B(G190GAT), .Z(n441) );
  XOR2_X1 U512 ( .A(n446), .B(n445), .Z(n542) );
  INV_X1 U513 ( .A(n542), .ZN(n528) );
  NAND2_X1 U514 ( .A1(n447), .A2(n528), .ZN(n448) );
  NAND2_X1 U515 ( .A1(n550), .A2(n586), .ZN(n452) );
  XOR2_X1 U516 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n450) );
  XNOR2_X1 U517 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n449) );
  XNOR2_X1 U518 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U519 ( .A(n452), .B(n451), .ZN(G1342GAT) );
  NAND2_X1 U520 ( .A1(n550), .A2(n562), .ZN(n455) );
  XOR2_X1 U521 ( .A(KEYINPUT51), .B(KEYINPUT122), .Z(n453) );
  XNOR2_X1 U522 ( .A(n455), .B(n454), .ZN(G1343GAT) );
  XOR2_X1 U523 ( .A(KEYINPUT54), .B(KEYINPUT124), .Z(n458) );
  INV_X1 U524 ( .A(n540), .ZN(n525) );
  NAND2_X1 U525 ( .A1(n456), .A2(n525), .ZN(n457) );
  XOR2_X1 U526 ( .A(n458), .B(n457), .Z(n459) );
  NAND2_X1 U527 ( .A1(n468), .A2(n576), .ZN(n460) );
  XNOR2_X1 U528 ( .A(n460), .B(KEYINPUT55), .ZN(n461) );
  NAND2_X1 U529 ( .A1(n461), .A2(n528), .ZN(n572) );
  NOR2_X1 U530 ( .A1(n495), .A2(n572), .ZN(n464) );
  XOR2_X1 U531 ( .A(KEYINPUT107), .B(KEYINPUT38), .Z(n486) );
  XNOR2_X1 U532 ( .A(n466), .B(n465), .ZN(n554) );
  INV_X1 U533 ( .A(n554), .ZN(n575) );
  NAND2_X1 U534 ( .A1(n575), .A2(n467), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n528), .A2(n525), .ZN(n469) );
  NAND2_X1 U536 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U537 ( .A(n470), .B(KEYINPUT97), .ZN(n471) );
  XNOR2_X1 U538 ( .A(n471), .B(KEYINPUT25), .ZN(n472) );
  NAND2_X1 U539 ( .A1(n473), .A2(n472), .ZN(n474) );
  INV_X1 U540 ( .A(n522), .ZN(n538) );
  NAND2_X1 U541 ( .A1(n474), .A2(n538), .ZN(n475) );
  XNOR2_X1 U542 ( .A(n475), .B(KEYINPUT98), .ZN(n479) );
  INV_X1 U543 ( .A(n530), .ZN(n545) );
  AND2_X1 U544 ( .A1(n476), .A2(n545), .ZN(n477) );
  NAND2_X1 U545 ( .A1(n477), .A2(n542), .ZN(n478) );
  NAND2_X1 U546 ( .A1(n479), .A2(n478), .ZN(n481) );
  NAND2_X1 U547 ( .A1(n498), .A2(n573), .ZN(n482) );
  XNOR2_X1 U548 ( .A(n482), .B(KEYINPUT105), .ZN(n483) );
  NAND2_X1 U549 ( .A1(n483), .A2(n590), .ZN(n484) );
  XNOR2_X1 U550 ( .A(n484), .B(KEYINPUT37), .ZN(n537) );
  NOR2_X1 U551 ( .A1(n577), .A2(n582), .ZN(n500) );
  NAND2_X1 U552 ( .A1(n537), .A2(n500), .ZN(n485) );
  XNOR2_X1 U553 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U554 ( .A(KEYINPUT106), .B(n487), .Z(n518) );
  NAND2_X1 U555 ( .A1(n518), .A2(n522), .ZN(n490) );
  XOR2_X1 U556 ( .A(KEYINPUT39), .B(KEYINPUT108), .Z(n488) );
  XNOR2_X1 U557 ( .A(n488), .B(G29GAT), .ZN(n489) );
  XNOR2_X1 U558 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n518), .A2(n528), .ZN(n494) );
  XOR2_X1 U560 ( .A(KEYINPUT40), .B(KEYINPUT110), .Z(n492) );
  NAND2_X1 U561 ( .A1(n586), .A2(n495), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n496), .B(KEYINPUT81), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n497), .B(KEYINPUT16), .ZN(n499) );
  AND2_X1 U564 ( .A1(n499), .A2(n498), .ZN(n521) );
  NAND2_X1 U565 ( .A1(n500), .A2(n521), .ZN(n508) );
  AND2_X1 U566 ( .A1(n508), .A2(G1GAT), .ZN(n503) );
  NOR2_X1 U567 ( .A1(n508), .A2(n501), .ZN(n502) );
  NOR2_X1 U568 ( .A1(n503), .A2(n502), .ZN(n507) );
  XOR2_X1 U569 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n505) );
  XNOR2_X1 U570 ( .A(KEYINPUT101), .B(KEYINPUT100), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U572 ( .A(n507), .B(n506), .Z(G1324GAT) );
  XOR2_X1 U573 ( .A(G8GAT), .B(KEYINPUT103), .Z(n510) );
  INV_X1 U574 ( .A(n508), .ZN(n513) );
  NAND2_X1 U575 ( .A1(n513), .A2(n525), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1325GAT) );
  XOR2_X1 U577 ( .A(G15GAT), .B(KEYINPUT35), .Z(n512) );
  NAND2_X1 U578 ( .A1(n513), .A2(n528), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(G1326GAT) );
  NAND2_X1 U580 ( .A1(n513), .A2(n530), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(KEYINPUT104), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G22GAT), .B(n515), .ZN(G1327GAT) );
  XOR2_X1 U583 ( .A(G36GAT), .B(KEYINPUT109), .Z(n517) );
  NAND2_X1 U584 ( .A1(n518), .A2(n525), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1329GAT) );
  NAND2_X1 U586 ( .A1(n518), .A2(n530), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n519), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U588 ( .A1(n555), .A2(n567), .ZN(n520) );
  XOR2_X1 U589 ( .A(KEYINPUT111), .B(n520), .Z(n536) );
  AND2_X1 U590 ( .A1(n536), .A2(n521), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n522), .A2(n531), .ZN(n523) );
  XNOR2_X1 U592 ( .A(KEYINPUT42), .B(n523), .ZN(n524) );
  XNOR2_X1 U593 ( .A(G57GAT), .B(n524), .ZN(G1332GAT) );
  NAND2_X1 U594 ( .A1(n531), .A2(n525), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n526), .B(KEYINPUT112), .ZN(n527) );
  XNOR2_X1 U596 ( .A(G64GAT), .B(n527), .ZN(G1333GAT) );
  NAND2_X1 U597 ( .A1(n528), .A2(n531), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n529), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT114), .B(KEYINPUT43), .Z(n533) );
  NAND2_X1 U600 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n535) );
  XOR2_X1 U602 ( .A(G78GAT), .B(KEYINPUT113), .Z(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(G1335GAT) );
  NAND2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n544) );
  NOR2_X1 U605 ( .A1(n538), .A2(n544), .ZN(n539) );
  XOR2_X1 U606 ( .A(G85GAT), .B(n539), .Z(G1336GAT) );
  NOR2_X1 U607 ( .A1(n540), .A2(n544), .ZN(n541) );
  XOR2_X1 U608 ( .A(G92GAT), .B(n541), .Z(G1337GAT) );
  NOR2_X1 U609 ( .A1(n542), .A2(n544), .ZN(n543) );
  XOR2_X1 U610 ( .A(G99GAT), .B(n543), .Z(G1338GAT) );
  NOR2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n547) );
  XNOR2_X1 U612 ( .A(KEYINPUT115), .B(KEYINPUT44), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G106GAT), .B(n548), .ZN(G1339GAT) );
  NAND2_X1 U615 ( .A1(n555), .A2(n550), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U617 ( .A(G120GAT), .B(KEYINPUT49), .Z(n552) );
  NAND2_X1 U618 ( .A1(n550), .A2(n557), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1341GAT) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n563), .A2(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  NAND2_X1 U624 ( .A1(n563), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n586), .A2(n563), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U629 ( .A(G162GAT), .B(KEYINPUT123), .Z(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1347GAT) );
  NOR2_X1 U632 ( .A1(n577), .A2(n572), .ZN(n566) );
  XOR2_X1 U633 ( .A(G169GAT), .B(n566), .Z(G1348GAT) );
  NOR2_X1 U634 ( .A1(n572), .A2(n567), .ZN(n571) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT57), .Z(n569) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(G183GAT), .B(n574), .Z(G1350GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n581) );
  NOR2_X1 U642 ( .A1(n577), .A2(n581), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n584) );
  INV_X1 U647 ( .A(n581), .ZN(n589) );
  NAND2_X1 U648 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(n585), .ZN(G1353GAT) );
  XOR2_X1 U651 ( .A(G211GAT), .B(KEYINPUT127), .Z(n588) );
  NAND2_X1 U652 ( .A1(n589), .A2(n586), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1354GAT) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

