

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XOR2_X1 U323 ( .A(n386), .B(n385), .Z(n291) );
  XNOR2_X1 U324 ( .A(n416), .B(KEYINPUT113), .ZN(n417) );
  XNOR2_X1 U325 ( .A(n418), .B(n417), .ZN(n421) );
  XNOR2_X1 U326 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n429) );
  XNOR2_X1 U327 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n426) );
  XNOR2_X1 U328 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U329 ( .A(n427), .B(n426), .ZN(n528) );
  XNOR2_X1 U330 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U331 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n450) );
  XNOR2_X1 U332 ( .A(n393), .B(n392), .ZN(n456) );
  XNOR2_X1 U333 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U334 ( .A(n307), .B(n338), .Z(n522) );
  XNOR2_X1 U335 ( .A(n453), .B(G176GAT), .ZN(n454) );
  XNOR2_X1 U336 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  XOR2_X1 U337 ( .A(G120GAT), .B(G71GAT), .Z(n389) );
  XOR2_X1 U338 ( .A(G15GAT), .B(G127GAT), .Z(n353) );
  XOR2_X1 U339 ( .A(n389), .B(n353), .Z(n293) );
  NAND2_X1 U340 ( .A1(G227GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U341 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U342 ( .A(G113GAT), .B(KEYINPUT0), .Z(n310) );
  XOR2_X1 U343 ( .A(n294), .B(n310), .Z(n302) );
  XOR2_X1 U344 ( .A(G190GAT), .B(G134GAT), .Z(n296) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(G99GAT), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U347 ( .A(G176GAT), .B(G183GAT), .Z(n298) );
  XNOR2_X1 U348 ( .A(KEYINPUT82), .B(KEYINPUT20), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n307) );
  XOR2_X1 U352 ( .A(KEYINPUT81), .B(KEYINPUT19), .Z(n304) );
  XNOR2_X1 U353 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n306) );
  XOR2_X1 U355 ( .A(KEYINPUT80), .B(KEYINPUT18), .Z(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n338) );
  INV_X1 U357 ( .A(n522), .ZN(n531) );
  XOR2_X1 U358 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n309) );
  XNOR2_X1 U359 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n314) );
  XOR2_X1 U361 ( .A(G134GAT), .B(KEYINPUT76), .Z(n369) );
  XOR2_X1 U362 ( .A(G85GAT), .B(n369), .Z(n312) );
  XNOR2_X1 U363 ( .A(n310), .B(G162GAT), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U365 ( .A(n314), .B(n313), .Z(n316) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U368 ( .A(n317), .B(KEYINPUT90), .Z(n321) );
  XOR2_X1 U369 ( .A(G155GAT), .B(KEYINPUT2), .Z(n319) );
  XNOR2_X1 U370 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n446) );
  XNOR2_X1 U372 ( .A(n446), .B(KEYINPUT87), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n329) );
  XOR2_X1 U374 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n323) );
  XNOR2_X1 U375 ( .A(G1GAT), .B(G57GAT), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U377 ( .A(G148GAT), .B(G127GAT), .Z(n325) );
  XNOR2_X1 U378 ( .A(G29GAT), .B(G120GAT), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U380 ( .A(n327), .B(n326), .Z(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n542) );
  XNOR2_X1 U382 ( .A(G8GAT), .B(G183GAT), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n330), .B(KEYINPUT78), .ZN(n352) );
  XOR2_X1 U384 ( .A(G176GAT), .B(G64GAT), .Z(n387) );
  XOR2_X1 U385 ( .A(n352), .B(n387), .Z(n332) );
  NAND2_X1 U386 ( .A1(G226GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n345) );
  XOR2_X1 U388 ( .A(KEYINPUT92), .B(KEYINPUT94), .Z(n334) );
  XNOR2_X1 U389 ( .A(KEYINPUT91), .B(KEYINPUT93), .ZN(n333) );
  XNOR2_X1 U390 ( .A(n334), .B(n333), .ZN(n337) );
  XOR2_X1 U391 ( .A(G92GAT), .B(G218GAT), .Z(n336) );
  XNOR2_X1 U392 ( .A(G36GAT), .B(G190GAT), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n368) );
  XOR2_X1 U394 ( .A(n337), .B(n368), .Z(n343) );
  INV_X1 U395 ( .A(n338), .ZN(n341) );
  XOR2_X1 U396 ( .A(G204GAT), .B(G211GAT), .Z(n340) );
  XNOR2_X1 U397 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n439) );
  XNOR2_X1 U399 ( .A(n341), .B(n439), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n520) );
  XOR2_X1 U402 ( .A(KEYINPUT119), .B(n520), .Z(n428) );
  XOR2_X1 U403 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n347) );
  NAND2_X1 U404 ( .A1(G231GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U406 ( .A(KEYINPUT14), .B(n348), .ZN(n360) );
  XOR2_X1 U407 ( .A(KEYINPUT79), .B(G64GAT), .Z(n350) );
  XNOR2_X1 U408 ( .A(G71GAT), .B(G155GAT), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U410 ( .A(n352), .B(n351), .Z(n355) );
  XOR2_X1 U411 ( .A(G57GAT), .B(KEYINPUT13), .Z(n388) );
  XNOR2_X1 U412 ( .A(n353), .B(n388), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U414 ( .A(n356), .B(G211GAT), .Z(n358) );
  XOR2_X1 U415 ( .A(G22GAT), .B(G1GAT), .Z(n394) );
  XNOR2_X1 U416 ( .A(n394), .B(G78GAT), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n484) );
  XOR2_X1 U419 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n362) );
  XNOR2_X1 U420 ( .A(KEYINPUT9), .B(KEYINPUT75), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n373) );
  XNOR2_X1 U422 ( .A(G99GAT), .B(G106GAT), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n363), .B(G85GAT), .ZN(n384) );
  INV_X1 U424 ( .A(KEYINPUT74), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n384), .B(n364), .ZN(n366) );
  NAND2_X1 U426 ( .A1(G232GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U428 ( .A(n368), .B(n367), .Z(n371) );
  XOR2_X1 U429 ( .A(G50GAT), .B(G162GAT), .Z(n435) );
  XNOR2_X1 U430 ( .A(n435), .B(n369), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n373), .B(n372), .ZN(n378) );
  XNOR2_X1 U433 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n374), .B(G29GAT), .ZN(n375) );
  XOR2_X1 U435 ( .A(n375), .B(KEYINPUT8), .Z(n377) );
  XNOR2_X1 U436 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n406) );
  XNOR2_X1 U438 ( .A(n378), .B(n406), .ZN(n419) );
  XNOR2_X1 U439 ( .A(KEYINPUT77), .B(n419), .ZN(n559) );
  XOR2_X1 U440 ( .A(KEYINPUT36), .B(n559), .Z(n581) );
  NOR2_X1 U441 ( .A1(n484), .A2(n581), .ZN(n379) );
  XNOR2_X1 U442 ( .A(n379), .B(KEYINPUT45), .ZN(n414) );
  XNOR2_X1 U443 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n381) );
  AND2_X1 U444 ( .A1(G230GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U446 ( .A(n382), .B(KEYINPUT31), .Z(n386) );
  XNOR2_X1 U447 ( .A(G78GAT), .B(KEYINPUT73), .ZN(n383) );
  XNOR2_X1 U448 ( .A(n383), .B(G148GAT), .ZN(n447) );
  XNOR2_X1 U449 ( .A(n447), .B(n384), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n291), .B(n387), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n391) );
  XNOR2_X1 U452 ( .A(G204GAT), .B(G92GAT), .ZN(n390) );
  INV_X1 U453 ( .A(n456), .ZN(n573) );
  XOR2_X1 U454 ( .A(G36GAT), .B(G50GAT), .Z(n396) );
  XNOR2_X1 U455 ( .A(n394), .B(KEYINPUT30), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n410) );
  XOR2_X1 U457 ( .A(G113GAT), .B(G141GAT), .Z(n398) );
  XNOR2_X1 U458 ( .A(G169GAT), .B(G197GAT), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U460 ( .A(KEYINPUT71), .B(KEYINPUT66), .Z(n400) );
  XNOR2_X1 U461 ( .A(G15GAT), .B(G8GAT), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U463 ( .A(n402), .B(n401), .Z(n408) );
  XOR2_X1 U464 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n404) );
  XNOR2_X1 U465 ( .A(KEYINPUT68), .B(KEYINPUT72), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U469 ( .A(n410), .B(n409), .Z(n412) );
  NAND2_X1 U470 ( .A1(G229GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n566) );
  INV_X1 U472 ( .A(n566), .ZN(n504) );
  NOR2_X1 U473 ( .A1(n573), .A2(n566), .ZN(n413) );
  NAND2_X1 U474 ( .A1(n414), .A2(n413), .ZN(n425) );
  XNOR2_X1 U475 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n415), .B(n573), .ZN(n547) );
  NAND2_X1 U477 ( .A1(n547), .A2(n566), .ZN(n418) );
  INV_X1 U478 ( .A(KEYINPUT46), .ZN(n416) );
  INV_X1 U479 ( .A(n419), .ZN(n553) );
  INV_X1 U480 ( .A(n484), .ZN(n576) );
  NOR2_X1 U481 ( .A1(n553), .A2(n576), .ZN(n420) );
  NAND2_X1 U482 ( .A1(n421), .A2(n420), .ZN(n423) );
  XOR2_X1 U483 ( .A(KEYINPUT114), .B(KEYINPUT47), .Z(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n424) );
  NAND2_X1 U485 ( .A1(n425), .A2(n424), .ZN(n427) );
  NAND2_X1 U486 ( .A1(n428), .A2(n528), .ZN(n430) );
  NOR2_X1 U487 ( .A1(n542), .A2(n431), .ZN(n565) );
  XOR2_X1 U488 ( .A(KEYINPUT84), .B(G106GAT), .Z(n433) );
  XNOR2_X1 U489 ( .A(G22GAT), .B(G218GAT), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U491 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U492 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U494 ( .A(n438), .B(KEYINPUT22), .Z(n441) );
  XNOR2_X1 U495 ( .A(n439), .B(KEYINPUT85), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U497 ( .A(KEYINPUT83), .B(KEYINPUT23), .Z(n443) );
  XNOR2_X1 U498 ( .A(KEYINPUT24), .B(KEYINPUT86), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U500 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n463) );
  NAND2_X1 U503 ( .A1(n565), .A2(n463), .ZN(n451) );
  NOR2_X1 U504 ( .A1(n531), .A2(n452), .ZN(n560) );
  NAND2_X1 U505 ( .A1(n560), .A2(n547), .ZN(n455) );
  XOR2_X1 U506 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n453) );
  XOR2_X1 U507 ( .A(KEYINPUT98), .B(KEYINPUT34), .Z(n474) );
  NAND2_X1 U508 ( .A1(n566), .A2(n456), .ZN(n489) );
  NOR2_X1 U509 ( .A1(n484), .A2(n559), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n457), .B(KEYINPUT16), .ZN(n471) );
  XOR2_X1 U511 ( .A(n463), .B(KEYINPUT28), .Z(n524) );
  XOR2_X1 U512 ( .A(n520), .B(KEYINPUT95), .Z(n458) );
  XNOR2_X1 U513 ( .A(n458), .B(KEYINPUT27), .ZN(n465) );
  NAND2_X1 U514 ( .A1(n465), .A2(n542), .ZN(n459) );
  NOR2_X1 U515 ( .A1(n524), .A2(n459), .ZN(n529) );
  NAND2_X1 U516 ( .A1(n531), .A2(n529), .ZN(n470) );
  INV_X1 U517 ( .A(n542), .ZN(n468) );
  NAND2_X1 U518 ( .A1(n522), .A2(n520), .ZN(n460) );
  NAND2_X1 U519 ( .A1(n460), .A2(n463), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(KEYINPUT96), .ZN(n462) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(n462), .Z(n466) );
  NOR2_X1 U522 ( .A1(n522), .A2(n463), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n464), .B(KEYINPUT26), .ZN(n564) );
  NAND2_X1 U524 ( .A1(n465), .A2(n564), .ZN(n544) );
  NAND2_X1 U525 ( .A1(n466), .A2(n544), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U527 ( .A1(n470), .A2(n469), .ZN(n483) );
  NAND2_X1 U528 ( .A1(n471), .A2(n483), .ZN(n505) );
  NOR2_X1 U529 ( .A1(n489), .A2(n505), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT97), .B(n472), .Z(n479) );
  NAND2_X1 U531 ( .A1(n479), .A2(n542), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U533 ( .A(G1GAT), .B(n475), .Z(G1324GAT) );
  NAND2_X1 U534 ( .A1(n520), .A2(n479), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U537 ( .A1(n479), .A2(n522), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n481) );
  NAND2_X1 U540 ( .A1(n479), .A2(n524), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  XOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  NAND2_X1 U544 ( .A1(n484), .A2(n483), .ZN(n485) );
  NOR2_X1 U545 ( .A1(n581), .A2(n485), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT102), .B(KEYINPUT37), .Z(n486) );
  XNOR2_X1 U547 ( .A(KEYINPUT101), .B(n486), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n517) );
  NOR2_X1 U549 ( .A1(n517), .A2(n489), .ZN(n490) );
  XOR2_X1 U550 ( .A(KEYINPUT38), .B(n490), .Z(n491) );
  XNOR2_X1 U551 ( .A(KEYINPUT103), .B(n491), .ZN(n499) );
  NAND2_X1 U552 ( .A1(n499), .A2(n542), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n495) );
  NAND2_X1 U555 ( .A1(n499), .A2(n520), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  NAND2_X1 U558 ( .A1(n499), .A2(n522), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U561 ( .A1(n499), .A2(n524), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT106), .ZN(n501) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(KEYINPUT108), .ZN(n503) );
  XOR2_X1 U566 ( .A(KEYINPUT107), .B(n503), .Z(n507) );
  NAND2_X1 U567 ( .A1(n504), .A2(n547), .ZN(n516) );
  NOR2_X1 U568 ( .A1(n505), .A2(n516), .ZN(n512) );
  NAND2_X1 U569 ( .A1(n512), .A2(n542), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  XOR2_X1 U571 ( .A(G64GAT), .B(KEYINPUT109), .Z(n509) );
  NAND2_X1 U572 ( .A1(n512), .A2(n520), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n522), .A2(n512), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(KEYINPUT110), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n511), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n514) );
  NAND2_X1 U578 ( .A1(n512), .A2(n524), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U580 ( .A(G78GAT), .B(n515), .Z(G1335GAT) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n519) );
  NOR2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n525), .A2(n542), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n520), .A2(n525), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n525), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  XOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT115), .Z(n533) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n538), .A2(n566), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U598 ( .A1(n538), .A2(n547), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NAND2_X1 U600 ( .A1(n576), .A2(n538), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n540) );
  NAND2_X1 U604 ( .A1(n538), .A2(n559), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(n541), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n542), .A2(n528), .ZN(n543) );
  NOR2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U609 ( .A(KEYINPUT117), .B(n545), .Z(n552) );
  NAND2_X1 U610 ( .A1(n552), .A2(n566), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  NAND2_X1 U613 ( .A1(n552), .A2(n547), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  NAND2_X1 U616 ( .A1(n576), .A2(n552), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT118), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n555), .ZN(G1347GAT) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n566), .A2(n560), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n576), .A2(n560), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n562) );
  XOR2_X1 U627 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n580) );
  INV_X1 U632 ( .A(n580), .ZN(n577) );
  NAND2_X1 U633 ( .A1(n577), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n571) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(n572), .Z(n575) );
  NAND2_X1 U640 ( .A1(n577), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(n582), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

