

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U555 ( .A(n702), .ZN(n719) );
  NOR2_X2 U556 ( .A1(n560), .A2(n559), .ZN(G164) );
  NOR2_X1 U557 ( .A1(n810), .A2(n809), .ZN(n811) );
  BUF_X1 U558 ( .A(n702), .Z(n740) );
  BUF_X1 U559 ( .A(n887), .Z(n521) );
  XNOR2_X1 U560 ( .A(n540), .B(KEYINPUT65), .ZN(n887) );
  XNOR2_X1 U561 ( .A(n730), .B(n729), .ZN(n738) );
  INV_X1 U562 ( .A(G8), .ZN(n690) );
  NOR2_X1 U563 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U564 ( .A1(G168), .A2(n695), .ZN(n696) );
  INV_X1 U565 ( .A(KEYINPUT29), .ZN(n729) );
  OR2_X1 U566 ( .A1(n732), .A2(n746), .ZN(n736) );
  NAND2_X1 U567 ( .A1(n779), .A2(n681), .ZN(n702) );
  NAND2_X1 U568 ( .A1(G8), .A2(n702), .ZN(n774) );
  NOR2_X1 U569 ( .A1(n635), .A2(n527), .ZN(n640) );
  NOR2_X1 U570 ( .A1(n635), .A2(G651), .ZN(n651) );
  NOR2_X1 U571 ( .A1(n580), .A2(n579), .ZN(n974) );
  NOR2_X1 U572 ( .A1(n545), .A2(n544), .ZN(G160) );
  NOR2_X1 U573 ( .A1(G543), .A2(G651), .ZN(n642) );
  NAND2_X1 U574 ( .A1(G89), .A2(n642), .ZN(n522) );
  XOR2_X1 U575 ( .A(KEYINPUT4), .B(n522), .Z(n523) );
  XNOR2_X1 U576 ( .A(n523), .B(KEYINPUT69), .ZN(n525) );
  XOR2_X1 U577 ( .A(KEYINPUT0), .B(G543), .Z(n635) );
  INV_X1 U578 ( .A(G651), .ZN(n527) );
  NAND2_X1 U579 ( .A1(G76), .A2(n640), .ZN(n524) );
  NAND2_X1 U580 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U581 ( .A(n526), .B(KEYINPUT5), .ZN(n533) );
  NOR2_X1 U582 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n528), .Z(n644) );
  NAND2_X1 U584 ( .A1(G63), .A2(n644), .ZN(n530) );
  NAND2_X1 U585 ( .A1(G51), .A2(n651), .ZN(n529) );
  NAND2_X1 U586 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U587 ( .A(KEYINPUT6), .B(n531), .Z(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U589 ( .A(n534), .B(KEYINPUT7), .ZN(G168) );
  INV_X1 U590 ( .A(G2104), .ZN(n541) );
  NOR2_X4 U591 ( .A1(G2105), .A2(n541), .ZN(n883) );
  NAND2_X1 U592 ( .A1(G101), .A2(n883), .ZN(n535) );
  XOR2_X1 U593 ( .A(KEYINPUT23), .B(n535), .Z(n536) );
  XNOR2_X1 U594 ( .A(n536), .B(KEYINPUT64), .ZN(n539) );
  NOR2_X1 U595 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  XOR2_X2 U596 ( .A(KEYINPUT17), .B(n537), .Z(n884) );
  NAND2_X1 U597 ( .A1(G137), .A2(n884), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n539), .A2(n538), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G2105), .A2(G2104), .ZN(n540) );
  NAND2_X1 U600 ( .A1(G113), .A2(n521), .ZN(n543) );
  AND2_X1 U601 ( .A1(n541), .A2(G2105), .ZN(n888) );
  NAND2_X1 U602 ( .A1(G125), .A2(n888), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U604 ( .A1(G85), .A2(n642), .ZN(n547) );
  NAND2_X1 U605 ( .A1(G72), .A2(n640), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U607 ( .A1(G60), .A2(n644), .ZN(n549) );
  NAND2_X1 U608 ( .A1(G47), .A2(n651), .ZN(n548) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n550) );
  OR2_X1 U610 ( .A1(n551), .A2(n550), .ZN(G290) );
  NAND2_X1 U611 ( .A1(n887), .A2(G114), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n552), .B(KEYINPUT82), .ZN(n554) );
  NAND2_X1 U613 ( .A1(G126), .A2(n888), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U615 ( .A(n555), .B(KEYINPUT83), .ZN(n557) );
  NAND2_X1 U616 ( .A1(G138), .A2(n884), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U618 ( .A1(G102), .A2(n883), .ZN(n558) );
  XOR2_X1 U619 ( .A(KEYINPUT84), .B(n558), .Z(n559) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  INV_X1 U622 ( .A(G132), .ZN(G219) );
  INV_X1 U623 ( .A(G82), .ZN(G220) );
  NAND2_X1 U624 ( .A1(G64), .A2(n644), .ZN(n562) );
  NAND2_X1 U625 ( .A1(G52), .A2(n651), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n567) );
  NAND2_X1 U627 ( .A1(G90), .A2(n642), .ZN(n564) );
  NAND2_X1 U628 ( .A1(G77), .A2(n640), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  NOR2_X1 U631 ( .A1(n567), .A2(n566), .ZN(G171) );
  XOR2_X1 U632 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U633 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n569) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G223) );
  INV_X1 U636 ( .A(G223), .ZN(n827) );
  NAND2_X1 U637 ( .A1(n827), .A2(G567), .ZN(n570) );
  XOR2_X1 U638 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  XOR2_X1 U639 ( .A(KEYINPUT68), .B(KEYINPUT14), .Z(n572) );
  NAND2_X1 U640 ( .A1(G56), .A2(n644), .ZN(n571) );
  XNOR2_X1 U641 ( .A(n572), .B(n571), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G68), .A2(n640), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n642), .A2(G81), .ZN(n573) );
  XNOR2_X1 U644 ( .A(n573), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U646 ( .A(n576), .B(KEYINPUT13), .ZN(n578) );
  NAND2_X1 U647 ( .A1(G43), .A2(n651), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n974), .A2(G860), .ZN(G153) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U652 ( .A1(G66), .A2(n644), .ZN(n582) );
  NAND2_X1 U653 ( .A1(G92), .A2(n642), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U655 ( .A1(G79), .A2(n640), .ZN(n584) );
  NAND2_X1 U656 ( .A1(G54), .A2(n651), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U659 ( .A(KEYINPUT15), .B(n587), .Z(n910) );
  INV_X1 U660 ( .A(n910), .ZN(n989) );
  INV_X1 U661 ( .A(G868), .ZN(n602) );
  NAND2_X1 U662 ( .A1(n989), .A2(n602), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G91), .A2(n642), .ZN(n591) );
  NAND2_X1 U665 ( .A1(G78), .A2(n640), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n644), .A2(G65), .ZN(n592) );
  XOR2_X1 U668 ( .A(KEYINPUT66), .B(n592), .Z(n593) );
  NOR2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n651), .A2(G53), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(G299) );
  NOR2_X1 U672 ( .A1(G286), .A2(n602), .ZN(n598) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U674 ( .A1(n598), .A2(n597), .ZN(G297) );
  INV_X1 U675 ( .A(G860), .ZN(n617) );
  NAND2_X1 U676 ( .A1(n617), .A2(G559), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n599), .A2(n910), .ZN(n600) );
  XNOR2_X1 U678 ( .A(n600), .B(KEYINPUT16), .ZN(n601) );
  XNOR2_X1 U679 ( .A(KEYINPUT70), .B(n601), .ZN(G148) );
  NAND2_X1 U680 ( .A1(n974), .A2(n602), .ZN(n603) );
  XNOR2_X1 U681 ( .A(KEYINPUT71), .B(n603), .ZN(n606) );
  NAND2_X1 U682 ( .A1(G868), .A2(n910), .ZN(n604) );
  NOR2_X1 U683 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U684 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G123), .A2(n888), .ZN(n607) );
  XNOR2_X1 U686 ( .A(n607), .B(KEYINPUT18), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n521), .A2(G111), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G99), .A2(n883), .ZN(n611) );
  NAND2_X1 U690 ( .A1(G135), .A2(n884), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n933) );
  XNOR2_X1 U693 ( .A(G2096), .B(n933), .ZN(n615) );
  INV_X1 U694 ( .A(G2100), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U696 ( .A1(G559), .A2(n910), .ZN(n616) );
  XNOR2_X1 U697 ( .A(n616), .B(n974), .ZN(n660) );
  NAND2_X1 U698 ( .A1(n617), .A2(n660), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G93), .A2(n642), .ZN(n619) );
  NAND2_X1 U700 ( .A1(G80), .A2(n640), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G55), .A2(n651), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n620), .B(KEYINPUT72), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n644), .A2(G67), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n663) );
  XOR2_X1 U707 ( .A(n625), .B(n663), .Z(G145) );
  NAND2_X1 U708 ( .A1(G88), .A2(n642), .ZN(n627) );
  NAND2_X1 U709 ( .A1(G75), .A2(n640), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G62), .A2(n644), .ZN(n629) );
  NAND2_X1 U712 ( .A1(G50), .A2(n651), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U714 ( .A1(n631), .A2(n630), .ZN(G166) );
  NAND2_X1 U715 ( .A1(G49), .A2(n651), .ZN(n633) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U718 ( .A(n634), .B(KEYINPUT73), .ZN(n637) );
  NAND2_X1 U719 ( .A1(G87), .A2(n635), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U721 ( .A1(n644), .A2(n638), .ZN(n639) );
  XOR2_X1 U722 ( .A(KEYINPUT74), .B(n639), .Z(G288) );
  NAND2_X1 U723 ( .A1(n640), .A2(G73), .ZN(n641) );
  XNOR2_X1 U724 ( .A(KEYINPUT2), .B(n641), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n642), .A2(G86), .ZN(n643) );
  XOR2_X1 U726 ( .A(KEYINPUT75), .B(n643), .Z(n646) );
  NAND2_X1 U727 ( .A1(n644), .A2(G61), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U729 ( .A(KEYINPUT76), .B(n647), .Z(n648) );
  NAND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n650), .B(KEYINPUT77), .ZN(n653) );
  NAND2_X1 U732 ( .A1(G48), .A2(n651), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(G305) );
  XNOR2_X1 U734 ( .A(G166), .B(KEYINPUT19), .ZN(n654) );
  XNOR2_X1 U735 ( .A(n654), .B(KEYINPUT78), .ZN(n657) );
  XNOR2_X1 U736 ( .A(G288), .B(G290), .ZN(n655) );
  XNOR2_X1 U737 ( .A(n655), .B(G299), .ZN(n656) );
  XNOR2_X1 U738 ( .A(n657), .B(n656), .ZN(n659) );
  XNOR2_X1 U739 ( .A(G305), .B(n663), .ZN(n658) );
  XNOR2_X1 U740 ( .A(n659), .B(n658), .ZN(n909) );
  XNOR2_X1 U741 ( .A(n909), .B(n660), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n661), .A2(G868), .ZN(n662) );
  XOR2_X1 U743 ( .A(KEYINPUT79), .B(n662), .Z(n665) );
  OR2_X1 U744 ( .A1(n663), .A2(G868), .ZN(n664) );
  NAND2_X1 U745 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U750 ( .A1(n669), .A2(G2072), .ZN(n670) );
  XNOR2_X1 U751 ( .A(KEYINPUT80), .B(n670), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U753 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U754 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U755 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U756 ( .A1(G96), .A2(n673), .ZN(n834) );
  NAND2_X1 U757 ( .A1(n834), .A2(G2106), .ZN(n677) );
  NAND2_X1 U758 ( .A1(G108), .A2(G120), .ZN(n674) );
  NOR2_X1 U759 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U760 ( .A1(G69), .A2(n675), .ZN(n835) );
  NAND2_X1 U761 ( .A1(n835), .A2(G567), .ZN(n676) );
  NAND2_X1 U762 ( .A1(n677), .A2(n676), .ZN(n846) );
  NAND2_X1 U763 ( .A1(G661), .A2(G483), .ZN(n678) );
  NOR2_X1 U764 ( .A1(n846), .A2(n678), .ZN(n679) );
  XOR2_X1 U765 ( .A(KEYINPUT81), .B(n679), .Z(n832) );
  NAND2_X1 U766 ( .A1(n832), .A2(G36), .ZN(G176) );
  XNOR2_X1 U767 ( .A(KEYINPUT85), .B(G166), .ZN(G303) );
  NOR2_X1 U768 ( .A1(G164), .A2(G1384), .ZN(n779) );
  NAND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n778) );
  INV_X1 U770 ( .A(n778), .ZN(n681) );
  NOR2_X1 U771 ( .A1(G1981), .A2(G305), .ZN(n682) );
  XOR2_X1 U772 ( .A(n682), .B(KEYINPUT24), .Z(n683) );
  NOR2_X1 U773 ( .A1(n774), .A2(n683), .ZN(n767) );
  XNOR2_X1 U774 ( .A(G1981), .B(KEYINPUT99), .ZN(n684) );
  XNOR2_X1 U775 ( .A(n684), .B(G305), .ZN(n984) );
  NOR2_X1 U776 ( .A1(G1976), .A2(G288), .ZN(n976) );
  NAND2_X1 U777 ( .A1(n976), .A2(KEYINPUT33), .ZN(n685) );
  NOR2_X1 U778 ( .A1(n774), .A2(n685), .ZN(n686) );
  XOR2_X1 U779 ( .A(KEYINPUT98), .B(n686), .Z(n687) );
  NAND2_X1 U780 ( .A1(n984), .A2(n687), .ZN(n765) );
  NOR2_X1 U781 ( .A1(G2084), .A2(n740), .ZN(n691) );
  AND2_X1 U782 ( .A1(G8), .A2(n691), .ZN(n688) );
  NOR2_X1 U783 ( .A1(G1966), .A2(n774), .ZN(n689) );
  OR2_X1 U784 ( .A1(n688), .A2(n689), .ZN(n732) );
  INV_X1 U785 ( .A(n689), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U787 ( .A(KEYINPUT30), .B(n694), .ZN(n695) );
  XNOR2_X1 U788 ( .A(n696), .B(KEYINPUT93), .ZN(n700) );
  XOR2_X1 U789 ( .A(G2078), .B(KEYINPUT25), .Z(n957) );
  NOR2_X1 U790 ( .A1(n957), .A2(n740), .ZN(n698) );
  NOR2_X1 U791 ( .A1(n719), .A2(G1961), .ZN(n697) );
  NOR2_X1 U792 ( .A1(n698), .A2(n697), .ZN(n731) );
  NAND2_X1 U793 ( .A1(n731), .A2(G301), .ZN(n699) );
  NAND2_X1 U794 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U795 ( .A(KEYINPUT31), .B(n701), .ZN(n746) );
  NAND2_X1 U796 ( .A1(n702), .A2(G1341), .ZN(n703) );
  XNOR2_X1 U797 ( .A(n703), .B(KEYINPUT90), .ZN(n704) );
  NAND2_X1 U798 ( .A1(n704), .A2(n974), .ZN(n708) );
  NAND2_X1 U799 ( .A1(n719), .A2(G1996), .ZN(n706) );
  INV_X1 U800 ( .A(KEYINPUT26), .ZN(n705) );
  XNOR2_X1 U801 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n715) );
  NAND2_X1 U803 ( .A1(n715), .A2(n910), .ZN(n713) );
  NAND2_X1 U804 ( .A1(G1348), .A2(n740), .ZN(n710) );
  NAND2_X1 U805 ( .A1(G2067), .A2(n719), .ZN(n709) );
  NAND2_X1 U806 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U807 ( .A(KEYINPUT91), .B(n711), .Z(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U809 ( .A(n714), .B(KEYINPUT92), .ZN(n717) );
  OR2_X1 U810 ( .A1(n715), .A2(n910), .ZN(n716) );
  NAND2_X1 U811 ( .A1(n717), .A2(n716), .ZN(n724) );
  INV_X1 U812 ( .A(G299), .ZN(n977) );
  NAND2_X1 U813 ( .A1(G1956), .A2(n740), .ZN(n718) );
  XNOR2_X1 U814 ( .A(KEYINPUT89), .B(n718), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n719), .A2(G2072), .ZN(n720) );
  XNOR2_X1 U816 ( .A(KEYINPUT27), .B(n720), .ZN(n721) );
  NOR2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n977), .A2(n725), .ZN(n723) );
  NAND2_X1 U819 ( .A1(n724), .A2(n723), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n977), .A2(n725), .ZN(n726) );
  XOR2_X1 U821 ( .A(n726), .B(KEYINPUT28), .Z(n727) );
  NAND2_X1 U822 ( .A1(n728), .A2(n727), .ZN(n730) );
  OR2_X1 U823 ( .A1(n731), .A2(G301), .ZN(n737) );
  INV_X1 U824 ( .A(n732), .ZN(n733) );
  AND2_X1 U825 ( .A1(n737), .A2(n733), .ZN(n734) );
  NAND2_X1 U826 ( .A1(n738), .A2(n734), .ZN(n735) );
  AND2_X1 U827 ( .A1(n736), .A2(n735), .ZN(n771) );
  NAND2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n987) );
  AND2_X1 U829 ( .A1(n771), .A2(n987), .ZN(n754) );
  NAND2_X1 U830 ( .A1(n738), .A2(n737), .ZN(n748) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n774), .ZN(n739) );
  XNOR2_X1 U832 ( .A(n739), .B(KEYINPUT94), .ZN(n742) );
  NOR2_X1 U833 ( .A1(n740), .A2(G2090), .ZN(n741) );
  NOR2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U835 ( .A1(n743), .A2(G303), .ZN(n744) );
  XOR2_X1 U836 ( .A(KEYINPUT95), .B(n744), .Z(n745) );
  OR2_X1 U837 ( .A1(n690), .A2(n745), .ZN(n749) );
  AND2_X1 U838 ( .A1(n746), .A2(n749), .ZN(n747) );
  NAND2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n752) );
  INV_X1 U840 ( .A(n749), .ZN(n750) );
  OR2_X1 U841 ( .A1(n750), .A2(G286), .ZN(n751) );
  NAND2_X1 U842 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U843 ( .A(n753), .B(KEYINPUT32), .ZN(n770) );
  NAND2_X1 U844 ( .A1(n754), .A2(n770), .ZN(n761) );
  INV_X1 U845 ( .A(n987), .ZN(n758) );
  NOR2_X1 U846 ( .A1(G1971), .A2(G303), .ZN(n755) );
  XNOR2_X1 U847 ( .A(KEYINPUT96), .B(n755), .ZN(n756) );
  NOR2_X1 U848 ( .A1(n976), .A2(n756), .ZN(n757) );
  OR2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n759) );
  OR2_X1 U850 ( .A1(n774), .A2(n759), .ZN(n760) );
  NAND2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U852 ( .A1(KEYINPUT33), .A2(n762), .ZN(n763) );
  XOR2_X1 U853 ( .A(KEYINPUT97), .B(n763), .Z(n764) );
  NOR2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n777) );
  NOR2_X1 U856 ( .A1(G2090), .A2(G303), .ZN(n768) );
  NAND2_X1 U857 ( .A1(G8), .A2(n768), .ZN(n769) );
  XNOR2_X1 U858 ( .A(n769), .B(KEYINPUT100), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n781) );
  NOR2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n823) );
  XNOR2_X1 U864 ( .A(G1986), .B(G290), .ZN(n979) );
  NAND2_X1 U865 ( .A1(n823), .A2(n979), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n810) );
  XNOR2_X1 U867 ( .A(KEYINPUT87), .B(KEYINPUT35), .ZN(n785) );
  NAND2_X1 U868 ( .A1(G116), .A2(n521), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G128), .A2(n888), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n785), .B(n784), .ZN(n791) );
  NAND2_X1 U872 ( .A1(n884), .A2(G140), .ZN(n786) );
  XNOR2_X1 U873 ( .A(n786), .B(KEYINPUT86), .ZN(n788) );
  NAND2_X1 U874 ( .A1(G104), .A2(n883), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U876 ( .A(KEYINPUT34), .B(n789), .ZN(n790) );
  NOR2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U878 ( .A(KEYINPUT36), .B(n792), .ZN(n905) );
  XNOR2_X1 U879 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NOR2_X1 U880 ( .A1(n905), .A2(n820), .ZN(n940) );
  NAND2_X1 U881 ( .A1(n823), .A2(n940), .ZN(n818) );
  NAND2_X1 U882 ( .A1(G119), .A2(n888), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G131), .A2(n884), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U885 ( .A1(G107), .A2(n521), .ZN(n796) );
  NAND2_X1 U886 ( .A1(G95), .A2(n883), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n797) );
  OR2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n900) );
  NAND2_X1 U889 ( .A1(G1991), .A2(n900), .ZN(n808) );
  NAND2_X1 U890 ( .A1(G117), .A2(n521), .ZN(n800) );
  NAND2_X1 U891 ( .A1(G129), .A2(n888), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U893 ( .A1(n883), .A2(G105), .ZN(n801) );
  XOR2_X1 U894 ( .A(KEYINPUT38), .B(n801), .Z(n802) );
  NOR2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U896 ( .A(n804), .B(KEYINPUT88), .ZN(n806) );
  NAND2_X1 U897 ( .A1(G141), .A2(n884), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n899) );
  NAND2_X1 U899 ( .A1(G1996), .A2(n899), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n936) );
  NAND2_X1 U901 ( .A1(n823), .A2(n936), .ZN(n812) );
  NAND2_X1 U902 ( .A1(n818), .A2(n812), .ZN(n809) );
  XNOR2_X1 U903 ( .A(n811), .B(KEYINPUT101), .ZN(n825) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n899), .ZN(n929) );
  INV_X1 U905 ( .A(n812), .ZN(n815) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n900), .ZN(n934) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U908 ( .A1(n934), .A2(n813), .ZN(n814) );
  NOR2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U910 ( .A1(n929), .A2(n816), .ZN(n817) );
  XNOR2_X1 U911 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n905), .A2(n820), .ZN(n943) );
  NAND2_X1 U914 ( .A1(n821), .A2(n943), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U917 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n827), .ZN(G217) );
  INV_X1 U919 ( .A(G661), .ZN(n829) );
  NAND2_X1 U920 ( .A1(G2), .A2(G15), .ZN(n828) );
  NOR2_X1 U921 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U922 ( .A(KEYINPUT104), .B(n830), .Z(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U924 ( .A1(n832), .A2(n831), .ZN(n833) );
  XOR2_X1 U925 ( .A(KEYINPUT105), .B(n833), .Z(G188) );
  XOR2_X1 U926 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  INV_X1 U928 ( .A(G108), .ZN(G238) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  NOR2_X1 U930 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U932 ( .A(G1348), .B(G2454), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n836), .B(G2430), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n837), .B(G1341), .ZN(n843) );
  XOR2_X1 U935 ( .A(G2443), .B(G2427), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2438), .B(G2446), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n841) );
  XOR2_X1 U938 ( .A(G2451), .B(G2435), .Z(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  NAND2_X1 U941 ( .A1(n844), .A2(G14), .ZN(n845) );
  XOR2_X1 U942 ( .A(KEYINPUT102), .B(n845), .Z(n919) );
  XOR2_X1 U943 ( .A(KEYINPUT103), .B(n919), .Z(G401) );
  INV_X1 U944 ( .A(n846), .ZN(G319) );
  XOR2_X1 U945 ( .A(G1976), .B(G1971), .Z(n848) );
  XNOR2_X1 U946 ( .A(G1961), .B(G1956), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U948 ( .A(n849), .B(KEYINPUT41), .Z(n851) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U951 ( .A(G2474), .B(G1981), .Z(n853) );
  XNOR2_X1 U952 ( .A(G1986), .B(G1966), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U955 ( .A(KEYINPUT107), .B(G2090), .Z(n857) );
  XNOR2_X1 U956 ( .A(G2078), .B(G2084), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(n858), .B(G2096), .Z(n860) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U961 ( .A(KEYINPUT43), .B(G2678), .Z(n862) );
  XNOR2_X1 U962 ( .A(KEYINPUT42), .B(G2100), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U964 ( .A(n864), .B(n863), .Z(G227) );
  NAND2_X1 U965 ( .A1(G124), .A2(n888), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n865), .B(KEYINPUT108), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G112), .A2(n521), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G100), .A2(n883), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G136), .A2(n884), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U973 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U974 ( .A1(G118), .A2(n521), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n873), .B(KEYINPUT110), .ZN(n882) );
  NAND2_X1 U976 ( .A1(n888), .A2(G130), .ZN(n874) );
  XNOR2_X1 U977 ( .A(KEYINPUT109), .B(n874), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G106), .A2(n883), .ZN(n876) );
  NAND2_X1 U979 ( .A1(G142), .A2(n884), .ZN(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(n877), .ZN(n878) );
  XNOR2_X1 U982 ( .A(KEYINPUT45), .B(n878), .ZN(n879) );
  NOR2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  NAND2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n898) );
  XOR2_X1 U985 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n896) );
  NAND2_X1 U986 ( .A1(G103), .A2(n883), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G139), .A2(n884), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n894) );
  NAND2_X1 U989 ( .A1(G115), .A2(n521), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G127), .A2(n888), .ZN(n889) );
  NAND2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U992 ( .A(KEYINPUT112), .B(n891), .Z(n892) );
  XNOR2_X1 U993 ( .A(KEYINPUT47), .B(n892), .ZN(n893) );
  NOR2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n923) );
  XNOR2_X1 U995 ( .A(n923), .B(G162), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n933), .B(n899), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(G160), .B(n902), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n905), .B(G164), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n908), .ZN(G395) );
  XOR2_X1 U1005 ( .A(KEYINPUT113), .B(n909), .Z(n912) );
  XNOR2_X1 U1006 ( .A(n910), .B(G286), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n914) );
  XOR2_X1 U1008 ( .A(n974), .B(G171), .Z(n913) );
  XNOR2_X1 U1009 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n915), .ZN(G397) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n916) );
  XOR2_X1 U1012 ( .A(KEYINPUT49), .B(n916), .Z(n917) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n917), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n922) );
  XNOR2_X1 U1020 ( .A(KEYINPUT116), .B(n922), .ZN(n926) );
  XOR2_X1 U1021 ( .A(n923), .B(KEYINPUT115), .Z(n924) );
  XOR2_X1 U1022 ( .A(G2072), .B(n924), .Z(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(KEYINPUT50), .B(n927), .ZN(n932) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT51), .B(n930), .Z(n931) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n945) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n938) );
  XOR2_X1 U1030 ( .A(G160), .B(G2084), .Z(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n941), .B(KEYINPUT114), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n946), .ZN(n947) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n970) );
  NAND2_X1 U1039 ( .A1(n947), .A2(n970), .ZN(n948) );
  NAND2_X1 U1040 ( .A1(n948), .A2(G29), .ZN(n1031) );
  XOR2_X1 U1041 ( .A(G2090), .B(G35), .Z(n963) );
  XOR2_X1 U1042 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n961) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G32), .B(G1996), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n956) );
  XOR2_X1 U1046 ( .A(G1991), .B(G25), .Z(n951) );
  NAND2_X1 U1047 ( .A1(n951), .A2(G28), .ZN(n954) );
  XOR2_X1 U1048 ( .A(KEYINPUT117), .B(G2072), .Z(n952) );
  XNOR2_X1 U1049 ( .A(G33), .B(n952), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(G27), .B(n957), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(n961), .B(n960), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(KEYINPUT119), .B(n964), .ZN(n968) );
  XOR2_X1 U1057 ( .A(G34), .B(KEYINPUT120), .Z(n966) );
  XNOR2_X1 U1058 ( .A(G2084), .B(KEYINPUT54), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(n966), .B(n965), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(n970), .B(n969), .ZN(n972) );
  INV_X1 U1062 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(G11), .A2(n973), .ZN(n1029) );
  XNOR2_X1 U1065 ( .A(G16), .B(KEYINPUT56), .ZN(n999) );
  XOR2_X1 U1066 ( .A(G1341), .B(n974), .Z(n975) );
  NOR2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n997) );
  XNOR2_X1 U1068 ( .A(n977), .B(G1956), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(G1971), .B(G303), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n995) );
  XOR2_X1 U1072 ( .A(G1966), .B(G168), .Z(n982) );
  XNOR2_X1 U1073 ( .A(KEYINPUT121), .B(n982), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(n986), .B(n985), .ZN(n993) );
  XNOR2_X1 U1077 ( .A(G171), .B(G1961), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(G1348), .B(n989), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1084 ( .A1(n999), .A2(n998), .ZN(n1027) );
  INV_X1 U1085 ( .A(G16), .ZN(n1025) );
  XNOR2_X1 U1086 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n1009) );
  XNOR2_X1 U1087 ( .A(KEYINPUT59), .B(G1348), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1000), .B(G4), .ZN(n1007) );
  XNOR2_X1 U1089 ( .A(G1956), .B(G20), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(G1341), .B(G19), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(G6), .B(G1981), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT123), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(n1009), .B(n1008), .ZN(n1021) );
  XOR2_X1 U1097 ( .A(G1986), .B(G24), .Z(n1013) );
  XNOR2_X1 U1098 ( .A(G1971), .B(G22), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(G23), .B(G1976), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(n1015), .B(n1014), .ZN(n1019) );
  XNOR2_X1 U1104 ( .A(G1966), .B(G21), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(G5), .B(G1961), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(n1023), .B(n1022), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1115 ( .A(n1032), .B(KEYINPUT62), .ZN(n1033) );
  XNOR2_X1 U1116 ( .A(KEYINPUT127), .B(n1033), .ZN(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

