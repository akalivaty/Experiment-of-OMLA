

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579;

  NOR2_X1 U322 ( .A1(n515), .A2(n446), .ZN(n560) );
  XOR2_X1 U323 ( .A(G134GAT), .B(G162GAT), .Z(n430) );
  INV_X1 U324 ( .A(KEYINPUT115), .ZN(n415) );
  XNOR2_X1 U325 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U326 ( .A(n384), .B(n383), .ZN(n385) );
  INV_X1 U327 ( .A(G190GAT), .ZN(n447) );
  XNOR2_X1 U328 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U329 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT18), .B(G190GAT), .Z(n291) );
  XNOR2_X1 U331 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U333 ( .A(KEYINPUT17), .B(n292), .Z(n328) );
  XOR2_X1 U334 ( .A(KEYINPUT89), .B(G71GAT), .Z(n294) );
  XNOR2_X1 U335 ( .A(G15GAT), .B(G99GAT), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U337 ( .A(n328), .B(n295), .ZN(n305) );
  XOR2_X1 U338 ( .A(KEYINPUT0), .B(G127GAT), .Z(n431) );
  XOR2_X1 U339 ( .A(n431), .B(G120GAT), .Z(n297) );
  NAND2_X1 U340 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U342 ( .A(n298), .B(G134GAT), .Z(n303) );
  XOR2_X1 U343 ( .A(KEYINPUT20), .B(G176GAT), .Z(n300) );
  XNOR2_X1 U344 ( .A(G169GAT), .B(G113GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(n301), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X2 U348 ( .A(n305), .B(n304), .ZN(n515) );
  XOR2_X1 U349 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n307) );
  XNOR2_X1 U350 ( .A(G106GAT), .B(KEYINPUT90), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U352 ( .A(G148GAT), .B(KEYINPUT91), .Z(n309) );
  XNOR2_X1 U353 ( .A(G141GAT), .B(KEYINPUT24), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U355 ( .A(n311), .B(n310), .Z(n322) );
  XNOR2_X1 U356 ( .A(G78GAT), .B(KEYINPUT78), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n312), .B(G204GAT), .ZN(n408) );
  XOR2_X1 U358 ( .A(n408), .B(G22GAT), .Z(n314) );
  NAND2_X1 U359 ( .A1(G228GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n314), .B(n313), .ZN(n320) );
  XOR2_X1 U361 ( .A(G155GAT), .B(KEYINPUT3), .Z(n316) );
  XNOR2_X1 U362 ( .A(KEYINPUT2), .B(KEYINPUT94), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n439) );
  XOR2_X1 U364 ( .A(G218GAT), .B(KEYINPUT84), .Z(n382) );
  XOR2_X1 U365 ( .A(n439), .B(n382), .Z(n318) );
  XNOR2_X1 U366 ( .A(G50GAT), .B(G162GAT), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U369 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U370 ( .A(KEYINPUT21), .B(KEYINPUT93), .Z(n324) );
  XNOR2_X1 U371 ( .A(KEYINPUT92), .B(G211GAT), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U373 ( .A(G197GAT), .B(n325), .Z(n327) );
  XOR2_X1 U374 ( .A(n326), .B(n327), .Z(n459) );
  XNOR2_X1 U375 ( .A(n328), .B(n327), .ZN(n338) );
  XOR2_X1 U376 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n330) );
  XNOR2_X1 U377 ( .A(G204GAT), .B(G92GAT), .ZN(n329) );
  XNOR2_X1 U378 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U379 ( .A(G176GAT), .B(G64GAT), .Z(n395) );
  XOR2_X1 U380 ( .A(n395), .B(G218GAT), .Z(n332) );
  XOR2_X1 U381 ( .A(G169GAT), .B(G8GAT), .Z(n346) );
  XNOR2_X1 U382 ( .A(G36GAT), .B(n346), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U384 ( .A(n334), .B(n333), .Z(n336) );
  NAND2_X1 U385 ( .A1(G226GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n338), .B(n337), .ZN(n513) );
  XOR2_X1 U388 ( .A(G43GAT), .B(G29GAT), .Z(n340) );
  XNOR2_X1 U389 ( .A(KEYINPUT72), .B(G50GAT), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U391 ( .A(n341), .B(KEYINPUT8), .Z(n343) );
  XNOR2_X1 U392 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n343), .B(n342), .ZN(n388) );
  XOR2_X1 U394 ( .A(KEYINPUT73), .B(KEYINPUT68), .Z(n345) );
  XNOR2_X1 U395 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n350) );
  XOR2_X1 U397 ( .A(KEYINPUT69), .B(G197GAT), .Z(n348) );
  XOR2_X1 U398 ( .A(G22GAT), .B(G15GAT), .Z(n368) );
  XNOR2_X1 U399 ( .A(n346), .B(n368), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U401 ( .A(n350), .B(n349), .Z(n352) );
  NAND2_X1 U402 ( .A1(G229GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U403 ( .A(n352), .B(n351), .ZN(n354) );
  INV_X1 U404 ( .A(KEYINPUT29), .ZN(n353) );
  XNOR2_X1 U405 ( .A(n354), .B(n353), .ZN(n357) );
  XNOR2_X1 U406 ( .A(G141GAT), .B(G113GAT), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n355), .B(G1GAT), .ZN(n427) );
  XNOR2_X1 U408 ( .A(n427), .B(KEYINPUT30), .ZN(n356) );
  XNOR2_X1 U409 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U410 ( .A(n388), .B(n358), .Z(n564) );
  XOR2_X1 U411 ( .A(KEYINPUT74), .B(n564), .Z(n552) );
  XOR2_X1 U412 ( .A(G155GAT), .B(G78GAT), .Z(n360) );
  XNOR2_X1 U413 ( .A(G127GAT), .B(G211GAT), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n374) );
  XOR2_X1 U415 ( .A(G57GAT), .B(G183GAT), .Z(n362) );
  XNOR2_X1 U416 ( .A(G1GAT), .B(G8GAT), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U418 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n364) );
  XNOR2_X1 U419 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U421 ( .A(n366), .B(n365), .ZN(n372) );
  XNOR2_X1 U422 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n367), .B(KEYINPUT75), .ZN(n396) );
  XOR2_X1 U424 ( .A(n396), .B(n368), .Z(n370) );
  NAND2_X1 U425 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n545) );
  INV_X1 U429 ( .A(KEYINPUT36), .ZN(n393) );
  XOR2_X1 U430 ( .A(KEYINPUT85), .B(KEYINPUT10), .Z(n376) );
  XNOR2_X1 U431 ( .A(G190GAT), .B(KEYINPUT66), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U433 ( .A(KEYINPUT65), .B(KEYINPUT11), .Z(n378) );
  XNOR2_X1 U434 ( .A(KEYINPUT64), .B(KEYINPUT9), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U436 ( .A(n380), .B(n379), .Z(n386) );
  XOR2_X1 U437 ( .A(n430), .B(KEYINPUT86), .Z(n384) );
  NAND2_X1 U438 ( .A1(G232GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U439 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U441 ( .A(KEYINPUT79), .B(G92GAT), .Z(n390) );
  XNOR2_X1 U442 ( .A(G99GAT), .B(G85GAT), .ZN(n389) );
  XNOR2_X1 U443 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U444 ( .A(G106GAT), .B(n391), .Z(n400) );
  XNOR2_X1 U445 ( .A(n392), .B(n400), .ZN(n549) );
  XNOR2_X1 U446 ( .A(KEYINPUT87), .B(n549), .ZN(n533) );
  XNOR2_X1 U447 ( .A(n393), .B(n533), .ZN(n577) );
  NOR2_X1 U448 ( .A1(n545), .A2(n577), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n394), .B(KEYINPUT45), .ZN(n413) );
  XOR2_X1 U450 ( .A(n396), .B(n395), .Z(n398) );
  NAND2_X1 U451 ( .A1(G230GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n400), .B(n399), .ZN(n412) );
  XOR2_X1 U454 ( .A(KEYINPUT76), .B(KEYINPUT81), .Z(n402) );
  XNOR2_X1 U455 ( .A(KEYINPUT82), .B(KEYINPUT32), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U457 ( .A(KEYINPUT80), .B(KEYINPUT31), .Z(n404) );
  XNOR2_X1 U458 ( .A(KEYINPUT33), .B(KEYINPUT77), .ZN(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U460 ( .A(n406), .B(n405), .Z(n410) );
  XNOR2_X1 U461 ( .A(G120GAT), .B(G148GAT), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n407), .B(G57GAT), .ZN(n426) );
  XNOR2_X1 U463 ( .A(n408), .B(n426), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U465 ( .A(n412), .B(n411), .ZN(n451) );
  NAND2_X1 U466 ( .A1(n413), .A2(n451), .ZN(n414) );
  NOR2_X1 U467 ( .A1(n552), .A2(n414), .ZN(n416) );
  XNOR2_X1 U468 ( .A(n416), .B(n415), .ZN(n423) );
  INV_X1 U469 ( .A(n545), .ZN(n572) );
  INV_X1 U470 ( .A(n451), .ZN(n569) );
  XNOR2_X1 U471 ( .A(KEYINPUT41), .B(n569), .ZN(n541) );
  NOR2_X1 U472 ( .A1(n564), .A2(n541), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n417), .B(KEYINPUT46), .ZN(n418) );
  NOR2_X1 U474 ( .A1(n572), .A2(n418), .ZN(n419) );
  NAND2_X1 U475 ( .A1(n419), .A2(n549), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n420), .B(KEYINPUT47), .ZN(n421) );
  XNOR2_X1 U477 ( .A(KEYINPUT114), .B(n421), .ZN(n422) );
  NOR2_X1 U478 ( .A1(n423), .A2(n422), .ZN(n424) );
  XNOR2_X1 U479 ( .A(KEYINPUT48), .B(n424), .ZN(n537) );
  NOR2_X1 U480 ( .A1(n513), .A2(n537), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n425), .B(KEYINPUT54), .ZN(n444) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n443) );
  XOR2_X1 U483 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n429) );
  XNOR2_X1 U484 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n435) );
  XOR2_X1 U486 ( .A(G85GAT), .B(n430), .Z(n433) );
  XNOR2_X1 U487 ( .A(G29GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U489 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n438), .B(KEYINPUT6), .Z(n441) );
  XNOR2_X1 U493 ( .A(n439), .B(KEYINPUT4), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n465) );
  XNOR2_X1 U496 ( .A(KEYINPUT97), .B(n465), .ZN(n511) );
  NAND2_X1 U497 ( .A1(n444), .A2(n511), .ZN(n562) );
  NOR2_X1 U498 ( .A1(n459), .A2(n562), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n445), .B(KEYINPUT55), .ZN(n446) );
  NAND2_X1 U500 ( .A1(n560), .A2(n533), .ZN(n450) );
  XOR2_X1 U501 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n448) );
  NAND2_X1 U502 ( .A1(n451), .A2(n552), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n452), .B(KEYINPUT83), .ZN(n483) );
  INV_X1 U504 ( .A(n515), .ZN(n523) );
  XNOR2_X1 U505 ( .A(n513), .B(KEYINPUT27), .ZN(n456) );
  NOR2_X1 U506 ( .A1(n511), .A2(n456), .ZN(n539) );
  XNOR2_X1 U507 ( .A(n459), .B(KEYINPUT28), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n453), .B(KEYINPUT67), .ZN(n518) );
  NAND2_X1 U509 ( .A1(n539), .A2(n518), .ZN(n521) );
  XNOR2_X1 U510 ( .A(KEYINPUT100), .B(n521), .ZN(n454) );
  NOR2_X1 U511 ( .A1(n523), .A2(n454), .ZN(n467) );
  NAND2_X1 U512 ( .A1(n459), .A2(n515), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n455), .B(KEYINPUT26), .ZN(n563) );
  NOR2_X1 U514 ( .A1(n563), .A2(n456), .ZN(n457) );
  XOR2_X1 U515 ( .A(KEYINPUT101), .B(n457), .Z(n462) );
  NOR2_X1 U516 ( .A1(n515), .A2(n513), .ZN(n458) );
  NOR2_X1 U517 ( .A1(n459), .A2(n458), .ZN(n460) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(n460), .Z(n461) );
  NOR2_X1 U519 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n463), .B(KEYINPUT102), .ZN(n464) );
  NOR2_X1 U521 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n479) );
  INV_X1 U523 ( .A(n533), .ZN(n468) );
  NAND2_X1 U524 ( .A1(n468), .A2(n572), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT16), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n470), .B(KEYINPUT88), .ZN(n471) );
  NOR2_X1 U527 ( .A1(n479), .A2(n471), .ZN(n498) );
  NAND2_X1 U528 ( .A1(n483), .A2(n498), .ZN(n477) );
  NOR2_X1 U529 ( .A1(n511), .A2(n477), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT34), .B(n472), .Z(n473) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(n473), .ZN(G1324GAT) );
  NOR2_X1 U532 ( .A1(n513), .A2(n477), .ZN(n474) );
  XOR2_X1 U533 ( .A(G8GAT), .B(n474), .Z(G1325GAT) );
  NOR2_X1 U534 ( .A1(n515), .A2(n477), .ZN(n476) );
  XNOR2_X1 U535 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(G1326GAT) );
  NOR2_X1 U537 ( .A1(n518), .A2(n477), .ZN(n478) );
  XOR2_X1 U538 ( .A(G22GAT), .B(n478), .Z(G1327GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n482) );
  NOR2_X1 U540 ( .A1(n479), .A2(n577), .ZN(n480) );
  NAND2_X1 U541 ( .A1(n480), .A2(n545), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n508) );
  NAND2_X1 U543 ( .A1(n483), .A2(n508), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(KEYINPUT38), .ZN(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT104), .B(n485), .ZN(n495) );
  NOR2_X1 U546 ( .A1(n495), .A2(n511), .ZN(n489) );
  XOR2_X1 U547 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n487) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  NOR2_X1 U551 ( .A1(n513), .A2(n495), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G36GAT), .B(KEYINPUT107), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1329GAT) );
  NOR2_X1 U554 ( .A1(n515), .A2(n495), .ZN(n493) );
  XNOR2_X1 U555 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U557 ( .A(G43GAT), .B(n494), .Z(G1330GAT) );
  NOR2_X1 U558 ( .A1(n518), .A2(n495), .ZN(n496) );
  XOR2_X1 U559 ( .A(G50GAT), .B(n496), .Z(G1331GAT) );
  XNOR2_X1 U560 ( .A(n541), .B(KEYINPUT109), .ZN(n557) );
  NAND2_X1 U561 ( .A1(n557), .A2(n564), .ZN(n497) );
  XOR2_X1 U562 ( .A(KEYINPUT110), .B(n497), .Z(n509) );
  NAND2_X1 U563 ( .A1(n498), .A2(n509), .ZN(n505) );
  NOR2_X1 U564 ( .A1(n511), .A2(n505), .ZN(n499) );
  XOR2_X1 U565 ( .A(G57GAT), .B(n499), .Z(n500) );
  XNOR2_X1 U566 ( .A(KEYINPUT42), .B(n500), .ZN(G1332GAT) );
  NOR2_X1 U567 ( .A1(n513), .A2(n505), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(KEYINPUT111), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n502), .B(n501), .ZN(G1333GAT) );
  NOR2_X1 U570 ( .A1(n515), .A2(n505), .ZN(n503) );
  XOR2_X1 U571 ( .A(KEYINPUT112), .B(n503), .Z(n504) );
  XNOR2_X1 U572 ( .A(G71GAT), .B(n504), .ZN(G1334GAT) );
  NOR2_X1 U573 ( .A1(n518), .A2(n505), .ZN(n507) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  NAND2_X1 U576 ( .A1(n509), .A2(n508), .ZN(n510) );
  XOR2_X1 U577 ( .A(KEYINPUT113), .B(n510), .Z(n517) );
  NOR2_X1 U578 ( .A1(n511), .A2(n517), .ZN(n512) );
  XOR2_X1 U579 ( .A(G85GAT), .B(n512), .Z(G1336GAT) );
  NOR2_X1 U580 ( .A1(n513), .A2(n517), .ZN(n514) );
  XOR2_X1 U581 ( .A(G92GAT), .B(n514), .Z(G1337GAT) );
  NOR2_X1 U582 ( .A1(n515), .A2(n517), .ZN(n516) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n516), .Z(G1338GAT) );
  NOR2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(n519), .Z(n520) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  XOR2_X1 U587 ( .A(G113GAT), .B(KEYINPUT117), .Z(n526) );
  NOR2_X1 U588 ( .A1(n537), .A2(n521), .ZN(n522) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U590 ( .A(KEYINPUT116), .B(n524), .Z(n534) );
  NAND2_X1 U591 ( .A1(n552), .A2(n534), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U594 ( .A1(n534), .A2(n557), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n532) );
  XOR2_X1 U597 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n530) );
  NAND2_X1 U598 ( .A1(n572), .A2(n534), .ZN(n529) );
  XNOR2_X1 U599 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U602 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  NOR2_X1 U604 ( .A1(n563), .A2(n537), .ZN(n538) );
  NAND2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n548) );
  NOR2_X1 U606 ( .A1(n564), .A2(n548), .ZN(n540) );
  XOR2_X1 U607 ( .A(G141GAT), .B(n540), .Z(G1344GAT) );
  NOR2_X1 U608 ( .A1(n541), .A2(n548), .ZN(n543) );
  XNOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(n544), .ZN(G1345GAT) );
  NOR2_X1 U612 ( .A1(n545), .A2(n548), .ZN(n546) );
  XOR2_X1 U613 ( .A(KEYINPUT120), .B(n546), .Z(n547) );
  XNOR2_X1 U614 ( .A(G155GAT), .B(n547), .ZN(G1346GAT) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1347GAT) );
  NAND2_X1 U618 ( .A1(n560), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n555) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U623 ( .A(KEYINPUT56), .B(n556), .Z(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n572), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT59), .Z(n566) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n573) );
  INV_X1 U630 ( .A(n573), .ZN(n576) );
  OR2_X1 U631 ( .A1(n576), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n571) );
  NAND2_X1 U636 ( .A1(n573), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(n578), .Z(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

