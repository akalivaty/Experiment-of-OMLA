//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1205, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  INV_X1    g0006(.A(G58), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n222), .B1(new_n207), .B2(new_n223), .C1(new_n208), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n203), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n206), .B(new_n215), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G226), .B(G232), .Z(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G1), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(G13), .A3(G20), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(KEYINPUT69), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT69), .ZN(new_n249));
  NAND4_X1  g0049(.A1(new_n249), .A2(new_n246), .A3(G13), .A4(G20), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n212), .B1(new_n203), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n213), .A2(G1), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(G50), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n213), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G150), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n213), .A2(new_n252), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n260), .A2(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G50), .A2(G58), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n213), .B1(new_n265), .B2(new_n208), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n253), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n259), .B(new_n267), .C1(G50), .C2(new_n251), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT68), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G222), .ZN(new_n277));
  INV_X1    g0077(.A(G223), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n275), .B(new_n277), .C1(new_n278), .C2(new_n276), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(G77), .B2(new_n275), .ZN(new_n280));
  INV_X1    g0080(.A(G226), .ZN(new_n281));
  INV_X1    g0081(.A(new_n271), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n246), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n274), .A2(new_n280), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(G274), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT66), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT66), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G45), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n246), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT67), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT67), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n292), .A2(new_n295), .A3(new_n246), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n286), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n285), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n269), .A2(new_n270), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(G200), .B2(new_n299), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n301), .B2(KEYINPUT74), .ZN(new_n304));
  XOR2_X1   g0104(.A(new_n302), .B(new_n304), .Z(new_n305));
  OR2_X1    g0105(.A1(new_n263), .A2(KEYINPUT71), .ZN(new_n306));
  INV_X1    g0106(.A(new_n260), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n263), .A2(KEYINPUT71), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT15), .B(G87), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n309), .B1(new_n213), .B2(new_n217), .C1(new_n261), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n253), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n256), .A2(G77), .A3(new_n258), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(G77), .C2(new_n251), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n275), .A2(G107), .ZN(new_n315));
  MUX2_X1   g0115(.A(new_n223), .B(new_n224), .S(G1698), .Z(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n275), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n282), .A2(new_n283), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n317), .A2(new_n273), .B1(new_n318), .B2(G244), .ZN(new_n319));
  INV_X1    g0119(.A(new_n286), .ZN(new_n320));
  INV_X1    g0120(.A(new_n296), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n295), .B1(new_n292), .B2(new_n246), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n314), .A2(new_n326), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n327), .A2(KEYINPUT73), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(KEYINPUT73), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n324), .A2(G179), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT72), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n299), .A2(new_n325), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n298), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n268), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n319), .A2(G190), .A3(new_n323), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n337), .A2(KEYINPUT70), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n319), .B2(new_n323), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n338), .A2(new_n314), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(KEYINPUT70), .B2(new_n337), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n332), .A2(new_n336), .A3(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n305), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G97), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n223), .A2(G1698), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(G226), .B2(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT3), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G33), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n345), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n273), .A2(new_n352), .B1(new_n318), .B2(G238), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n323), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT13), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n354), .A2(KEYINPUT13), .ZN(new_n357));
  OAI21_X1  g0157(.A(G169), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n353), .A2(new_n323), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT13), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n355), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n358), .A2(KEYINPUT14), .B1(new_n334), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n325), .B1(new_n361), .B2(new_n355), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT14), .ZN(new_n365));
  OR3_X1    g0165(.A1(new_n364), .A2(KEYINPUT76), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT76), .B1(new_n364), .B2(new_n365), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n256), .A2(G68), .A3(new_n258), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT75), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n251), .A2(G68), .ZN(new_n371));
  INV_X1    g0171(.A(G50), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n263), .A2(new_n372), .B1(new_n213), .B2(G68), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n261), .A2(new_n217), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n253), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT11), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n371), .A2(KEYINPUT12), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n371), .A2(KEYINPUT12), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n377), .B(new_n378), .C1(new_n376), .C2(new_n375), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n370), .A2(new_n379), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n368), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n362), .A2(G200), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n382), .B(new_n380), .C1(new_n300), .C2(new_n362), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n209), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G20), .ZN(new_n387));
  INV_X1    g0187(.A(new_n263), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G159), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(KEYINPUT77), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT77), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n213), .B1(new_n209), .B2(new_n385), .ZN(new_n392));
  INV_X1    g0192(.A(G159), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n263), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n391), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n275), .B2(G20), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n351), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n208), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n254), .B1(new_n401), .B2(KEYINPUT16), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n349), .A2(KEYINPUT78), .A3(G33), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n348), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT78), .B1(new_n349), .B2(G33), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT7), .B(new_n213), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n208), .B1(new_n407), .B2(new_n398), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n403), .B1(new_n408), .B2(new_n396), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n402), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n260), .A2(new_n257), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n248), .A2(new_n250), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n256), .A2(new_n411), .B1(new_n412), .B2(new_n260), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n278), .A2(G1698), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT80), .B1(new_n275), .B2(new_n415), .ZN(new_n416));
  AND4_X1   g0216(.A1(KEYINPUT80), .A2(new_n415), .A3(new_n348), .A4(new_n350), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(G226), .A2(G1698), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n348), .A2(new_n350), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT79), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n348), .A2(new_n350), .A3(new_n419), .A4(KEYINPUT79), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G87), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n273), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n284), .A2(new_n223), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n428), .A3(new_n323), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G169), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n297), .A2(new_n427), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(G179), .A3(new_n426), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n414), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT18), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n414), .A2(new_n436), .A3(new_n433), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n426), .A2(new_n300), .A3(new_n428), .A4(new_n323), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT81), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT81), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n431), .A2(new_n441), .A3(new_n300), .A4(new_n426), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n429), .A2(new_n339), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n413), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n402), .B2(new_n409), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT82), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n444), .A2(KEYINPUT82), .A3(new_n446), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(KEYINPUT17), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n444), .A2(new_n446), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT83), .B(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n438), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n344), .A2(new_n384), .A3(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n351), .A2(new_n220), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n276), .ZN(new_n458));
  INV_X1    g0258(.A(G257), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(new_n276), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n275), .A2(new_n460), .B1(G33), .B2(G294), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n273), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n246), .B(G45), .C1(new_n291), .C2(KEYINPUT5), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n464), .A2(KEYINPUT84), .B1(KEYINPUT5), .B2(new_n291), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n287), .A2(G1), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT84), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n466), .B(new_n467), .C1(KEYINPUT5), .C2(new_n291), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n271), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G264), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n320), .A2(new_n468), .A3(new_n465), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n463), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G169), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(KEYINPUT91), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n470), .A2(KEYINPUT91), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n471), .B(new_n463), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n473), .B1(new_n477), .B2(new_n334), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n213), .A2(KEYINPUT23), .A3(G107), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT90), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n479), .A2(new_n480), .B1(KEYINPUT23), .B2(G107), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G116), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT23), .ZN(new_n484));
  AOI21_X1  g0284(.A(G20), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n275), .A2(new_n213), .A3(G87), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n487), .A2(KEYINPUT22), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(KEYINPUT22), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n481), .B(new_n486), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n490), .A2(KEYINPUT24), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(KEYINPUT24), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n253), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n251), .A2(KEYINPUT25), .A3(G107), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT25), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n495), .B1(new_n412), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n251), .B(new_n254), .C1(G1), .C2(new_n252), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AOI211_X1 g0299(.A(new_n494), .B(new_n497), .C1(new_n499), .C2(G107), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n478), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  OR2_X1    g0303(.A1(new_n472), .A2(G190), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n477), .A2(new_n339), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  INV_X1    g0308(.A(G97), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n508), .B(new_n213), .C1(G33), .C2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n510), .B(new_n253), .C1(new_n213), .C2(G116), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT20), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G116), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n412), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n513), .B(new_n515), .C1(new_n498), .C2(new_n514), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G264), .A2(G1698), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n275), .B(new_n517), .C1(new_n459), .C2(G1698), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n273), .B(new_n518), .C1(G303), .C2(new_n275), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n469), .A2(G270), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n471), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n516), .A2(G169), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT21), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n521), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(G179), .A3(new_n516), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n516), .A2(KEYINPUT21), .A3(new_n521), .A4(G169), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n516), .B1(new_n521), .B2(G200), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n300), .B2(new_n521), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n351), .B2(new_n218), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n275), .A2(KEYINPUT4), .A3(G244), .A4(new_n276), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n534), .A2(new_n508), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(G1698), .B1(new_n457), .B2(new_n533), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n274), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n469), .A2(G257), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n471), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n325), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n407), .A2(new_n398), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n496), .A2(KEYINPUT6), .A3(G97), .ZN(new_n546));
  XOR2_X1   g0346(.A(G97), .B(G107), .Z(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(KEYINPUT6), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(G20), .B1(G77), .B2(new_n388), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n254), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n412), .A2(new_n509), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n498), .B2(new_n509), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n541), .A2(new_n334), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n543), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(G200), .B1(new_n538), .B2(new_n540), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n553), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(G190), .B2(new_n541), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g0361(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n562), .B(KEYINPUT87), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n213), .B1(new_n345), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n275), .A2(new_n213), .A3(G68), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n564), .B1(new_n261), .B2(new_n509), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT88), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n566), .A2(KEYINPUT88), .A3(new_n567), .A4(new_n568), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n253), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n310), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n499), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n412), .A2(new_n310), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n275), .A2(G238), .A3(new_n276), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT86), .ZN(new_n579));
  XNOR2_X1  g0379(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n275), .A2(G244), .A3(G1698), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n581), .A2(new_n483), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n274), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n466), .A2(new_n220), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n282), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT85), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n282), .A2(KEYINPUT85), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n320), .A2(new_n466), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n334), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n325), .B1(new_n583), .B2(new_n591), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n577), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n499), .A2(G87), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n596), .B(KEYINPUT89), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n573), .A3(new_n576), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n592), .A2(G190), .ZN(new_n599));
  OAI21_X1  g0399(.A(G200), .B1(new_n583), .B2(new_n591), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n595), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n507), .A2(new_n532), .A3(new_n561), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n456), .A2(new_n604), .ZN(G372));
  INV_X1    g0405(.A(new_n456), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT94), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n595), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n577), .A2(new_n593), .A3(KEYINPUT94), .A4(new_n594), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n573), .A2(new_n576), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n611), .A2(new_n597), .A3(new_n600), .A4(new_n599), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n557), .A2(new_n595), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n610), .B1(new_n613), .B2(KEYINPUT26), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT93), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n524), .B2(new_n528), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n522), .A2(new_n523), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(KEYINPUT93), .A3(new_n526), .A4(new_n527), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n502), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n505), .A2(new_n504), .ZN(new_n620));
  INV_X1    g0420(.A(new_n501), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n560), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n557), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n612), .A2(new_n595), .A3(KEYINPUT92), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT92), .B1(new_n612), .B2(new_n595), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n614), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n606), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g0429(.A(new_n629), .B(KEYINPUT95), .Z(new_n630));
  INV_X1    g0430(.A(new_n336), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n435), .A2(new_n437), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n383), .A2(new_n328), .A3(new_n329), .A4(new_n331), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n381), .A2(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n444), .A2(KEYINPUT82), .A3(new_n446), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT82), .B1(new_n444), .B2(new_n446), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT17), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n452), .A2(new_n453), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n632), .B1(new_n634), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT96), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n305), .B(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n631), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n630), .A2(new_n644), .ZN(G369));
  NAND2_X1  g0445(.A1(new_n616), .A2(new_n618), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n246), .A2(new_n213), .A3(G13), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n516), .A2(new_n652), .ZN(new_n653));
  MUX2_X1   g0453(.A(new_n646), .B(new_n532), .S(new_n653), .Z(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G330), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n501), .A2(new_n652), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT97), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n656), .B(new_n657), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n658), .A2(new_n507), .B1(new_n503), .B2(new_n652), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n529), .A2(new_n652), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(new_n507), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n502), .B2(new_n652), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n660), .A2(new_n663), .ZN(G399));
  OR2_X1    g0464(.A1(new_n563), .A2(G116), .ZN(new_n665));
  INV_X1    g0465(.A(new_n204), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G41), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G1), .ZN(new_n669));
  OAI22_X1  g0469(.A1(new_n665), .A2(new_n669), .B1(new_n210), .B2(new_n668), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  INV_X1    g0471(.A(new_n652), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n628), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT29), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n602), .A2(new_n556), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n610), .B1(new_n676), .B2(new_n624), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n529), .A2(new_n502), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n625), .B2(new_n626), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n622), .A2(new_n556), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT92), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n602), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n612), .A2(new_n595), .A3(KEYINPUT92), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n624), .B1(new_n685), .B2(new_n557), .ZN(new_n686));
  OAI211_X1 g0486(.A(KEYINPUT29), .B(new_n672), .C1(new_n681), .C2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n675), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n592), .A2(new_n525), .A3(G179), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT98), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n477), .A2(new_n542), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n477), .B2(new_n542), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT99), .ZN(new_n694));
  INV_X1    g0494(.A(new_n476), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n695), .A2(new_n474), .B1(new_n273), .B2(new_n462), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n521), .A2(new_n334), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n697), .A3(new_n592), .A4(new_n541), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT30), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT31), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT99), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n701), .B(new_n689), .C1(new_n691), .C2(new_n692), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n694), .A2(new_n699), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(KEYINPUT31), .A2(new_n604), .B1(new_n703), .B2(new_n652), .ZN(new_n704));
  AOI211_X1 g0504(.A(new_n700), .B(new_n672), .C1(new_n699), .C2(new_n693), .ZN(new_n705));
  OAI21_X1  g0505(.A(G330), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n688), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n671), .B1(new_n707), .B2(G1), .ZN(G364));
  AOI21_X1  g0508(.A(new_n212), .B1(G20), .B2(new_n325), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n213), .A2(new_n334), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G200), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n300), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n351), .B1(new_n712), .B2(G50), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n710), .B(KEYINPUT101), .Z(new_n714));
  NOR3_X1   g0514(.A1(new_n714), .A2(new_n300), .A3(G200), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n714), .A2(G190), .A3(G200), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI221_X1 g0518(.A(new_n713), .B1(new_n716), .B2(new_n207), .C1(new_n217), .C2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n339), .A2(G179), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT102), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n300), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G87), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G179), .A2(G200), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(G20), .A3(new_n300), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G159), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n711), .A2(G190), .ZN(new_n729));
  AOI22_X1  g0529(.A1(KEYINPUT32), .A2(new_n728), .B1(new_n729), .B2(G68), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n724), .B(new_n730), .C1(KEYINPUT32), .C2(new_n728), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n213), .B1(new_n725), .B2(G190), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n732), .A2(KEYINPUT103), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(KEYINPUT103), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n509), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n722), .A2(G190), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n739), .B2(new_n496), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n719), .A2(new_n731), .A3(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(G283), .A2(new_n738), .B1(new_n723), .B2(G303), .ZN(new_n742));
  INV_X1    g0542(.A(G294), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(new_n743), .B2(new_n735), .ZN(new_n744));
  INV_X1    g0544(.A(G311), .ZN(new_n745));
  INV_X1    g0545(.A(G322), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n718), .B1(new_n716), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(KEYINPUT33), .A2(G317), .ZN(new_n748));
  AND2_X1   g0548(.A1(KEYINPUT33), .A2(G317), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n729), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n275), .B1(new_n727), .B2(G329), .ZN(new_n751));
  INV_X1    g0551(.A(G326), .ZN(new_n752));
  INV_X1    g0552(.A(new_n712), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n750), .B(new_n751), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n744), .A2(new_n747), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n709), .B1(new_n741), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G13), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n246), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n667), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n275), .A2(new_n204), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT100), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n764), .A2(G355), .B1(new_n514), .B2(new_n666), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n244), .A2(new_n287), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n666), .A2(new_n275), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n288), .A2(new_n290), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n767), .B1(new_n769), .B2(new_n210), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n765), .B1(new_n766), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G13), .A2(G33), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n709), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n762), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n774), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n756), .B(new_n776), .C1(new_n654), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n655), .A2(new_n762), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n654), .A2(G330), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(G396));
  NAND2_X1  g0581(.A1(new_n314), .A2(new_n652), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n332), .A2(new_n342), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n332), .B2(new_n782), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n673), .B(new_n784), .Z(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n706), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n761), .B1(new_n785), .B2(new_n706), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n784), .A2(new_n773), .ZN(new_n789));
  INV_X1    g0589(.A(new_n709), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n729), .A2(G150), .B1(new_n712), .B2(G137), .ZN(new_n791));
  INV_X1    g0591(.A(G143), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n791), .B1(new_n716), .B2(new_n792), .C1(new_n393), .C2(new_n718), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT34), .ZN(new_n794));
  INV_X1    g0594(.A(G132), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n275), .B1(new_n795), .B2(new_n726), .C1(new_n735), .C2(new_n207), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n739), .A2(new_n208), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(G50), .C2(new_n723), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n351), .B1(new_n726), .B2(new_n745), .C1(new_n753), .C2(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n514), .A2(new_n718), .B1(new_n716), .B2(new_n743), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n801), .B(new_n802), .C1(G283), .C2(new_n729), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n723), .A2(G107), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n738), .A2(G87), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n803), .A2(new_n737), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n790), .B1(new_n799), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n709), .A2(new_n772), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n762), .B(new_n807), .C1(new_n217), .C2(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G384));
  NOR2_X1   g0611(.A1(new_n758), .A2(new_n246), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT38), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT37), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n430), .A2(new_n432), .A3(new_n650), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n414), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n449), .A2(new_n814), .A3(new_n450), .A4(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n447), .A2(new_n816), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n455), .A2(new_n446), .A3(new_n650), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT106), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR4_X1   g0622(.A1(new_n455), .A2(KEYINPUT106), .A3(new_n446), .A4(new_n650), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n813), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT104), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n401), .A2(KEYINPUT16), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n403), .B1(new_n396), .B2(new_n400), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n826), .A2(new_n827), .A3(new_n253), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n413), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n815), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n635), .A2(new_n636), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n825), .B1(new_n831), .B2(new_n814), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n449), .A2(new_n450), .ZN(new_n833));
  OAI211_X1 g0633(.A(KEYINPUT104), .B(KEYINPUT37), .C1(new_n833), .C2(new_n830), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n832), .A2(new_n834), .A3(new_n817), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n632), .B1(new_n638), .B2(new_n639), .ZN(new_n836));
  INV_X1    g0636(.A(new_n650), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(new_n837), .A3(new_n829), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n835), .A2(new_n838), .A3(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT108), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT108), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n835), .A2(new_n838), .A3(new_n841), .A4(KEYINPUT38), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n824), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n652), .B1(new_n370), .B2(new_n379), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n383), .B(new_n844), .C1(new_n368), .C2(new_n380), .ZN(new_n845));
  INV_X1    g0645(.A(new_n844), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n366), .A2(new_n367), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(new_n363), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n784), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n604), .A2(KEYINPUT31), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n703), .A2(new_n652), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n694), .A2(new_n699), .A3(new_n702), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n850), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n843), .A2(KEYINPUT40), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT38), .B1(new_n835), .B2(new_n838), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT105), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n839), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI211_X1 g0661(.A(KEYINPUT105), .B(KEYINPUT38), .C1(new_n835), .C2(new_n838), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n856), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  XOR2_X1   g0663(.A(KEYINPUT109), .B(KEYINPUT40), .Z(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT110), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT110), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n863), .A2(new_n867), .A3(new_n864), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n858), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n853), .A2(new_n855), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(new_n606), .A3(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n869), .B1(new_n606), .B2(new_n870), .ZN(new_n873));
  INV_X1    g0673(.A(G330), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT111), .Z(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT39), .B1(new_n861), .B2(new_n862), .ZN(new_n878));
  XNOR2_X1  g0678(.A(KEYINPUT107), .B(KEYINPUT39), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n824), .A2(new_n840), .A3(new_n842), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n381), .A2(new_n652), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n861), .A2(new_n862), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n628), .A2(new_n672), .A3(new_n784), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n332), .A2(new_n652), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n849), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n884), .A2(new_n890), .B1(new_n438), .B2(new_n650), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n606), .A2(new_n675), .A3(new_n687), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n644), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n892), .B(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n812), .B1(new_n877), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n877), .B2(new_n895), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n548), .A2(KEYINPUT35), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n548), .A2(KEYINPUT35), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n898), .A2(G116), .A3(new_n214), .A4(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT36), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n211), .A2(G77), .A3(new_n385), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(G50), .B2(new_n208), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(G1), .A3(new_n757), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n897), .A2(new_n901), .A3(new_n904), .ZN(G367));
  INV_X1    g0705(.A(new_n767), .ZN(new_n906));
  OAI221_X1 g0706(.A(new_n775), .B1(new_n204), .B2(new_n310), .C1(new_n236), .C2(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n907), .A2(new_n761), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n598), .A2(new_n652), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n608), .B2(new_n609), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n685), .B2(new_n909), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(G137), .ZN(new_n913));
  INV_X1    g0713(.A(new_n729), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n275), .B1(new_n726), .B2(new_n913), .C1(new_n914), .C2(new_n393), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n372), .A2(new_n718), .B1(new_n716), .B2(new_n262), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n915), .B(new_n916), .C1(G143), .C2(new_n712), .ZN(new_n917));
  INV_X1    g0717(.A(new_n735), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(G68), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n723), .A2(G58), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n738), .A2(G77), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n917), .A2(new_n919), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(G317), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n351), .B1(new_n726), .B2(new_n923), .C1(new_n753), .C2(new_n745), .ZN(new_n924));
  INV_X1    g0724(.A(G283), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n925), .A2(new_n718), .B1(new_n716), .B2(new_n800), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n924), .B(new_n926), .C1(G294), .C2(new_n729), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n927), .B1(new_n509), .B2(new_n739), .C1(new_n496), .C2(new_n735), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n723), .A2(G116), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT46), .Z(new_n930));
  OAI21_X1  g0730(.A(new_n922), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT47), .Z(new_n932));
  OAI221_X1 g0732(.A(new_n908), .B1(new_n777), .B2(new_n912), .C1(new_n932), .C2(new_n790), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n561), .B1(new_n553), .B2(new_n672), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n557), .A2(new_n652), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(new_n662), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT113), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n556), .B1(new_n934), .B2(new_n502), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT112), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n652), .B1(new_n940), .B2(new_n941), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n938), .A2(KEYINPUT42), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT43), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n911), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n660), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(new_n936), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n939), .A2(new_n944), .A3(new_n946), .A4(new_n911), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT114), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n949), .A2(new_n952), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n955), .B(new_n956), .C1(new_n951), .C2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n663), .A2(new_n936), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT45), .Z(new_n960));
  NAND2_X1  g0760(.A1(new_n663), .A2(new_n936), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT44), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(new_n660), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n659), .B1(new_n529), .B2(new_n652), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n662), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(new_n655), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n707), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n667), .B(KEYINPUT41), .Z(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n760), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n933), .B1(new_n958), .B2(new_n971), .ZN(G387));
  OR2_X1    g0772(.A1(new_n233), .A2(new_n768), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n973), .A2(new_n767), .B1(new_n665), .B2(new_n764), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n307), .A2(new_n372), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT50), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n287), .B1(new_n208), .B2(new_n217), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n976), .A2(new_n665), .A3(new_n977), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n974), .A2(new_n978), .B1(G107), .B2(new_n204), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n762), .B1(new_n979), .B2(new_n775), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n372), .A2(new_n716), .B1(new_n718), .B2(new_n208), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n723), .A2(G77), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n918), .A2(new_n574), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(new_n739), .C2(new_n509), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n753), .A2(new_n393), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n275), .B1(new_n726), .B2(new_n262), .C1(new_n914), .C2(new_n260), .ZN(new_n986));
  NOR4_X1   g0786(.A1(new_n981), .A2(new_n984), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n729), .A2(G311), .B1(new_n712), .B2(G322), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n716), .B2(new_n923), .C1(new_n800), .C2(new_n718), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT48), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n723), .A2(G294), .B1(new_n918), .B2(G283), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT49), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n351), .B1(new_n752), .B2(new_n726), .C1(new_n739), .C2(new_n514), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n995), .B2(KEYINPUT49), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n987), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n980), .B1(new_n999), .B2(new_n790), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n659), .B2(new_n774), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n967), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1001), .B1(new_n1002), .B2(new_n760), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n707), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n667), .B(KEYINPUT115), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1002), .A2(new_n707), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1003), .B1(new_n1006), .B2(new_n1007), .ZN(G393));
  XNOR2_X1  g0808(.A(new_n963), .B(new_n950), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n760), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n241), .A2(new_n906), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n775), .B1(new_n509), .B2(new_n204), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n761), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n715), .A2(G311), .B1(G317), .B2(new_n712), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT52), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n351), .B1(new_n726), .B2(new_n746), .C1(new_n914), .C2(new_n800), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n717), .B2(G294), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n723), .A2(G283), .B1(new_n918), .B2(G116), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n496), .C2(new_n739), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n715), .A2(G159), .B1(G150), .B2(new_n712), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT51), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n275), .B1(new_n726), .B2(new_n792), .C1(new_n914), .C2(new_n372), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n717), .B2(new_n307), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n918), .A2(G77), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n723), .A2(G68), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1023), .A2(new_n805), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1015), .A2(new_n1019), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1013), .B1(new_n1027), .B2(new_n709), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n936), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n777), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1010), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1004), .ZN(new_n1032));
  OAI21_X1  g0832(.A(KEYINPUT116), .B1(new_n1009), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT116), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n964), .A2(new_n1034), .A3(new_n1004), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1005), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n1009), .B2(new_n1032), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1031), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(G390));
  INV_X1    g0840(.A(new_n882), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n888), .B2(new_n889), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n878), .A2(new_n880), .A3(new_n1042), .ZN(new_n1043));
  OAI211_X1 g0843(.A(G330), .B(new_n784), .C1(new_n704), .C2(new_n705), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1044), .A2(new_n889), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n672), .B(new_n784), .C1(new_n681), .C2(new_n686), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n887), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n882), .B1(new_n1047), .B2(new_n849), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1045), .B1(new_n843), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT117), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n1043), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1050), .B1(new_n1043), .B2(new_n1049), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n843), .A2(new_n1048), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1043), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n874), .B1(new_n853), .B2(new_n855), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n850), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1053), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n760), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n808), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n761), .B1(new_n1062), .B2(new_n307), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n351), .B1(new_n726), .B2(new_n743), .C1(new_n753), .C2(new_n925), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n509), .A2(new_n718), .B1(new_n716), .B2(new_n514), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(G107), .C2(new_n729), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n797), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1066), .A2(new_n724), .A3(new_n1067), .A4(new_n1024), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n723), .A2(G150), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT53), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(KEYINPUT54), .B(G143), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n718), .A2(new_n1071), .B1(new_n913), .B2(new_n914), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT118), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n351), .B1(new_n727), .B2(G125), .ZN(new_n1074));
  INV_X1    g0874(.A(G128), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n753), .C1(new_n716), .C2(new_n795), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G159), .B2(new_n918), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1073), .B(new_n1077), .C1(new_n372), .C2(new_n739), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1068), .B1(new_n1070), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1063), .B1(new_n1079), .B2(new_n709), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n881), .B2(new_n773), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1061), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1056), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n893), .B(new_n644), .C1(new_n456), .C2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n849), .B1(new_n1056), .B2(new_n784), .ZN(new_n1085));
  OR3_X1    g0885(.A1(new_n1085), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n888), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1044), .A2(new_n889), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1087), .B1(new_n1059), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1084), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1060), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1091), .A2(new_n1037), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1093), .B(new_n1090), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1082), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(G378));
  AOI22_X1  g0896(.A1(new_n729), .A2(G132), .B1(new_n712), .B2(G125), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n716), .B2(new_n1075), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n723), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1099), .A2(new_n1071), .B1(new_n262), .B2(new_n735), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(G137), .C2(new_n717), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1102), .A2(KEYINPUT59), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(KEYINPUT59), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n738), .A2(G159), .ZN(new_n1105));
  AOI211_X1 g0905(.A(G33), .B(G41), .C1(new_n727), .C2(G124), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n496), .A2(new_n716), .B1(new_n718), .B2(new_n310), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n738), .A2(G58), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n982), .A2(new_n1109), .A3(new_n919), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n275), .A2(G41), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G283), .B2(new_n727), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n509), .B2(new_n914), .C1(new_n514), .C2(new_n753), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1108), .A2(new_n1110), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT58), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1112), .B(new_n372), .C1(G33), .C2(G41), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1115), .A2(KEYINPUT58), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1107), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n709), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n762), .B1(new_n372), .B2(new_n808), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n643), .A2(new_n336), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1123), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n643), .A2(new_n336), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n268), .A2(new_n837), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1124), .A2(new_n268), .A3(new_n837), .A4(new_n1126), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1120), .B(new_n1121), .C1(new_n1131), .C2(new_n773), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n863), .A2(new_n867), .A3(new_n864), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n867), .B1(new_n863), .B2(new_n864), .ZN(new_n1135));
  OAI211_X1 g0935(.A(G330), .B(new_n857), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1131), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n866), .A2(new_n868), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1139), .A2(G330), .A3(new_n857), .A4(new_n1131), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT119), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n883), .B2(new_n891), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1138), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1133), .B1(new_n1145), .B2(new_n760), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1084), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1094), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT120), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1094), .A2(KEYINPUT120), .A3(new_n1147), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT57), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1131), .B1(new_n869), .B2(G330), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n892), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1138), .A2(new_n1140), .A3(new_n883), .A4(new_n891), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1153), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1037), .B1(new_n1152), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT57), .B1(new_n1152), .B2(new_n1145), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT121), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI211_X1 g0962(.A(KEYINPUT121), .B(KEYINPUT57), .C1(new_n1152), .C2(new_n1145), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1146), .B1(new_n1162), .B2(new_n1163), .ZN(G375));
  NAND2_X1  g0964(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n760), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1166), .A2(KEYINPUT122), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1166), .A2(KEYINPUT122), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n889), .A2(new_n772), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n761), .B1(new_n1062), .B2(G68), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n351), .B1(new_n726), .B2(new_n800), .C1(new_n753), .C2(new_n743), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n496), .A2(new_n718), .B1(new_n716), .B2(new_n925), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(G116), .C2(new_n729), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n723), .A2(G97), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1173), .A2(new_n921), .A3(new_n983), .A4(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n723), .A2(G159), .B1(G128), .B2(new_n727), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT123), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n914), .A2(new_n1071), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n351), .B(new_n1178), .C1(G132), .C2(new_n712), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G137), .A2(new_n715), .B1(new_n717), .B2(G150), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n918), .A2(G50), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1109), .A4(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1175), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1170), .B1(new_n1183), .B2(new_n709), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1167), .B(new_n1168), .C1(new_n1169), .C2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1165), .A2(new_n1147), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1090), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n970), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1185), .B1(new_n1186), .B2(new_n1188), .ZN(G381));
  OAI211_X1 g0989(.A(new_n1039), .B(new_n933), .C1(new_n971), .C2(new_n958), .ZN(new_n1190));
  OR2_X1    g0990(.A1(G393), .A2(G396), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1190), .A2(G381), .A3(G384), .A4(new_n1191), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1094), .A2(KEYINPUT120), .A3(new_n1147), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT120), .B1(new_n1094), .B2(new_n1147), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1144), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1138), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1153), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT121), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1200), .A2(new_n1201), .A3(new_n1159), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1192), .A2(new_n1202), .A3(new_n1095), .A4(new_n1146), .ZN(G407));
  NOR2_X1   g1003(.A1(new_n1192), .A2(new_n651), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1095), .A3(new_n1146), .ZN(new_n1205));
  OAI21_X1  g1005(.A(G213), .B1(new_n1204), .B2(new_n1205), .ZN(G409));
  AND2_X1   g1006(.A1(new_n651), .A2(G213), .ZN(new_n1207));
  OAI211_X1 g1007(.A(G378), .B(new_n1146), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1195), .A2(new_n1198), .A3(new_n969), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1132), .B1(new_n1210), .B2(new_n759), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1095), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1207), .B1(new_n1208), .B2(new_n1212), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1037), .B(new_n1090), .C1(new_n1186), .C2(KEYINPUT60), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(KEYINPUT60), .B2(new_n1186), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1185), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n810), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1185), .A2(G384), .A3(new_n1215), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1213), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT63), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1207), .A2(G2897), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1219), .B(new_n1225), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1213), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1213), .A2(KEYINPUT63), .A3(new_n1220), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G387), .A2(G390), .ZN(new_n1229));
  XOR2_X1   g1029(.A(G393), .B(G396), .Z(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1190), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1231), .B1(new_n1229), .B2(new_n1190), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1233), .A2(new_n1234), .A3(KEYINPUT61), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1223), .A2(new_n1227), .A3(new_n1228), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT62), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1213), .A2(new_n1237), .A3(new_n1220), .ZN(new_n1238));
  XOR2_X1   g1038(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1213), .B2(new_n1226), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1237), .B1(new_n1213), .B2(new_n1220), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT125), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1234), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(KEYINPUT125), .A3(new_n1232), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1236), .B1(new_n1242), .B2(new_n1247), .ZN(G405));
  NAND2_X1  g1048(.A1(G375), .A2(new_n1095), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1249), .A2(new_n1208), .A3(new_n1219), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1219), .B1(new_n1249), .B2(new_n1208), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1247), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT127), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1247), .B(KEYINPUT127), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1208), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G378), .B1(new_n1202), .B2(new_n1146), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1220), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1249), .A2(new_n1208), .A3(new_n1219), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT126), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1258), .A2(new_n1259), .A3(KEYINPUT126), .A4(new_n1260), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1254), .A2(new_n1255), .B1(new_n1263), .B2(new_n1264), .ZN(G402));
endmodule


