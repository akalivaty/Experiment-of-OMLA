

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747;

  AND2_X1 U364 ( .A1(n367), .A2(n386), .ZN(n366) );
  AND2_X1 U365 ( .A1(n558), .A2(n557), .ZN(n389) );
  XNOR2_X1 U366 ( .A(n390), .B(n538), .ZN(n559) );
  XNOR2_X1 U367 ( .A(n603), .B(n602), .ZN(n695) );
  XNOR2_X1 U368 ( .A(n578), .B(KEYINPUT38), .ZN(n697) );
  AND2_X1 U369 ( .A1(n383), .A2(n532), .ZN(n604) );
  XNOR2_X1 U370 ( .A(n357), .B(n440), .ZN(n552) );
  AND2_X1 U371 ( .A1(n403), .A2(n402), .ZN(n401) );
  NAND2_X1 U372 ( .A1(n555), .A2(n580), .ZN(n384) );
  XNOR2_X2 U373 ( .A(n677), .B(KEYINPUT104), .ZN(n555) );
  NAND2_X1 U374 ( .A1(n343), .A2(n593), .ZN(n396) );
  INV_X1 U375 ( .A(n344), .ZN(n343) );
  NAND2_X1 U376 ( .A1(n630), .A2(KEYINPUT72), .ZN(n344) );
  AND2_X2 U377 ( .A1(n567), .A2(n520), .ZN(n521) );
  XNOR2_X2 U378 ( .A(n519), .B(KEYINPUT92), .ZN(n567) );
  XNOR2_X2 U379 ( .A(G101), .B(G119), .ZN(n421) );
  NOR2_X1 U380 ( .A1(G953), .A2(G237), .ZN(n491) );
  INV_X1 U381 ( .A(G953), .ZN(n359) );
  AND2_X2 U382 ( .A1(n532), .A2(n353), .ZN(n519) );
  NAND2_X2 U383 ( .A1(n381), .A2(n373), .ZN(n649) );
  NAND2_X4 U384 ( .A1(n401), .A2(n398), .ZN(n677) );
  XNOR2_X2 U385 ( .A(n467), .B(n430), .ZN(n631) );
  INV_X1 U386 ( .A(n649), .ZN(n639) );
  AND2_X1 U387 ( .A1(n379), .A2(n620), .ZN(n373) );
  NAND2_X1 U388 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U389 ( .A1(n414), .A2(n412), .ZN(n746) );
  OR2_X1 U390 ( .A1(n584), .A2(n486), .ZN(n611) );
  XNOR2_X1 U391 ( .A(n482), .B(KEYINPUT87), .ZN(n483) );
  XNOR2_X1 U392 ( .A(n441), .B(G902), .ZN(n620) );
  XNOR2_X2 U393 ( .A(G116), .B(KEYINPUT3), .ZN(n422) );
  INV_X1 U394 ( .A(n389), .ZN(n385) );
  NOR2_X1 U395 ( .A1(n389), .A2(n388), .ZN(n387) );
  XNOR2_X1 U396 ( .A(G134), .B(G131), .ZN(n418) );
  OR2_X1 U397 ( .A1(n651), .A2(G902), .ZN(n468) );
  NAND2_X1 U398 ( .A1(n400), .A2(n513), .ZN(n399) );
  XNOR2_X1 U399 ( .A(KEYINPUT86), .B(G110), .ZN(n464) );
  NAND2_X1 U400 ( .A1(n363), .A2(n365), .ZN(n379) );
  NAND2_X1 U401 ( .A1(n376), .A2(n382), .ZN(n381) );
  INV_X1 U402 ( .A(KEYINPUT2), .ZN(n382) );
  AND2_X1 U403 ( .A1(n365), .A2(n577), .ZN(n377) );
  INV_X1 U404 ( .A(KEYINPUT34), .ZN(n374) );
  OR2_X1 U405 ( .A1(n579), .A2(n348), .ZN(n413) );
  NAND2_X1 U406 ( .A1(n416), .A2(n348), .ZN(n415) );
  XNOR2_X1 U407 ( .A(n409), .B(n408), .ZN(n407) );
  INV_X1 U408 ( .A(KEYINPUT30), .ZN(n408) );
  XNOR2_X1 U409 ( .A(n446), .B(n439), .ZN(n357) );
  NAND2_X1 U410 ( .A1(n381), .A2(n379), .ZN(n361) );
  AND2_X1 U411 ( .A1(n598), .A2(n397), .ZN(n395) );
  NAND2_X1 U412 ( .A1(KEYINPUT47), .A2(KEYINPUT72), .ZN(n397) );
  INV_X1 U413 ( .A(KEYINPUT44), .ZN(n388) );
  INV_X1 U414 ( .A(KEYINPUT69), .ZN(n420) );
  INV_X1 U415 ( .A(G237), .ZN(n481) );
  INV_X1 U416 ( .A(G472), .ZN(n400) );
  NAND2_X1 U417 ( .A1(G902), .A2(G472), .ZN(n402) );
  XNOR2_X1 U418 ( .A(G119), .B(G128), .ZN(n431) );
  XOR2_X1 U419 ( .A(G122), .B(G107), .Z(n503) );
  NAND2_X1 U420 ( .A1(G234), .A2(G237), .ZN(n447) );
  NAND2_X1 U421 ( .A1(n555), .A2(n696), .ZN(n409) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n410) );
  INV_X1 U423 ( .A(KEYINPUT19), .ZN(n355) );
  NOR2_X1 U424 ( .A1(n578), .A2(n486), .ZN(n356) );
  BUF_X1 U425 ( .A(n469), .Z(n429) );
  XOR2_X1 U426 ( .A(G104), .B(G122), .Z(n488) );
  XNOR2_X1 U427 ( .A(G113), .B(G143), .ZN(n487) );
  XOR2_X1 U428 ( .A(KEYINPUT11), .B(KEYINPUT95), .Z(n495) );
  XOR2_X1 U429 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n493) );
  XNOR2_X1 U430 ( .A(n537), .B(n536), .ZN(n709) );
  XNOR2_X1 U431 ( .A(n384), .B(n459), .ZN(n383) );
  NAND2_X1 U432 ( .A1(n695), .A2(n699), .ZN(n405) );
  AND2_X2 U433 ( .A1(n410), .A2(n604), .ZN(n595) );
  XNOR2_X1 U434 ( .A(n358), .B(n438), .ZN(n720) );
  XNOR2_X1 U435 ( .A(n437), .B(n436), .ZN(n358) );
  XNOR2_X1 U436 ( .A(n467), .B(n466), .ZN(n651) );
  XNOR2_X1 U437 ( .A(n627), .B(KEYINPUT85), .ZN(n722) );
  INV_X1 U438 ( .A(n587), .ZN(n391) );
  AND2_X1 U439 ( .A1(n411), .A2(n415), .ZN(n414) );
  XNOR2_X1 U440 ( .A(n360), .B(KEYINPUT122), .ZN(n713) );
  NAND2_X1 U441 ( .A1(n361), .A2(n346), .ZN(n360) );
  XNOR2_X1 U442 ( .A(n389), .B(n372), .ZN(G12) );
  INV_X1 U443 ( .A(G110), .ZN(n372) );
  XNOR2_X1 U444 ( .A(G146), .B(G125), .ZN(n473) );
  XOR2_X1 U445 ( .A(KEYINPUT23), .B(G110), .Z(n345) );
  NOR2_X1 U446 ( .A1(n712), .A2(n711), .ZN(n346) );
  OR2_X1 U447 ( .A1(n417), .A2(n413), .ZN(n347) );
  XNOR2_X1 U448 ( .A(KEYINPUT75), .B(KEYINPUT32), .ZN(n348) );
  XOR2_X1 U449 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n349) );
  XOR2_X1 U450 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n350) );
  AND2_X1 U451 ( .A1(n577), .A2(KEYINPUT2), .ZN(n351) );
  NAND2_X1 U452 ( .A1(n454), .A2(G217), .ZN(n444) );
  XNOR2_X1 U453 ( .A(n443), .B(KEYINPUT20), .ZN(n454) );
  XNOR2_X1 U454 ( .A(n523), .B(KEYINPUT39), .ZN(n542) );
  INV_X1 U455 ( .A(n684), .ZN(n353) );
  NOR2_X2 U456 ( .A1(n620), .A2(n640), .ZN(n484) );
  XNOR2_X2 U457 ( .A(n468), .B(G469), .ZN(n532) );
  BUF_X1 U458 ( .A(n559), .Z(n354) );
  AND2_X1 U459 ( .A1(n601), .A2(n671), .ZN(n608) );
  NAND2_X1 U460 ( .A1(n362), .A2(n351), .ZN(n364) );
  NAND2_X1 U461 ( .A1(n364), .A2(n380), .ZN(n363) );
  AND2_X1 U462 ( .A1(n365), .A2(n359), .ZN(n727) );
  XNOR2_X2 U463 ( .A(n576), .B(n349), .ZN(n365) );
  INV_X1 U464 ( .A(n619), .ZN(n362) );
  NAND2_X1 U465 ( .A1(n366), .A2(n368), .ZN(n575) );
  NAND2_X1 U466 ( .A1(n369), .A2(n388), .ZN(n367) );
  NAND2_X1 U467 ( .A1(n370), .A2(n387), .ZN(n368) );
  NAND2_X1 U468 ( .A1(n371), .A2(n385), .ZN(n369) );
  NOR2_X1 U469 ( .A1(n746), .A2(n559), .ZN(n370) );
  INV_X1 U470 ( .A(n559), .ZN(n371) );
  XNOR2_X1 U471 ( .A(n375), .B(n374), .ZN(n392) );
  NAND2_X1 U472 ( .A1(n569), .A2(n709), .ZN(n375) );
  XNOR2_X2 U473 ( .A(n393), .B(n530), .ZN(n569) );
  NAND2_X1 U474 ( .A1(n378), .A2(n377), .ZN(n376) );
  INV_X1 U475 ( .A(n734), .ZN(n378) );
  XNOR2_X1 U476 ( .A(n619), .B(KEYINPUT78), .ZN(n734) );
  NAND2_X1 U477 ( .A1(n619), .A2(KEYINPUT79), .ZN(n380) );
  NAND2_X1 U478 ( .A1(n746), .A2(n388), .ZN(n386) );
  NAND2_X1 U479 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U480 ( .A1(n410), .A2(n529), .ZN(n393) );
  NAND2_X1 U481 ( .A1(n599), .A2(n394), .ZN(n600) );
  NAND2_X1 U482 ( .A1(n396), .A2(n395), .ZN(n394) );
  OR2_X1 U483 ( .A1(n631), .A2(n399), .ZN(n398) );
  NAND2_X1 U484 ( .A1(n631), .A2(G472), .ZN(n403) );
  XNOR2_X2 U485 ( .A(n404), .B(KEYINPUT42), .ZN(n747) );
  NAND2_X1 U486 ( .A1(n710), .A2(n604), .ZN(n404) );
  XNOR2_X2 U487 ( .A(n405), .B(KEYINPUT41), .ZN(n710) );
  XNOR2_X2 U488 ( .A(n406), .B(G143), .ZN(n509) );
  XNOR2_X2 U489 ( .A(G128), .B(KEYINPUT76), .ZN(n406) );
  INV_X1 U490 ( .A(n589), .ZN(n522) );
  NAND2_X1 U491 ( .A1(n521), .A2(n407), .ZN(n589) );
  OR2_X1 U492 ( .A1(n554), .A2(n347), .ZN(n412) );
  XNOR2_X2 U493 ( .A(n551), .B(KEYINPUT22), .ZN(n554) );
  NAND2_X1 U494 ( .A1(n554), .A2(n348), .ZN(n411) );
  NOR2_X1 U495 ( .A1(n554), .A2(n579), .ZN(n560) );
  NAND2_X1 U496 ( .A1(n553), .A2(n582), .ZN(n416) );
  INV_X1 U497 ( .A(n553), .ZN(n417) );
  BUF_X1 U498 ( .A(n578), .Z(n614) );
  XNOR2_X2 U499 ( .A(n509), .B(KEYINPUT4), .ZN(n477) );
  XNOR2_X1 U500 ( .A(n472), .B(n471), .ZN(n723) );
  INV_X1 U501 ( .A(n473), .ZN(n474) );
  INV_X1 U502 ( .A(KEYINPUT89), .ZN(n432) );
  INV_X1 U503 ( .A(KEYINPUT110), .ZN(n602) );
  XNOR2_X1 U504 ( .A(n432), .B(KEYINPUT24), .ZN(n433) );
  XNOR2_X1 U505 ( .A(n434), .B(n433), .ZN(n437) );
  BUF_X1 U506 ( .A(n723), .Z(n724) );
  INV_X1 U507 ( .A(n735), .ZN(n438) );
  XNOR2_X1 U508 ( .A(n512), .B(n511), .ZN(n716) );
  XNOR2_X1 U509 ( .A(n418), .B(KEYINPUT67), .ZN(n419) );
  XNOR2_X2 U510 ( .A(n477), .B(n419), .ZN(n736) );
  XNOR2_X2 U511 ( .A(n736), .B(G146), .ZN(n467) );
  XNOR2_X1 U512 ( .A(n421), .B(n420), .ZN(n424) );
  XNOR2_X1 U513 ( .A(n422), .B(G113), .ZN(n423) );
  XNOR2_X1 U514 ( .A(n424), .B(n423), .ZN(n469) );
  NAND2_X1 U515 ( .A1(n491), .A2(G210), .ZN(n425) );
  XNOR2_X1 U516 ( .A(n425), .B(KEYINPUT5), .ZN(n427) );
  XNOR2_X1 U517 ( .A(G137), .B(KEYINPUT93), .ZN(n426) );
  XNOR2_X1 U518 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U519 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U520 ( .A(n345), .B(n431), .ZN(n434) );
  NAND2_X1 U521 ( .A1(G234), .A2(n359), .ZN(n435) );
  XOR2_X1 U522 ( .A(KEYINPUT8), .B(n435), .Z(n504) );
  NAND2_X1 U523 ( .A1(n504), .A2(G221), .ZN(n436) );
  XNOR2_X1 U524 ( .A(n473), .B(KEYINPUT10), .ZN(n490) );
  XNOR2_X1 U525 ( .A(G137), .B(G140), .ZN(n462) );
  XNOR2_X1 U526 ( .A(n490), .B(n462), .ZN(n735) );
  NOR2_X1 U527 ( .A1(G902), .A2(n720), .ZN(n440) );
  XNOR2_X1 U528 ( .A(KEYINPUT90), .B(KEYINPUT25), .ZN(n439) );
  XOR2_X1 U529 ( .A(KEYINPUT91), .B(KEYINPUT73), .Z(n445) );
  INV_X1 U530 ( .A(KEYINPUT15), .ZN(n441) );
  INV_X1 U531 ( .A(n620), .ZN(n442) );
  NAND2_X1 U532 ( .A1(G234), .A2(n442), .ZN(n443) );
  XNOR2_X1 U533 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U534 ( .A(n447), .B(KEYINPUT14), .ZN(n451) );
  AND2_X1 U535 ( .A1(G953), .A2(G902), .ZN(n448) );
  NAND2_X1 U536 ( .A1(n451), .A2(n448), .ZN(n525) );
  XOR2_X1 U537 ( .A(KEYINPUT105), .B(n525), .Z(n449) );
  NOR2_X1 U538 ( .A1(G900), .A2(n449), .ZN(n450) );
  XNOR2_X1 U539 ( .A(n450), .B(KEYINPUT106), .ZN(n452) );
  NAND2_X1 U540 ( .A1(G952), .A2(n451), .ZN(n708) );
  NOR2_X1 U541 ( .A1(G953), .A2(n708), .ZN(n528) );
  NOR2_X1 U542 ( .A1(n452), .A2(n528), .ZN(n453) );
  XNOR2_X1 U543 ( .A(n453), .B(KEYINPUT77), .ZN(n520) );
  NAND2_X1 U544 ( .A1(n454), .A2(G221), .ZN(n455) );
  XNOR2_X1 U545 ( .A(n455), .B(KEYINPUT21), .ZN(n675) );
  INV_X1 U546 ( .A(n675), .ZN(n456) );
  AND2_X1 U547 ( .A1(n520), .A2(n456), .ZN(n457) );
  XNOR2_X1 U548 ( .A(n457), .B(KEYINPUT68), .ZN(n458) );
  AND2_X1 U549 ( .A1(n552), .A2(n458), .ZN(n580) );
  INV_X1 U550 ( .A(KEYINPUT28), .ZN(n459) );
  XNOR2_X1 U551 ( .A(G101), .B(G107), .ZN(n461) );
  NAND2_X1 U552 ( .A1(n359), .A2(G227), .ZN(n460) );
  XNOR2_X1 U553 ( .A(n461), .B(n460), .ZN(n463) );
  XNOR2_X1 U554 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X1 U555 ( .A(n464), .B(G104), .ZN(n470) );
  XNOR2_X1 U556 ( .A(n465), .B(n470), .ZN(n466) );
  XNOR2_X1 U557 ( .A(n469), .B(n503), .ZN(n472) );
  XOR2_X1 U558 ( .A(n470), .B(KEYINPUT16), .Z(n471) );
  XNOR2_X1 U559 ( .A(n723), .B(KEYINPUT17), .ZN(n480) );
  NAND2_X1 U560 ( .A1(G224), .A2(n359), .ZN(n475) );
  XNOR2_X1 U561 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U562 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U563 ( .A(n478), .B(KEYINPUT18), .Z(n479) );
  XNOR2_X1 U564 ( .A(n480), .B(n479), .ZN(n640) );
  INV_X1 U565 ( .A(G902), .ZN(n513) );
  NAND2_X1 U566 ( .A1(n513), .A2(n481), .ZN(n485) );
  NAND2_X1 U567 ( .A1(G210), .A2(n485), .ZN(n482) );
  XNOR2_X2 U568 ( .A(n484), .B(n483), .ZN(n578) );
  NAND2_X1 U569 ( .A1(n485), .A2(G214), .ZN(n696) );
  INV_X1 U570 ( .A(n696), .ZN(n486) );
  XNOR2_X1 U571 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n501) );
  XNOR2_X1 U572 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U573 ( .A(n490), .B(n489), .ZN(n499) );
  NAND2_X1 U574 ( .A1(G214), .A2(n491), .ZN(n492) );
  XNOR2_X1 U575 ( .A(n493), .B(n492), .ZN(n497) );
  XNOR2_X1 U576 ( .A(G131), .B(G140), .ZN(n494) );
  XNOR2_X1 U577 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U578 ( .A(n497), .B(n496), .Z(n498) );
  XNOR2_X1 U579 ( .A(n499), .B(n498), .ZN(n623) );
  NOR2_X1 U580 ( .A1(G902), .A2(n623), .ZN(n500) );
  XNOR2_X1 U581 ( .A(n501), .B(n500), .ZN(n502) );
  INV_X1 U582 ( .A(G475), .ZN(n621) );
  XNOR2_X1 U583 ( .A(n502), .B(n621), .ZN(n547) );
  XOR2_X1 U584 ( .A(G134), .B(n503), .Z(n506) );
  NAND2_X1 U585 ( .A1(G217), .A2(n504), .ZN(n505) );
  XNOR2_X1 U586 ( .A(n506), .B(n505), .ZN(n512) );
  XOR2_X1 U587 ( .A(KEYINPUT9), .B(KEYINPUT98), .Z(n508) );
  XNOR2_X1 U588 ( .A(G116), .B(KEYINPUT7), .ZN(n507) );
  XNOR2_X1 U589 ( .A(n508), .B(n507), .ZN(n510) );
  XNOR2_X1 U590 ( .A(n509), .B(n510), .ZN(n511) );
  NAND2_X1 U591 ( .A1(n716), .A2(n513), .ZN(n515) );
  XOR2_X1 U592 ( .A(KEYINPUT99), .B(G478), .Z(n514) );
  XNOR2_X1 U593 ( .A(n515), .B(n514), .ZN(n546) );
  INV_X1 U594 ( .A(n546), .ZN(n539) );
  OR2_X1 U595 ( .A1(n547), .A2(n539), .ZN(n516) );
  XNOR2_X1 U596 ( .A(n516), .B(KEYINPUT101), .ZN(n666) );
  NAND2_X1 U597 ( .A1(n595), .A2(n666), .ZN(n593) );
  XOR2_X1 U598 ( .A(KEYINPUT29), .B(KEYINPUT115), .Z(n517) );
  XOR2_X1 U599 ( .A(n517), .B(G128), .Z(n518) );
  XNOR2_X1 U600 ( .A(n593), .B(n518), .ZN(G30) );
  XNOR2_X1 U601 ( .A(G134), .B(KEYINPUT118), .ZN(n524) );
  OR2_X2 U602 ( .A1(n552), .A2(n675), .ZN(n684) );
  NAND2_X1 U603 ( .A1(n522), .A2(n697), .ZN(n523) );
  AND2_X1 U604 ( .A1(n542), .A2(n666), .ZN(n616) );
  XOR2_X1 U605 ( .A(n524), .B(n616), .Z(G36) );
  NOR2_X1 U606 ( .A1(G898), .A2(n525), .ZN(n526) );
  XNOR2_X1 U607 ( .A(n526), .B(KEYINPUT88), .ZN(n527) );
  OR2_X1 U608 ( .A1(n528), .A2(n527), .ZN(n529) );
  INV_X1 U609 ( .A(KEYINPUT0), .ZN(n530) );
  INV_X1 U610 ( .A(KEYINPUT1), .ZN(n531) );
  XNOR2_X2 U611 ( .A(n532), .B(n531), .ZN(n683) );
  NOR2_X1 U612 ( .A1(n684), .A2(n683), .ZN(n534) );
  INV_X1 U613 ( .A(KEYINPUT6), .ZN(n533) );
  XNOR2_X1 U614 ( .A(n677), .B(n533), .ZN(n579) );
  NAND2_X1 U615 ( .A1(n534), .A2(n579), .ZN(n537) );
  XNOR2_X1 U616 ( .A(KEYINPUT82), .B(KEYINPUT33), .ZN(n535) );
  XNOR2_X1 U617 ( .A(n535), .B(KEYINPUT70), .ZN(n536) );
  NAND2_X1 U618 ( .A1(n547), .A2(n546), .ZN(n587) );
  XNOR2_X1 U619 ( .A(KEYINPUT74), .B(KEYINPUT35), .ZN(n538) );
  XOR2_X1 U620 ( .A(n354), .B(G122), .Z(G24) );
  NAND2_X1 U621 ( .A1(n539), .A2(n547), .ZN(n541) );
  INV_X1 U622 ( .A(KEYINPUT100), .ZN(n540) );
  XNOR2_X2 U623 ( .A(n541), .B(n540), .ZN(n664) );
  NAND2_X1 U624 ( .A1(n542), .A2(n664), .ZN(n545) );
  INV_X1 U625 ( .A(KEYINPUT109), .ZN(n543) );
  XNOR2_X1 U626 ( .A(n543), .B(KEYINPUT40), .ZN(n544) );
  XNOR2_X2 U627 ( .A(n545), .B(n544), .ZN(n605) );
  XNOR2_X1 U628 ( .A(n605), .B(G131), .ZN(G33) );
  NOR2_X1 U629 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U630 ( .A(n548), .B(KEYINPUT102), .ZN(n699) );
  INV_X1 U631 ( .A(n699), .ZN(n549) );
  NOR2_X1 U632 ( .A1(n675), .A2(n549), .ZN(n550) );
  NAND2_X1 U633 ( .A1(n569), .A2(n550), .ZN(n551) );
  INV_X1 U634 ( .A(n552), .ZN(n561) );
  NOR2_X1 U635 ( .A1(n561), .A2(n683), .ZN(n553) );
  INV_X1 U636 ( .A(n554), .ZN(n558) );
  NAND2_X1 U637 ( .A1(n683), .A2(n552), .ZN(n556) );
  NOR2_X1 U638 ( .A1(n556), .A2(n555), .ZN(n557) );
  AND2_X1 U639 ( .A1(n561), .A2(n683), .ZN(n562) );
  NAND2_X1 U640 ( .A1(n560), .A2(n562), .ZN(n563) );
  XNOR2_X1 U641 ( .A(n563), .B(KEYINPUT103), .ZN(n745) );
  INV_X1 U642 ( .A(n677), .ZN(n566) );
  NOR2_X1 U643 ( .A1(n684), .A2(n566), .ZN(n564) );
  INV_X1 U644 ( .A(n683), .ZN(n681) );
  AND2_X1 U645 ( .A1(n564), .A2(n681), .ZN(n690) );
  NAND2_X1 U646 ( .A1(n569), .A2(n690), .ZN(n565) );
  XNOR2_X1 U647 ( .A(KEYINPUT31), .B(n565), .ZN(n667) );
  AND2_X1 U648 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U649 ( .A1(n569), .A2(n568), .ZN(n571) );
  INV_X1 U650 ( .A(KEYINPUT94), .ZN(n570) );
  XNOR2_X1 U651 ( .A(n571), .B(n570), .ZN(n656) );
  NOR2_X1 U652 ( .A1(n667), .A2(n656), .ZN(n572) );
  OR2_X1 U653 ( .A1(n666), .A2(n664), .ZN(n694) );
  INV_X1 U654 ( .A(n694), .ZN(n594) );
  NOR2_X1 U655 ( .A1(n572), .A2(n594), .ZN(n573) );
  NOR2_X1 U656 ( .A1(n745), .A2(n573), .ZN(n574) );
  NAND2_X1 U657 ( .A1(n575), .A2(n574), .ZN(n576) );
  INV_X1 U658 ( .A(KEYINPUT79), .ZN(n577) );
  INV_X1 U659 ( .A(n579), .ZN(n582) );
  NAND2_X1 U660 ( .A1(n580), .A2(n664), .ZN(n581) );
  NOR2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U662 ( .A(n583), .B(KEYINPUT107), .ZN(n584) );
  NOR2_X1 U663 ( .A1(n614), .A2(n611), .ZN(n585) );
  XNOR2_X1 U664 ( .A(n585), .B(KEYINPUT36), .ZN(n586) );
  NAND2_X1 U665 ( .A1(n586), .A2(n681), .ZN(n671) );
  OR2_X1 U666 ( .A1(n614), .A2(n587), .ZN(n588) );
  NOR2_X1 U667 ( .A1(n589), .A2(n588), .ZN(n663) );
  AND2_X1 U668 ( .A1(n694), .A2(KEYINPUT72), .ZN(n590) );
  NAND2_X1 U669 ( .A1(n595), .A2(n590), .ZN(n591) );
  AND2_X1 U670 ( .A1(n591), .A2(KEYINPUT47), .ZN(n592) );
  NOR2_X1 U671 ( .A1(n663), .A2(n592), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n595), .A2(n664), .ZN(n630) );
  NAND2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n597) );
  INV_X1 U674 ( .A(KEYINPUT72), .ZN(n596) );
  NAND2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U676 ( .A(n600), .B(KEYINPUT71), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n697), .A2(n696), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n605), .A2(n747), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(n350), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n610) );
  XNOR2_X1 U681 ( .A(KEYINPUT81), .B(KEYINPUT48), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n610), .B(n609), .ZN(n618) );
  XOR2_X1 U683 ( .A(KEYINPUT108), .B(n611), .Z(n612) );
  NAND2_X1 U684 ( .A1(n612), .A2(n683), .ZN(n613) );
  XNOR2_X1 U685 ( .A(n613), .B(KEYINPUT43), .ZN(n615) );
  AND2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n673) );
  NOR2_X1 U687 ( .A1(n673), .A2(n616), .ZN(n617) );
  NOR2_X1 U688 ( .A1(n649), .A2(n621), .ZN(n625) );
  XNOR2_X1 U689 ( .A(KEYINPUT66), .B(KEYINPUT59), .ZN(n622) );
  XNOR2_X1 U690 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U691 ( .A(n625), .B(n624), .ZN(n628) );
  INV_X1 U692 ( .A(G952), .ZN(n626) );
  NAND2_X1 U693 ( .A1(n626), .A2(G953), .ZN(n627) );
  NOR2_X1 U694 ( .A1(n628), .A2(n722), .ZN(n629) );
  XNOR2_X1 U695 ( .A(n629), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U696 ( .A(n630), .B(G146), .ZN(G48) );
  NAND2_X1 U697 ( .A1(n639), .A2(G472), .ZN(n635) );
  XNOR2_X1 U698 ( .A(KEYINPUT83), .B(KEYINPUT111), .ZN(n632) );
  XNOR2_X1 U699 ( .A(n632), .B(KEYINPUT62), .ZN(n633) );
  XNOR2_X1 U700 ( .A(n631), .B(n633), .ZN(n634) );
  XNOR2_X1 U701 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X2 U702 ( .A1(n636), .A2(n722), .ZN(n638) );
  XOR2_X1 U703 ( .A(KEYINPUT84), .B(KEYINPUT63), .Z(n637) );
  XNOR2_X1 U704 ( .A(n638), .B(n637), .ZN(G57) );
  NAND2_X1 U705 ( .A1(n639), .A2(G210), .ZN(n645) );
  BUF_X1 U706 ( .A(n640), .Z(n641) );
  XNOR2_X1 U707 ( .A(KEYINPUT123), .B(KEYINPUT54), .ZN(n642) );
  XNOR2_X1 U708 ( .A(n642), .B(KEYINPUT55), .ZN(n643) );
  XNOR2_X1 U709 ( .A(n641), .B(n643), .ZN(n644) );
  XNOR2_X1 U710 ( .A(n645), .B(n644), .ZN(n646) );
  NOR2_X2 U711 ( .A1(n646), .A2(n722), .ZN(n648) );
  XNOR2_X1 U712 ( .A(KEYINPUT80), .B(KEYINPUT56), .ZN(n647) );
  XNOR2_X1 U713 ( .A(n648), .B(n647), .ZN(G51) );
  INV_X1 U714 ( .A(n649), .ZN(n718) );
  NAND2_X1 U715 ( .A1(n718), .A2(G469), .ZN(n653) );
  XOR2_X1 U716 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n650) );
  XNOR2_X1 U717 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U718 ( .A(n653), .B(n652), .ZN(n654) );
  NOR2_X1 U719 ( .A1(n654), .A2(n722), .ZN(G54) );
  NAND2_X1 U720 ( .A1(n656), .A2(n664), .ZN(n655) );
  XNOR2_X1 U721 ( .A(n655), .B(G104), .ZN(G6) );
  NAND2_X1 U722 ( .A1(n656), .A2(n666), .ZN(n662) );
  XOR2_X1 U723 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n658) );
  XNOR2_X1 U724 ( .A(KEYINPUT112), .B(KEYINPUT27), .ZN(n657) );
  XNOR2_X1 U725 ( .A(n658), .B(n657), .ZN(n660) );
  XOR2_X1 U726 ( .A(G107), .B(KEYINPUT26), .Z(n659) );
  XNOR2_X1 U727 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U728 ( .A(n662), .B(n661), .ZN(G9) );
  XOR2_X1 U729 ( .A(G143), .B(n663), .Z(G45) );
  NAND2_X1 U730 ( .A1(n664), .A2(n667), .ZN(n665) );
  XNOR2_X1 U731 ( .A(n665), .B(G113), .ZN(G15) );
  XOR2_X1 U732 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n669) );
  NAND2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U734 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U735 ( .A(G116), .B(n670), .ZN(G18) );
  XOR2_X1 U736 ( .A(G125), .B(n671), .Z(n672) );
  XNOR2_X1 U737 ( .A(n672), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U738 ( .A(G140), .B(n673), .ZN(n674) );
  XNOR2_X1 U739 ( .A(n674), .B(KEYINPUT119), .ZN(G42) );
  NAND2_X1 U740 ( .A1(n675), .A2(n552), .ZN(n676) );
  XNOR2_X1 U741 ( .A(KEYINPUT49), .B(n676), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U743 ( .A(KEYINPUT120), .B(n679), .Z(n689) );
  INV_X1 U744 ( .A(KEYINPUT50), .ZN(n680) );
  NAND2_X1 U745 ( .A1(n684), .A2(n680), .ZN(n682) );
  NOR2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n687) );
  NAND2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n685) );
  AND2_X1 U748 ( .A1(n685), .A2(KEYINPUT50), .ZN(n686) );
  NOR2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n689), .A2(n688), .ZN(n691) );
  NOR2_X1 U751 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U752 ( .A(n692), .B(KEYINPUT51), .ZN(n693) );
  NAND2_X1 U753 ( .A1(n693), .A2(n710), .ZN(n705) );
  NAND2_X1 U754 ( .A1(n695), .A2(n694), .ZN(n702) );
  NOR2_X1 U755 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U756 ( .A(n698), .B(KEYINPUT121), .ZN(n700) );
  NAND2_X1 U757 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U758 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U759 ( .A1(n703), .A2(n709), .ZN(n704) );
  NAND2_X1 U760 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U761 ( .A(KEYINPUT52), .B(n706), .Z(n707) );
  NOR2_X1 U762 ( .A1(n708), .A2(n707), .ZN(n712) );
  AND2_X1 U763 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n713), .A2(G953), .ZN(n714) );
  XNOR2_X1 U765 ( .A(n714), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U766 ( .A1(n718), .A2(G478), .ZN(n715) );
  XOR2_X1 U767 ( .A(n716), .B(n715), .Z(n717) );
  NOR2_X1 U768 ( .A1(n722), .A2(n717), .ZN(G63) );
  NAND2_X1 U769 ( .A1(n718), .A2(G217), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U771 ( .A1(n722), .A2(n721), .ZN(G66) );
  NOR2_X1 U772 ( .A1(G898), .A2(n359), .ZN(n726) );
  XOR2_X1 U773 ( .A(n724), .B(KEYINPUT125), .Z(n725) );
  NOR2_X1 U774 ( .A1(n726), .A2(n725), .ZN(n733) );
  XOR2_X1 U775 ( .A(KEYINPUT124), .B(n727), .Z(n731) );
  NAND2_X1 U776 ( .A1(G953), .A2(G224), .ZN(n728) );
  XNOR2_X1 U777 ( .A(KEYINPUT61), .B(n728), .ZN(n729) );
  NAND2_X1 U778 ( .A1(n729), .A2(G898), .ZN(n730) );
  NAND2_X1 U779 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U780 ( .A(n733), .B(n732), .ZN(G69) );
  XNOR2_X1 U781 ( .A(n736), .B(n735), .ZN(n739) );
  XNOR2_X1 U782 ( .A(n734), .B(n739), .ZN(n737) );
  NAND2_X1 U783 ( .A1(n737), .A2(n359), .ZN(n738) );
  XNOR2_X1 U784 ( .A(KEYINPUT126), .B(n738), .ZN(n744) );
  XNOR2_X1 U785 ( .A(n739), .B(G227), .ZN(n740) );
  NAND2_X1 U786 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U787 ( .A1(G953), .A2(n741), .ZN(n742) );
  XOR2_X1 U788 ( .A(KEYINPUT127), .B(n742), .Z(n743) );
  NAND2_X1 U789 ( .A1(n744), .A2(n743), .ZN(G72) );
  XOR2_X1 U790 ( .A(G101), .B(n745), .Z(G3) );
  XOR2_X1 U791 ( .A(n746), .B(G119), .Z(G21) );
  XNOR2_X1 U792 ( .A(n747), .B(G137), .ZN(G39) );
endmodule

