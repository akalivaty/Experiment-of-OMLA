//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n202));
  OR2_X1    g001(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(G190gat), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(G169gat), .A3(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G169gat), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n205), .A2(new_n210), .A3(new_n212), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G176gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT23), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G169gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n202), .B1(new_n218), .B2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  OAI22_X1  g028(.A1(new_n229), .A2(KEYINPUT23), .B1(new_n204), .B2(G190gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n230), .B1(new_n207), .B2(new_n209), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT67), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n234), .A3(KEYINPUT23), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n231), .A2(KEYINPUT25), .A3(new_n205), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n228), .A2(new_n236), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n207), .A2(new_n209), .B1(new_n215), .B2(KEYINPUT26), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n232), .A2(new_n234), .A3(new_n239), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n238), .A2(new_n240), .B1(G183gat), .B2(G190gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT27), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n244), .A2(G183gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(G183gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n243), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(G183gat), .ZN(new_n248));
  AOI21_X1  g047(.A(G190gat), .B1(new_n248), .B2(KEYINPUT68), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT28), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT27), .B(G183gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT28), .A3(new_n211), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI22_X1  g052(.A1(new_n241), .A2(new_n242), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n215), .A2(KEYINPUT26), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n210), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(KEYINPUT69), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n237), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G127gat), .B(G134gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263));
  INV_X1    g062(.A(G127gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(G134gat), .ZN(new_n265));
  INV_X1    g064(.A(G134gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(G127gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n263), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G113gat), .ZN(new_n270));
  INV_X1    g069(.A(G120gat), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(new_n270), .B2(new_n271), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n261), .A2(new_n272), .ZN(new_n274));
  XOR2_X1   g073(.A(KEYINPUT71), .B(G120gat), .Z(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G113gat), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n269), .A2(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G227gat), .ZN(new_n279));
  INV_X1    g078(.A(G233gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n258), .A2(KEYINPUT69), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n211), .B1(new_n245), .B2(new_n243), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n252), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n241), .A2(new_n242), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n282), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n269), .A2(new_n273), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n276), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n292), .A3(new_n237), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n278), .A2(new_n281), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT32), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT33), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G71gat), .B(G99gat), .Z(new_n298));
  XNOR2_X1  g097(.A(G15gat), .B(G43gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n295), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT72), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(KEYINPUT33), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n294), .A2(KEYINPUT32), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT73), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n294), .A2(new_n306), .A3(KEYINPUT32), .A4(new_n303), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n295), .A2(new_n297), .A3(new_n309), .A4(new_n300), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n302), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT34), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n278), .A2(new_n293), .ZN(new_n313));
  INV_X1    g112(.A(new_n281), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI211_X1 g114(.A(KEYINPUT34), .B(new_n281), .C1(new_n278), .C2(new_n293), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n311), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n302), .A2(new_n308), .A3(new_n317), .A4(new_n310), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT36), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n311), .A2(KEYINPUT74), .A3(new_n318), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n319), .A2(KEYINPUT36), .A3(new_n321), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G155gat), .B(G162gat), .ZN(new_n328));
  OR2_X1    g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n334));
  OAI21_X1  g133(.A(G155gat), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT2), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n331), .B1(new_n336), .B2(KEYINPUT78), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n338), .A3(KEYINPUT2), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n329), .A2(new_n340), .A3(new_n330), .ZN(new_n341));
  INV_X1    g140(.A(new_n328), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n337), .A2(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G211gat), .B(G218gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT76), .B(G211gat), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT22), .B1(new_n346), .B2(G218gat), .ZN(new_n347));
  INV_X1    g146(.A(G204gat), .ZN(new_n348));
  AND2_X1   g147(.A1(KEYINPUT75), .A2(G197gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(KEYINPUT75), .A2(G197gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n352));
  INV_X1    g151(.A(G197gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(KEYINPUT75), .A2(G197gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(G204gat), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n345), .B1(new_n347), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n360));
  OAI21_X1  g159(.A(G218gat), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT22), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n363), .A2(new_n356), .A3(new_n351), .A4(new_n344), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n343), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G155gat), .ZN(new_n370));
  OR2_X1    g169(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n370), .B1(new_n371), .B2(new_n332), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT78), .B1(new_n372), .B2(new_n340), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n339), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n342), .A2(new_n341), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n368), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n365), .B1(new_n377), .B2(new_n366), .ZN(new_n378));
  INV_X1    g177(.A(G228gat), .ZN(new_n379));
  OAI22_X1  g178(.A1(new_n369), .A2(new_n378), .B1(new_n379), .B2(new_n280), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT29), .B1(new_n343), .B2(new_n368), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT83), .B1(new_n383), .B2(new_n365), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n379), .A2(new_n280), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n368), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(new_n376), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n378), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n384), .A2(new_n385), .A3(new_n388), .A4(new_n390), .ZN(new_n391));
  OAI221_X1 g190(.A(KEYINPUT82), .B1(new_n379), .B2(new_n280), .C1(new_n369), .C2(new_n378), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n382), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT84), .B1(new_n393), .B2(G22gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(G50gat), .ZN(new_n396));
  XOR2_X1   g195(.A(G78gat), .B(G106gat), .Z(new_n397));
  XOR2_X1   g196(.A(new_n396), .B(new_n397), .Z(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(G22gat), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT3), .B1(new_n365), .B2(new_n366), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n385), .B1(new_n401), .B2(new_n343), .ZN(new_n402));
  AOI211_X1 g201(.A(KEYINPUT83), .B(new_n365), .C1(new_n377), .C2(new_n366), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n404), .A2(new_n384), .B1(new_n380), .B2(new_n381), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n400), .B1(new_n405), .B2(new_n392), .ZN(new_n406));
  AND4_X1   g205(.A1(new_n400), .A2(new_n382), .A3(new_n391), .A4(new_n392), .ZN(new_n407));
  OAI22_X1  g206(.A1(new_n394), .A2(new_n399), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n400), .A3(new_n392), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n393), .A2(G22gat), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT84), .A4(new_n398), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n365), .ZN(new_n413));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n237), .B(new_n414), .C1(new_n254), .C2(new_n259), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n289), .B2(new_n237), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n413), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(KEYINPUT69), .A2(new_n258), .B1(new_n286), .B2(new_n252), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n420), .A2(new_n288), .B1(new_n228), .B2(new_n236), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n365), .B(new_n415), .C1(new_n421), .C2(new_n417), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  NAND3_X1  g224(.A1(new_n419), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT37), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n419), .A2(new_n428), .A3(new_n422), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT85), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n419), .A2(new_n431), .A3(new_n422), .A4(new_n428), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n419), .A2(new_n422), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n425), .B1(new_n434), .B2(KEYINPUT37), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n427), .B1(new_n436), .B2(KEYINPUT38), .ZN(new_n437));
  XNOR2_X1  g236(.A(G1gat), .B(G29gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT0), .ZN(new_n439));
  XNOR2_X1  g238(.A(G57gat), .B(G85gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  NAND2_X1  g240(.A1(new_n377), .A2(new_n292), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n368), .B1(new_n375), .B2(new_n376), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT79), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n387), .A2(KEYINPUT3), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT79), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n292), .A4(new_n377), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G225gat), .A2(G233gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n277), .A2(new_n376), .A3(new_n375), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT4), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n343), .A2(KEYINPUT4), .A3(new_n277), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n448), .A2(new_n449), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n449), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n343), .A2(new_n277), .ZN(new_n458));
  INV_X1    g257(.A(new_n450), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT5), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n454), .B1(new_n444), .B2(new_n447), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT5), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n449), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n441), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT6), .ZN(new_n468));
  INV_X1    g267(.A(new_n441), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n456), .A2(KEYINPUT5), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n461), .B1(new_n464), .B2(new_n449), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n463), .A2(new_n441), .A3(new_n466), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT38), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n433), .A2(new_n476), .A3(new_n435), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n437), .A2(new_n468), .A3(new_n475), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n448), .A2(new_n455), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT39), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n480), .A3(new_n457), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n458), .A2(new_n459), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n480), .B1(new_n482), .B2(new_n449), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n464), .B2(new_n449), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n481), .A2(new_n484), .A3(KEYINPUT40), .A4(new_n441), .ZN(new_n485));
  INV_X1    g284(.A(new_n425), .ZN(new_n486));
  OR3_X1    g285(.A1(new_n434), .A2(KEYINPUT30), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n434), .A2(new_n486), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(KEYINPUT30), .A3(new_n426), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n472), .A2(new_n485), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n481), .A2(new_n441), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT40), .B1(new_n491), .B2(new_n484), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n412), .B1(new_n478), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n473), .B(new_n474), .C1(new_n467), .C2(KEYINPUT80), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n467), .A2(KEYINPUT80), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n468), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n489), .A2(new_n487), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n412), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n327), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n499), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT84), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n410), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n504), .A2(new_n398), .B1(new_n409), .B2(new_n410), .ZN(new_n505));
  AND4_X1   g304(.A1(KEYINPUT84), .A2(new_n409), .A3(new_n410), .A4(new_n398), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n319), .B(new_n321), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT35), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n322), .A2(new_n324), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n475), .A2(new_n468), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n499), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n512), .B1(new_n411), .B2(new_n408), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n501), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT86), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT86), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n520), .B(KEYINPUT13), .Z(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(G15gat), .B(G22gat), .Z(new_n523));
  INV_X1    g322(.A(G1gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(G1gat), .ZN(new_n528));
  INV_X1    g327(.A(G8gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT90), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n525), .A2(new_n528), .A3(KEYINPUT89), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n533), .B(G8gat), .C1(KEYINPUT89), .C2(new_n525), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT14), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G29gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT88), .B(G36gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT15), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n538), .B(KEYINPUT15), .C1(new_n539), .C2(new_n540), .ZN(new_n544));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n544), .A2(new_n545), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n535), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT91), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n548), .A3(KEYINPUT91), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n554));
  INV_X1    g353(.A(new_n535), .ZN(new_n555));
  INV_X1    g354(.A(new_n548), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n553), .A2(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n551), .A2(KEYINPUT92), .A3(new_n552), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n522), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n548), .A2(KEYINPUT17), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n546), .B2(new_n547), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n555), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n553), .A2(new_n520), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT18), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n559), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G197gat), .ZN(new_n570));
  XOR2_X1   g369(.A(KEYINPUT11), .B(G169gat), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n572), .B(new_n573), .Z(new_n574));
  NAND2_X1  g373(.A1(new_n564), .A2(new_n565), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n564), .A2(KEYINPUT93), .A3(new_n565), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n553), .A2(new_n554), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n555), .A2(new_n556), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n558), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n521), .ZN(new_n583));
  INV_X1    g382(.A(new_n567), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI22_X1  g384(.A1(new_n568), .A2(new_n574), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT8), .ZN(new_n587));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(KEYINPUT96), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n589), .B1(KEYINPUT96), .B2(new_n588), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT7), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT97), .B(G92gat), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n590), .B(new_n592), .C1(G85gat), .C2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G99gat), .B(G106gat), .Z(new_n595));
  OR2_X1    g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n560), .B2(new_n562), .ZN(new_n599));
  XOR2_X1   g398(.A(G190gat), .B(G218gat), .Z(new_n600));
  AND2_X1   g399(.A1(new_n596), .A2(new_n597), .ZN(new_n601));
  AND2_X1   g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n601), .A2(new_n548), .B1(KEYINPUT41), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n599), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT98), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n599), .A2(new_n603), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n606), .A2(new_n600), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(KEYINPUT99), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n608), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n605), .B(new_n607), .C1(KEYINPUT99), .C2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G57gat), .B(G64gat), .Z(new_n617));
  INV_X1    g416(.A(KEYINPUT9), .ZN(new_n618));
  INV_X1    g417(.A(G71gat), .ZN(new_n619));
  INV_X1    g418(.A(G78gat), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G71gat), .B(G78gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(new_n264), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n624), .B(KEYINPUT94), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n535), .B1(new_n630), .B2(KEYINPUT21), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n629), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G183gat), .B(G211gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT95), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n370), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n632), .B(new_n637), .Z(new_n638));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n639), .B1(new_n596), .B2(new_n597), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n596), .A2(new_n639), .A3(new_n597), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(new_n624), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n624), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n640), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT10), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n630), .A2(KEYINPUT10), .A3(new_n601), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(G230gat), .ZN(new_n649));
  OAI22_X1  g448(.A1(new_n646), .A2(new_n648), .B1(new_n649), .B2(new_n280), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n280), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n645), .A2(new_n643), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(G120gat), .B(G148gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT101), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n650), .A2(new_n652), .A3(new_n657), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n616), .A2(new_n638), .A3(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n517), .A2(new_n519), .A3(new_n586), .A4(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n498), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(new_n524), .ZN(G1324gat));
  XNOR2_X1  g464(.A(KEYINPUT16), .B(G8gat), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n663), .A2(new_n499), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n669));
  OR3_X1    g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n663), .ZN(new_n671));
  INV_X1    g470(.A(new_n499), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI22_X1  g472(.A1(G8gat), .A2(new_n673), .B1(new_n667), .B2(KEYINPUT42), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n668), .B1(new_n667), .B2(new_n669), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n670), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n670), .A2(new_n674), .A3(KEYINPUT104), .A4(new_n675), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(G1325gat));
  INV_X1    g479(.A(G15gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n671), .A2(new_n681), .A3(new_n509), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n325), .A2(new_n683), .A3(new_n326), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n325), .B2(new_n326), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n663), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n682), .B1(new_n681), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT106), .Z(G1326gat));
  NAND2_X1  g488(.A1(new_n408), .A2(new_n411), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n663), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(new_n616), .ZN(new_n694));
  INV_X1    g493(.A(new_n661), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n638), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n517), .A2(new_n519), .A3(new_n586), .A4(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(G29gat), .A3(new_n498), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n699), .A2(KEYINPUT45), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(KEYINPUT45), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n501), .A2(new_n515), .A3(new_n518), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n518), .B1(new_n501), .B2(new_n515), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n694), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n702), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n327), .A2(KEYINPUT105), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n412), .A2(new_n498), .A3(new_n499), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n433), .A2(new_n476), .A3(new_n435), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n476), .B1(new_n433), .B2(new_n435), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n710), .A2(new_n711), .A3(new_n427), .ZN(new_n712));
  INV_X1    g511(.A(new_n510), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n493), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n709), .B1(new_n714), .B2(new_n412), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n325), .A2(new_n683), .A3(new_n326), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n708), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n515), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT44), .B1(new_n718), .B2(new_n616), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n707), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n586), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n696), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n721), .A2(new_n498), .A3(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n700), .B(new_n701), .C1(new_n725), .C2(new_n539), .ZN(G1328gat));
  NAND2_X1  g525(.A1(new_n672), .A2(new_n540), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT46), .B1(new_n698), .B2(new_n727), .ZN(new_n728));
  OR3_X1    g527(.A1(new_n698), .A2(KEYINPUT46), .A3(new_n727), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n721), .A2(new_n499), .A3(new_n724), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n540), .ZN(G1329gat));
  INV_X1    g530(.A(G43gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n509), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n698), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT107), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n708), .A2(new_n716), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n736), .A3(new_n723), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G43gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n735), .A2(KEYINPUT47), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1330gat));
  OR3_X1    g542(.A1(new_n698), .A2(G50gat), .A3(new_n690), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n412), .A2(new_n713), .A3(new_n512), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n319), .A2(new_n321), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n746), .A2(new_n498), .A3(new_n690), .A4(new_n499), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n509), .A2(new_n745), .B1(new_n747), .B2(KEYINPUT35), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(new_n686), .B2(new_n715), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n704), .B1(new_n749), .B2(new_n694), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n517), .A2(new_n519), .A3(new_n705), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n750), .A2(new_n751), .A3(new_n412), .A4(new_n723), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G50gat), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n753), .ZN(new_n756));
  OAI211_X1 g555(.A(KEYINPUT48), .B(new_n744), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n752), .A2(G50gat), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n758), .A2(new_n744), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(KEYINPUT48), .B2(new_n759), .ZN(G1331gat));
  XNOR2_X1  g559(.A(new_n632), .B(new_n637), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n722), .A2(new_n694), .A3(new_n761), .A4(new_n661), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n749), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n498), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g565(.A(new_n499), .B(KEYINPUT109), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT49), .B(G64gat), .Z(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(G1333gat));
  NAND3_X1  g570(.A1(new_n763), .A2(G71gat), .A3(new_n736), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n763), .A2(new_n509), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n619), .B1(new_n773), .B2(KEYINPUT110), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n772), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g576(.A1(new_n763), .A2(new_n412), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g578(.A1(new_n586), .A2(new_n761), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT111), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(new_n661), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n720), .A2(new_n764), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G85gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n718), .A2(new_n616), .A3(new_n781), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n695), .A2(G85gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n764), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n784), .A2(new_n789), .ZN(G1336gat));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n786), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n785), .A2(new_n791), .A3(KEYINPUT51), .ZN(new_n794));
  INV_X1    g593(.A(new_n767), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n795), .A2(G92gat), .A3(new_n695), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT113), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n793), .A2(new_n799), .A3(new_n794), .A4(new_n796), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n720), .A2(new_n672), .A3(new_n782), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n593), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n798), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT52), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(new_n787), .B2(new_n796), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n720), .A2(new_n767), .A3(new_n782), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n593), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n804), .A2(new_n808), .ZN(G1337gat));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810));
  XNOR2_X1  g609(.A(KEYINPUT115), .B(G99gat), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n750), .A2(new_n751), .A3(new_n736), .A4(new_n782), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(KEYINPUT114), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(KEYINPUT114), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n695), .B1(new_n322), .B2(new_n324), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n812), .B1(new_n787), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n810), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n720), .A2(new_n821), .A3(new_n736), .A4(new_n782), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n813), .A2(KEYINPUT114), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n811), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(KEYINPUT116), .A3(new_n818), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n820), .A2(new_n825), .ZN(G1338gat));
  NOR3_X1   g625(.A1(new_n695), .A2(new_n690), .A3(G106gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n787), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n750), .A2(new_n751), .A3(new_n412), .A4(new_n782), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G106gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n793), .A2(new_n794), .A3(new_n827), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n831), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n833), .B1(new_n835), .B2(KEYINPUT53), .ZN(new_n836));
  AOI211_X1 g635(.A(KEYINPUT117), .B(new_n829), .C1(new_n834), .C2(new_n831), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n832), .B1(new_n836), .B2(new_n837), .ZN(G1339gat));
  INV_X1    g637(.A(KEYINPUT10), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n644), .A2(new_n640), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n601), .A2(new_n639), .A3(new_n624), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n651), .B1(new_n842), .B2(new_n647), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n657), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n842), .A2(new_n651), .A3(new_n647), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n650), .A2(KEYINPUT54), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n847), .A3(KEYINPUT55), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n660), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n845), .A2(new_n847), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI211_X1 g653(.A(KEYINPUT118), .B(KEYINPUT55), .C1(new_n845), .C2(new_n847), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n586), .B(new_n850), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n553), .A2(new_n563), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n582), .A2(new_n521), .B1(new_n520), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n572), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n859), .B(new_n661), .C1(new_n579), .C2(new_n585), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n616), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n559), .A2(new_n567), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(new_n574), .A3(new_n577), .A4(new_n578), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n863), .A2(new_n613), .A3(new_n615), .A4(new_n859), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n854), .A2(new_n855), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n864), .A2(new_n865), .A3(new_n849), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n638), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n662), .A2(new_n722), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n869), .A2(new_n498), .A3(new_n507), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(new_n795), .ZN(new_n871));
  AOI21_X1  g670(.A(G113gat), .B1(new_n871), .B2(new_n586), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n869), .A2(new_n412), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n509), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n767), .A2(new_n498), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n722), .A2(new_n270), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(G1340gat));
  INV_X1    g678(.A(new_n877), .ZN(new_n880));
  OAI21_X1  g679(.A(G120gat), .B1(new_n880), .B2(new_n695), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n695), .A2(new_n275), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n871), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1341gat));
  OAI21_X1  g683(.A(G127gat), .B1(new_n880), .B2(new_n638), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n871), .A2(new_n264), .A3(new_n761), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1342gat));
  AND4_X1   g686(.A1(new_n266), .A2(new_n870), .A3(new_n499), .A4(new_n616), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n888), .A2(KEYINPUT119), .A3(new_n889), .ZN(new_n893));
  INV_X1    g692(.A(new_n874), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n616), .A3(new_n875), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT56), .B1(new_n895), .B2(G134gat), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n892), .B(new_n893), .C1(new_n896), .C2(new_n888), .ZN(G1343gat));
  NOR2_X1   g696(.A1(new_n869), .A2(new_n498), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n736), .A2(new_n690), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n722), .A2(G141gat), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n898), .A2(new_n795), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT58), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT120), .B1(new_n902), .B2(KEYINPUT121), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n662), .A2(new_n722), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n854), .A2(new_n855), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n863), .A2(new_n859), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n906), .A2(new_n907), .A3(new_n616), .A4(new_n850), .ZN(new_n908));
  INV_X1    g707(.A(new_n860), .ZN(new_n909));
  INV_X1    g708(.A(new_n574), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n585), .B2(new_n566), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n849), .B1(new_n911), .B2(new_n863), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n852), .A2(new_n853), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n908), .B1(new_n914), .B2(new_n616), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n905), .B1(new_n915), .B2(new_n638), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT57), .B1(new_n916), .B2(new_n690), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n867), .A2(new_n868), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(new_n919), .A3(new_n412), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n736), .A2(new_n876), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n586), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n904), .B1(G141gat), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT121), .B1(new_n923), .B2(G141gat), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n898), .A2(new_n899), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n926), .A2(KEYINPUT120), .A3(new_n795), .A4(new_n900), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n924), .B1(new_n928), .B2(new_n902), .ZN(G1344gat));
  INV_X1    g728(.A(G148gat), .ZN(new_n930));
  AOI211_X1 g729(.A(KEYINPUT59), .B(new_n930), .C1(new_n922), .C2(new_n661), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n919), .B1(new_n916), .B2(new_n690), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n918), .A2(KEYINPUT57), .A3(new_n412), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n661), .A3(new_n921), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n932), .B1(new_n936), .B2(G148gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n926), .A2(new_n795), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n661), .A2(new_n930), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n931), .A2(new_n937), .B1(new_n938), .B2(new_n939), .ZN(G1345gat));
  INV_X1    g739(.A(new_n922), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n941), .A2(new_n370), .A3(new_n638), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n926), .A2(new_n761), .A3(new_n795), .ZN(new_n943));
  AOI21_X1  g742(.A(G155gat), .B1(new_n943), .B2(KEYINPUT122), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n945), .B1(new_n938), .B2(new_n638), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n942), .B1(new_n944), .B2(new_n946), .ZN(G1346gat));
  NOR2_X1   g746(.A1(new_n333), .A2(new_n334), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n926), .A2(new_n948), .A3(new_n499), .A4(new_n616), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n941), .A2(new_n694), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(new_n948), .ZN(G1347gat));
  NOR2_X1   g750(.A1(new_n869), .A2(new_n764), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n795), .A2(new_n507), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n954), .A2(new_n226), .A3(new_n722), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n764), .A2(new_n499), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n874), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(new_n586), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G169gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n957), .A2(new_n962), .ZN(G1348gat));
  OAI21_X1  g762(.A(new_n214), .B1(new_n954), .B2(new_n695), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n219), .A2(new_n221), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n873), .A2(new_n965), .A3(new_n817), .A4(new_n958), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n967), .B(new_n968), .ZN(G1349gat));
  NAND4_X1  g768(.A1(new_n873), .A2(new_n509), .A3(new_n761), .A4(new_n958), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(G183gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n761), .A2(new_n251), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n954), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT60), .ZN(G1350gat));
  AOI211_X1 g773(.A(KEYINPUT61), .B(new_n211), .C1(new_n960), .C2(new_n616), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT61), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n894), .A2(new_n616), .A3(new_n958), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n976), .B1(new_n977), .B2(G190gat), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n616), .A2(new_n211), .ZN(new_n979));
  OAI22_X1  g778(.A1(new_n975), .A2(new_n978), .B1(new_n954), .B2(new_n979), .ZN(G1351gat));
  NOR3_X1   g779(.A1(new_n736), .A2(new_n690), .A3(new_n795), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n981), .A2(KEYINPUT125), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(KEYINPUT125), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n952), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n984), .A2(new_n353), .A3(new_n586), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT126), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n736), .A2(new_n959), .ZN(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n989), .B1(new_n933), .B2(new_n934), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(new_n586), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT126), .B1(new_n991), .B2(G197gat), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n987), .B1(new_n992), .B2(new_n985), .ZN(G1352gat));
  NAND3_X1  g792(.A1(new_n984), .A2(new_n348), .A3(new_n661), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n995));
  INV_X1    g794(.A(new_n990), .ZN(new_n996));
  OAI21_X1  g795(.A(G204gat), .B1(new_n996), .B2(new_n695), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n995), .A2(new_n997), .A3(new_n998), .ZN(G1353gat));
  INV_X1    g798(.A(KEYINPUT63), .ZN(new_n1000));
  AOI211_X1 g799(.A(new_n919), .B(new_n690), .C1(new_n867), .C2(new_n868), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n586), .A2(new_n850), .A3(new_n913), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n616), .B1(new_n1002), .B2(new_n860), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n638), .B1(new_n1003), .B2(new_n866), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(new_n868), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT57), .B1(new_n1005), .B2(new_n412), .ZN(new_n1006));
  OAI211_X1 g805(.A(new_n761), .B(new_n988), .C1(new_n1001), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n1008));
  OAI21_X1  g807(.A(G211gat), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g808(.A(KEYINPUT127), .B1(new_n990), .B2(new_n761), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1000), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n990), .A2(KEYINPUT127), .A3(new_n761), .ZN(new_n1013));
  NAND4_X1  g812(.A1(new_n1012), .A2(new_n1013), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g814(.A(new_n346), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n984), .A2(new_n1016), .A3(new_n761), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1015), .A2(new_n1017), .ZN(G1354gat));
  OAI21_X1  g817(.A(G218gat), .B1(new_n996), .B2(new_n694), .ZN(new_n1019));
  INV_X1    g818(.A(G218gat), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n984), .A2(new_n1020), .A3(new_n616), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1019), .A2(new_n1021), .ZN(G1355gat));
endmodule


