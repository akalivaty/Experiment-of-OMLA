//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  XOR2_X1   g001(.A(G127gat), .B(G134gat), .Z(new_n203));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(KEYINPUT1), .B2(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G113gat), .B(G120gat), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  AND3_X1   g009(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(KEYINPUT23), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222));
  NOR3_X1   g021(.A1(new_n222), .A2(G169gat), .A3(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(KEYINPUT23), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n226), .B2(KEYINPUT64), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT25), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n229), .A2(KEYINPUT68), .A3(new_n230), .A4(new_n231), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT24), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n238), .B1(G183gat), .B2(G190gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT66), .ZN(new_n242));
  INV_X1    g041(.A(new_n211), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n238), .A2(G183gat), .A3(G190gat), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT24), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n236), .A2(new_n242), .A3(new_n243), .A4(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n219), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n251));
  NOR4_X1   g050(.A1(new_n226), .A2(new_n223), .A3(new_n250), .A4(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n228), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n225), .B(KEYINPUT26), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n219), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n212), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT28), .ZN(new_n257));
  NOR2_X1   g056(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT67), .B(G183gat), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(KEYINPUT27), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n257), .B1(new_n260), .B2(G190gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT27), .B(G183gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(KEYINPUT28), .A3(new_n230), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n256), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n210), .B1(new_n253), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G227gat), .ZN(new_n266));
  INV_X1    g065(.A(G233gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n205), .A2(new_n209), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n261), .A2(new_n263), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n255), .A2(new_n212), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n252), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n246), .B(KEYINPUT66), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n211), .B1(new_n234), .B2(new_n235), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n269), .B(new_n272), .C1(new_n276), .C2(new_n228), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n265), .A2(new_n268), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT33), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT69), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n282), .A3(new_n279), .ZN(new_n283));
  XNOR2_X1  g082(.A(G15gat), .B(G43gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT70), .ZN(new_n285));
  XNOR2_X1  g084(.A(G71gat), .B(G99gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n278), .B2(KEYINPUT32), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n281), .A2(new_n283), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n268), .B1(new_n265), .B2(new_n277), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT34), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI211_X1 g091(.A(KEYINPUT34), .B(new_n268), .C1(new_n265), .C2(new_n277), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n287), .B(KEYINPUT71), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n278), .B(KEYINPUT32), .C1(new_n279), .C2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n289), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n289), .A2(KEYINPUT72), .A3(new_n294), .A4(new_n296), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n294), .B1(new_n289), .B2(new_n296), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT90), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n302), .B1(new_n299), .B2(new_n300), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT90), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G197gat), .B(G204gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT22), .ZN(new_n311));
  INV_X1    g110(.A(G211gat), .ZN(new_n312));
  INV_X1    g111(.A(G218gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G211gat), .B(G218gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n310), .A3(new_n314), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n272), .B1(new_n276), .B2(new_n228), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n321), .A2(KEYINPUT74), .A3(G226gat), .A4(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(new_n253), .B2(new_n264), .ZN(new_n325));
  NAND2_X1  g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n253), .A2(new_n264), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(new_n326), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n320), .B(new_n322), .C1(new_n327), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT75), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n321), .A2(G226gat), .A3(G233gat), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n321), .A2(new_n324), .B1(G226gat), .B2(G233gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(new_n323), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n334), .A2(new_n335), .A3(new_n320), .A4(new_n322), .ZN(new_n336));
  INV_X1    g135(.A(new_n320), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n325), .A2(new_n326), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n332), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n331), .A2(new_n336), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT30), .ZN(new_n341));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n336), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n339), .A2(new_n337), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n345), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT30), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n340), .A2(new_n345), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n346), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT35), .ZN(new_n353));
  INV_X1    g152(.A(G148gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n356));
  INV_X1    g155(.A(G141gat), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n356), .B1(new_n357), .B2(G148gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(G148gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n361), .B1(new_n363), .B2(KEYINPUT2), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n361), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT76), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n361), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n361), .A2(KEYINPUT2), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G141gat), .B(G148gat), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n367), .B(new_n369), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n365), .A2(new_n373), .A3(KEYINPUT78), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(KEYINPUT3), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n357), .A2(G148gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n354), .A2(G141gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n382), .A2(new_n370), .B1(KEYINPUT76), .B2(new_n366), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n383), .A2(new_n369), .B1(new_n360), .B2(new_n364), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n210), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n210), .A2(new_n384), .A3(KEYINPUT4), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n374), .B2(new_n269), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n269), .A3(new_n377), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n210), .A2(new_n384), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT5), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT0), .ZN(new_n402));
  XNOR2_X1  g201(.A(G57gat), .B(G85gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n392), .B(new_n393), .C1(new_n398), .C2(new_n397), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n400), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n400), .A2(new_n406), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT88), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT88), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n400), .A2(new_n413), .A3(new_n406), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n404), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT6), .B1(new_n411), .B2(new_n404), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n410), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n324), .B1(new_n374), .B2(KEYINPUT3), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n337), .ZN(new_n420));
  NAND2_X1  g219(.A1(G228gat), .A2(G233gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n376), .A2(new_n377), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT3), .B1(new_n320), .B2(new_n324), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT83), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n421), .B1(new_n419), .B2(new_n337), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n428), .B(new_n429), .C1(new_n424), .C2(new_n425), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT82), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n431), .B1(new_n320), .B2(new_n324), .ZN(new_n432));
  AOI211_X1 g231(.A(KEYINPUT82), .B(KEYINPUT29), .C1(new_n318), .C2(new_n319), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n379), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n434), .A2(new_n374), .B1(new_n337), .B2(new_n419), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n421), .B(KEYINPUT81), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n427), .B(new_n430), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G22gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n320), .A2(new_n324), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT82), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n320), .A2(new_n431), .A3(new_n324), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT3), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n420), .B1(new_n442), .B2(new_n384), .ZN(new_n443));
  INV_X1    g242(.A(new_n436), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n428), .B1(new_n424), .B2(new_n425), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n443), .A2(new_n444), .B1(new_n445), .B2(KEYINPUT83), .ZN(new_n446));
  INV_X1    g245(.A(G22gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n447), .A3(new_n430), .ZN(new_n448));
  XOR2_X1   g247(.A(G78gat), .B(G106gat), .Z(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT31), .B(G50gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n448), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n447), .B1(new_n446), .B2(new_n430), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n451), .ZN(new_n456));
  INV_X1    g255(.A(new_n453), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n446), .A2(new_n447), .A3(new_n430), .A4(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n454), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n457), .B1(new_n437), .B2(G22gat), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n462), .A2(new_n448), .B1(new_n455), .B2(new_n451), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(KEYINPUT85), .A3(new_n458), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n352), .A2(new_n353), .A3(new_n418), .A4(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n202), .B1(new_n309), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n416), .A2(new_n407), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT80), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT80), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n416), .A2(new_n470), .A3(new_n407), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n471), .A3(new_n410), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n352), .A2(new_n472), .A3(new_n465), .A4(new_n306), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT35), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT85), .B1(new_n463), .B2(new_n458), .ZN(new_n475));
  AND4_X1   g274(.A1(KEYINPUT85), .A2(new_n454), .A3(new_n458), .A4(new_n456), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n418), .B(new_n353), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  AND4_X1   g276(.A1(new_n341), .A2(new_n347), .A3(new_n348), .A4(new_n345), .ZN(new_n478));
  INV_X1    g277(.A(new_n340), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n344), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n341), .B1(new_n340), .B2(new_n345), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n307), .B1(new_n301), .B2(new_n303), .ZN(new_n484));
  AOI211_X1 g283(.A(KEYINPUT90), .B(new_n302), .C1(new_n299), .C2(new_n300), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(KEYINPUT91), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n467), .A2(new_n474), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n400), .A2(new_n413), .A3(new_n406), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n413), .B1(new_n400), .B2(new_n406), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n405), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n409), .B1(new_n491), .B2(new_n416), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n349), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n334), .A2(new_n337), .A3(new_n322), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT37), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n339), .B2(new_n320), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n345), .A2(KEYINPUT38), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n495), .B2(new_n340), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT89), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n344), .B1(new_n479), .B2(KEYINPUT37), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n340), .A2(new_n495), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT38), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n500), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT89), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n505), .A2(new_n492), .A3(new_n506), .A4(new_n349), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n501), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n465), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT87), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n386), .A2(new_n390), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(new_n391), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n395), .A2(new_n391), .A3(new_n396), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT39), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n511), .A2(KEYINPUT39), .A3(new_n391), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n404), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n515), .A2(KEYINPUT86), .A3(new_n404), .A4(new_n517), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n510), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT40), .ZN(new_n523));
  OR2_X1    g322(.A1(KEYINPUT86), .A2(KEYINPUT87), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n518), .B2(new_n524), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n522), .A2(new_n415), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n509), .B1(new_n526), .B2(new_n482), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n508), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n306), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n465), .B1(new_n352), .B2(new_n472), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n488), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G183gat), .B(G211gat), .Z(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT16), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(G1gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541));
  MUX2_X1   g340(.A(G1gat), .B(new_n540), .S(new_n541), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G8gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT21), .ZN(new_n544));
  INV_X1    g343(.A(G64gat), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n545), .A2(G57gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT97), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n545), .A2(G57gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n549), .A2(KEYINPUT97), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n550), .B2(new_n546), .ZN(new_n551));
  NAND2_X1  g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  INV_X1    g351(.A(G71gat), .ZN(new_n553));
  INV_X1    g352(.A(G78gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT9), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT9), .B1(new_n546), .B2(new_n549), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(new_n552), .A3(new_n555), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n543), .B1(new_n544), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT99), .ZN(new_n563));
  XOR2_X1   g362(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n544), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT98), .ZN(new_n566));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  XNOR2_X1  g368(.A(G127gat), .B(G155gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n570), .B1(new_n568), .B2(new_n569), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n564), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n573), .ZN(new_n575));
  INV_X1    g374(.A(new_n564), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n571), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n563), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n574), .A2(new_n577), .A3(new_n563), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n538), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n580), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n582), .A2(new_n578), .A3(new_n537), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT102), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT7), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT101), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT101), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n594), .A3(KEYINPUT7), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n593), .B(new_n595), .C1(KEYINPUT7), .C2(new_n591), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G99gat), .B(G106gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT103), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n597), .A2(KEYINPUT103), .A3(new_n598), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n597), .A2(new_n598), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G43gat), .B(G50gat), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n606), .A2(KEYINPUT15), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(G29gat), .B2(G36gat), .ZN(new_n608));
  INV_X1    g407(.A(G29gat), .ZN(new_n609));
  INV_X1    g408(.A(G36gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT14), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n608), .B(new_n612), .C1(KEYINPUT15), .C2(new_n606), .ZN(new_n613));
  OAI22_X1  g412(.A1(new_n612), .A2(KEYINPUT92), .B1(new_n609), .B2(new_n610), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n612), .A2(KEYINPUT92), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n607), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n605), .A2(new_n617), .B1(KEYINPUT41), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n613), .A2(new_n616), .A3(KEYINPUT17), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n617), .A2(KEYINPUT93), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT93), .B1(new_n617), .B2(new_n621), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n620), .B(new_n604), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n619), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n630));
  XNOR2_X1  g429(.A(G134gat), .B(G162gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n627), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(KEYINPUT104), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT104), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n619), .A2(new_n624), .A3(new_n635), .A4(new_n628), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n636), .A3(new_n627), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n632), .B(KEYINPUT100), .Z(new_n639));
  AND3_X1   g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n638), .B1(new_n637), .B2(new_n639), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n633), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n585), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n543), .A2(KEYINPUT94), .ZN(new_n645));
  INV_X1    g444(.A(G8gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n542), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT94), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n620), .B(new_n650), .C1(new_n622), .C2(new_n623), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n617), .A2(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(G229gat), .A2(G233gat), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n651), .A2(KEYINPUT18), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n617), .B(new_n647), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n653), .B(KEYINPUT13), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n663));
  XNOR2_X1  g462(.A(G113gat), .B(G141gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT11), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(new_n216), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G197gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT12), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n659), .B(new_n662), .C1(new_n663), .C2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n663), .A3(new_n657), .ZN(new_n671));
  INV_X1    g470(.A(new_n662), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n671), .B(new_n668), .C1(new_n672), .C2(new_n658), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n558), .A2(KEYINPUT10), .A3(new_n560), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n604), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n561), .B1(new_n597), .B2(new_n598), .ZN(new_n678));
  AOI22_X1  g477(.A1(new_n604), .A2(new_n561), .B1(new_n603), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT10), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(G230gat), .A2(G233gat), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT106), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n604), .A2(new_n561), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n603), .A2(new_n678), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n686), .A2(new_n680), .A3(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n685), .B(new_n682), .C1(new_n688), .C2(new_n677), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n679), .A2(new_n682), .ZN(new_n690));
  XNOR2_X1  g489(.A(G120gat), .B(G148gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(G176gat), .B(G204gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n684), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n681), .A2(new_n683), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n696), .B2(new_n690), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n644), .A2(new_n675), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n536), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n472), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g503(.A1(new_n700), .A2(new_n352), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT42), .B1(new_n705), .B2(new_n646), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT16), .B(G8gat), .Z(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  MUX2_X1   g507(.A(KEYINPUT42), .B(new_n706), .S(new_n708), .Z(G1325gat));
  AOI21_X1  g508(.A(G15gat), .B1(new_n701), .B2(new_n486), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n532), .A2(G15gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT107), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n710), .B1(new_n701), .B2(new_n712), .ZN(G1326gat));
  NOR2_X1   g512(.A1(new_n700), .A2(new_n465), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT43), .B(G22gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n536), .A2(new_n717), .A3(new_n642), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT108), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n643), .B1(new_n488), .B2(new_n535), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n721), .A3(new_n717), .ZN(new_n722));
  INV_X1    g521(.A(new_n720), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n719), .A2(new_n722), .B1(KEYINPUT44), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n698), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n584), .A2(new_n674), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n728), .B2(new_n472), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n723), .A2(new_n726), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n609), .A3(new_n702), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT45), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(G1328gat));
  OAI21_X1  g532(.A(G36gat), .B1(new_n728), .B2(new_n352), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n730), .A2(new_n610), .A3(new_n482), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT46), .Z(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(G1329gat));
  AOI21_X1  g536(.A(G43gat), .B1(new_n730), .B2(new_n486), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n532), .A2(G43gat), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n727), .B2(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g540(.A(G50gat), .B1(new_n730), .B2(new_n509), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n509), .A2(G50gat), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n727), .B2(new_n743), .ZN(new_n744));
  XOR2_X1   g543(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1331gat));
  NOR3_X1   g545(.A1(new_n644), .A2(new_n674), .A3(new_n725), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n536), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n472), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(G57gat), .Z(G1332gat));
  OR2_X1    g549(.A1(new_n352), .A2(KEYINPUT110), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n352), .A2(KEYINPUT110), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI211_X1 g552(.A(new_n753), .B(new_n748), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1333gat));
  OAI21_X1  g555(.A(new_n553), .B1(new_n748), .B2(new_n309), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n532), .A2(G71gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n748), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g559(.A1(new_n748), .A2(new_n465), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(new_n554), .ZN(G1335gat));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n536), .A2(new_n764), .A3(new_n642), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n584), .A2(new_n675), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n720), .A2(new_n764), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n763), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n723), .A2(KEYINPUT112), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n766), .B1(new_n720), .B2(new_n764), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n772), .A3(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n774), .A2(new_n587), .A3(new_n702), .A4(new_n698), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n766), .A2(new_n725), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT111), .B1(new_n724), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n723), .A2(KEYINPUT44), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n720), .A2(new_n721), .A3(new_n717), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n721), .B1(new_n720), .B2(new_n717), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n783), .A3(new_n776), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n778), .A2(new_n702), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n775), .B1(new_n785), .B2(new_n587), .ZN(G1336gat));
  NAND3_X1  g585(.A1(new_n778), .A2(new_n784), .A3(new_n482), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT113), .B1(new_n771), .B2(new_n772), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(new_n763), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n753), .A2(G92gat), .A3(new_n725), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n787), .A2(G92gat), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n724), .A2(new_n777), .ZN(new_n793));
  INV_X1    g592(.A(new_n753), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n588), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n774), .ZN(new_n796));
  INV_X1    g595(.A(new_n790), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n792), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n791), .A2(new_n792), .B1(new_n795), .B2(new_n798), .ZN(G1337gat));
  NAND3_X1  g598(.A1(new_n778), .A2(new_n784), .A3(new_n532), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G99gat), .ZN(new_n801));
  OR3_X1    g600(.A1(new_n309), .A2(G99gat), .A3(new_n725), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n796), .B2(new_n802), .ZN(G1338gat));
  NAND3_X1  g602(.A1(new_n778), .A2(new_n784), .A3(new_n509), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n465), .A2(new_n725), .A3(G106gat), .ZN(new_n805));
  AOI22_X1  g604(.A1(new_n804), .A2(G106gat), .B1(new_n789), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT53), .B1(new_n774), .B2(new_n805), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n782), .A2(new_n509), .A3(new_n776), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G106gat), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n808), .A2(KEYINPUT114), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT114), .B1(new_n808), .B2(new_n810), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n806), .A2(new_n807), .B1(new_n811), .B2(new_n812), .ZN(G1339gat));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n681), .B2(new_n683), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n684), .A2(new_n815), .A3(new_n689), .ZN(new_n816));
  INV_X1    g615(.A(new_n693), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n696), .B2(new_n814), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n818), .A3(KEYINPUT55), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n816), .A2(new_n818), .A3(KEYINPUT115), .A4(KEYINPUT55), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n684), .A2(new_n689), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n821), .A2(new_n822), .B1(new_n823), .B2(new_n694), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n659), .A2(new_n669), .A3(new_n662), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n653), .B1(new_n651), .B2(new_n652), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n655), .A2(new_n656), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n667), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n816), .A2(new_n818), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n824), .A2(new_n642), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n725), .A2(new_n829), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n830), .A2(new_n831), .B1(new_n670), .B2(new_n673), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n824), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n833), .B1(new_n836), .B2(new_n642), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n584), .ZN(new_n838));
  NOR4_X1   g637(.A1(new_n584), .A2(new_n642), .A3(new_n674), .A4(new_n698), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n794), .A2(new_n472), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(new_n509), .A3(new_n304), .ZN(new_n844));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n674), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n843), .A2(new_n509), .A3(new_n309), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n674), .A2(G113gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(G1340gat));
  INV_X1    g647(.A(new_n846), .ZN(new_n849));
  OAI21_X1  g648(.A(G120gat), .B1(new_n849), .B2(new_n725), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n725), .A2(G120gat), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT116), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n844), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(G1341gat));
  AND3_X1   g653(.A1(new_n846), .A2(G127gat), .A3(new_n585), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n844), .A2(new_n585), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(G127gat), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(G1342gat));
  AOI21_X1  g659(.A(new_n839), .B1(new_n837), .B2(new_n584), .ZN(new_n861));
  NOR4_X1   g660(.A1(new_n861), .A2(new_n472), .A3(new_n482), .A4(new_n643), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n509), .A2(new_n304), .A3(G134gat), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n864), .B(new_n865), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT56), .ZN(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n849), .B2(new_n643), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1343gat));
  NOR2_X1   g668(.A1(new_n532), .A2(new_n465), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n674), .A2(new_n357), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n843), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n532), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n842), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n841), .A2(KEYINPUT57), .A3(new_n509), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n878), .B1(new_n861), .B2(new_n465), .ZN(new_n879));
  AOI211_X1 g678(.A(new_n675), .B(new_n876), .C1(new_n877), .C2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n874), .B1(new_n880), .B2(new_n357), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT58), .B1(new_n881), .B2(KEYINPUT119), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n876), .B1(new_n877), .B2(new_n879), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n357), .B1(new_n883), .B2(new_n674), .ZN(new_n884));
  NOR4_X1   g683(.A1(new_n884), .A2(KEYINPUT119), .A3(KEYINPUT120), .A4(new_n873), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  INV_X1    g685(.A(new_n876), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n841), .B2(new_n509), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n861), .A2(new_n878), .A3(new_n465), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n674), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n873), .B1(new_n890), .B2(G141gat), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n882), .B1(new_n885), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n892), .B(new_n874), .C1(new_n880), .C2(new_n357), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT120), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n897), .B1(new_n891), .B2(new_n892), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n891), .A2(new_n892), .A3(new_n886), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n894), .A2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n821), .A2(new_n822), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n695), .A3(new_n835), .ZN(new_n904));
  INV_X1    g703(.A(new_n834), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n642), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n824), .A2(new_n642), .A3(new_n832), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT122), .B(new_n833), .C1(new_n836), .C2(new_n642), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n585), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n509), .B1(new_n910), .B2(new_n839), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n889), .B1(new_n911), .B2(new_n878), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n887), .A2(new_n698), .ZN(new_n913));
  OAI21_X1  g712(.A(G148gat), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  XOR2_X1   g713(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT123), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n914), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n354), .A2(KEYINPUT59), .ZN(new_n920));
  INV_X1    g719(.A(new_n883), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n725), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n843), .A2(new_n871), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n354), .A3(new_n698), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1345gat));
  OAI21_X1  g725(.A(G155gat), .B1(new_n921), .B2(new_n584), .ZN(new_n927));
  INV_X1    g726(.A(G155gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n928), .A3(new_n585), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1346gat));
  OAI21_X1  g729(.A(G162gat), .B1(new_n921), .B2(new_n643), .ZN(new_n931));
  INV_X1    g730(.A(G162gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n862), .A2(new_n932), .A3(new_n870), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n702), .A2(new_n352), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n486), .A2(new_n935), .A3(new_n465), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n861), .A2(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(new_n216), .A3(new_n675), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n861), .A2(new_n702), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n753), .A2(new_n509), .A3(new_n304), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n674), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n938), .B1(new_n943), .B2(new_n216), .ZN(G1348gat));
  OAI21_X1  g743(.A(G176gat), .B1(new_n937), .B2(new_n725), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n698), .A2(new_n217), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n941), .B2(new_n946), .ZN(G1349gat));
  OAI21_X1  g746(.A(new_n259), .B1(new_n937), .B2(new_n584), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n585), .A2(new_n262), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n941), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g750(.A(G190gat), .B1(new_n937), .B2(new_n643), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT61), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n942), .A2(new_n230), .A3(new_n642), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n955), .B(new_n956), .ZN(G1351gat));
  NOR4_X1   g756(.A1(new_n861), .A2(new_n702), .A3(new_n753), .A4(new_n871), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n674), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n875), .A2(new_n935), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n960), .B(KEYINPUT125), .Z(new_n961));
  NOR2_X1   g760(.A1(new_n912), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n674), .A2(G197gat), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G1352gat));
  XOR2_X1   g763(.A(KEYINPUT126), .B(G204gat), .Z(new_n965));
  NAND3_X1  g764(.A1(new_n958), .A2(new_n698), .A3(new_n965), .ZN(new_n966));
  XOR2_X1   g765(.A(new_n966), .B(KEYINPUT62), .Z(new_n967));
  NOR3_X1   g766(.A1(new_n912), .A2(new_n725), .A3(new_n961), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n965), .B2(new_n968), .ZN(G1353gat));
  NAND3_X1  g768(.A1(new_n585), .A2(new_n875), .A3(new_n935), .ZN(new_n970));
  OAI21_X1  g769(.A(G211gat), .B1(new_n912), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g770(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  NAND3_X1  g771(.A1(new_n958), .A2(new_n312), .A3(new_n585), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1354gat));
  AOI21_X1  g773(.A(G218gat), .B1(new_n958), .B2(new_n642), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT127), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n643), .A2(new_n313), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n976), .B1(new_n962), .B2(new_n977), .ZN(G1355gat));
endmodule


