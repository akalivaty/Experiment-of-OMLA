//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n792, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1035, new_n1036;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  INV_X1    g006(.A(G127gat), .ZN(new_n208));
  INV_X1    g007(.A(G134gat), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n212));
  OAI21_X1  g011(.A(G127gat), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT69), .B1(new_n204), .B2(G120gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT70), .B1(new_n202), .B2(G113gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(new_n202), .A3(G113gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(new_n204), .A3(G120gat), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n214), .A2(new_n215), .A3(new_n217), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n207), .A2(KEYINPUT71), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT71), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n209), .ZN(new_n224));
  NAND2_X1  g023(.A1(G127gat), .A2(G134gat), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n221), .A2(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n210), .A2(new_n213), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(KEYINPUT74), .A2(G162gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(KEYINPUT74), .A2(G162gat), .ZN(new_n229));
  OAI21_X1  g028(.A(G155gat), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT2), .ZN(new_n231));
  INV_X1    g030(.A(G162gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G155gat), .ZN(new_n233));
  OR2_X1    g032(.A1(G141gat), .A2(G148gat), .ZN(new_n234));
  INV_X1    g033(.A(G155gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G162gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(G141gat), .A2(G148gat), .ZN(new_n237));
  AND4_X1   g036(.A1(new_n233), .A2(new_n234), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n233), .A2(new_n236), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT2), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n234), .A2(new_n240), .A3(new_n237), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n231), .A2(new_n238), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT4), .B1(new_n227), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n220), .A2(new_n226), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G120gat), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n213), .B(new_n224), .C1(KEYINPUT1), .C2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n241), .A2(new_n239), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT74), .B(G162gat), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n240), .B1(new_n250), .B2(G155gat), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n234), .A2(new_n233), .A3(new_n236), .A4(new_n237), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n249), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n244), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n227), .A2(new_n242), .A3(KEYINPUT77), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n243), .B1(new_n256), .B2(KEYINPUT4), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT5), .ZN(new_n258));
  NAND2_X1  g057(.A1(G225gat), .A2(G233gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n261), .B(new_n249), .C1(new_n251), .C2(new_n252), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT75), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n231), .A2(new_n238), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT75), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n261), .A4(new_n249), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n227), .B1(KEYINPUT3), .B2(new_n253), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n260), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n257), .A2(new_n258), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT4), .B1(new_n248), .B2(new_n253), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT76), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n227), .A2(new_n242), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT4), .B1(new_n254), .B2(new_n255), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n269), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n248), .A2(new_n253), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n254), .A2(new_n255), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n258), .B1(new_n281), .B2(new_n260), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n279), .A2(KEYINPUT78), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT78), .B1(new_n279), .B2(new_n282), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n271), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G1gat), .B(G29gat), .Z(new_n286));
  XNOR2_X1  g085(.A(G57gat), .B(G85gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n269), .A2(new_n258), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n291), .B1(new_n294), .B2(new_n257), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n283), .B2(new_n284), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT80), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT80), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n299), .B(new_n295), .C1(new_n283), .C2(new_n284), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n292), .A2(new_n297), .A3(new_n298), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT81), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n291), .A2(new_n285), .B1(new_n296), .B2(KEYINPUT80), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n300), .A2(new_n298), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT81), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n279), .A2(new_n282), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT78), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n279), .A2(KEYINPUT78), .A3(new_n282), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n290), .B1(new_n311), .B2(new_n271), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT6), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n302), .A2(new_n306), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G8gat), .B(G36gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(G64gat), .B(G92gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G226gat), .A2(G233gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G183gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT27), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G183gat), .ZN(new_n324));
  INV_X1    g123(.A(G190gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT66), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT28), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT28), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334));
  OR3_X1    g133(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT67), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT67), .B1(new_n333), .B2(new_n334), .ZN(new_n336));
  INV_X1    g135(.A(new_n334), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n335), .B(new_n336), .C1(KEYINPUT26), .C2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n330), .A2(new_n332), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT65), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(KEYINPUT23), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(KEYINPUT65), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n337), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n325), .ZN(new_n345));
  NAND2_X1  g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(KEYINPUT24), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT24), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n329), .A2(new_n348), .B1(G169gat), .B2(G176gat), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n344), .A2(KEYINPUT64), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n334), .A2(KEYINPUT23), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n344), .A2(new_n347), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n350), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n339), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n320), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G197gat), .B(G204gat), .ZN(new_n359));
  INV_X1    g158(.A(G211gat), .ZN(new_n360));
  INV_X1    g159(.A(G218gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(KEYINPUT22), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G211gat), .B(G218gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n344), .A2(new_n347), .A3(new_n349), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n366), .B(new_n351), .C1(KEYINPUT64), .C2(KEYINPUT25), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n319), .B1(new_n369), .B2(new_n339), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n358), .A2(new_n365), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n365), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n331), .A2(new_n328), .A3(new_n329), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n367), .A2(new_n368), .B1(new_n373), .B2(new_n338), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n319), .B1(new_n374), .B2(KEYINPUT29), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n320), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n318), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n365), .B1(new_n358), .B2(new_n370), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(new_n372), .A3(new_n376), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n317), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(KEYINPUT30), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n379), .A2(new_n380), .A3(new_n383), .A4(new_n317), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n372), .B1(new_n267), .B2(new_n357), .ZN(new_n387));
  OAI211_X1 g186(.A(G228gat), .B(G233gat), .C1(new_n387), .C2(KEYINPUT82), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n387), .ZN(new_n390));
  INV_X1    g189(.A(G22gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n261), .B1(new_n365), .B2(KEYINPUT29), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n253), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n391), .B1(new_n390), .B2(new_n393), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n389), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n390), .A2(new_n393), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G22gat), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(new_n394), .A3(new_n388), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G78gat), .B(G106gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT31), .B(G50gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n374), .A2(new_n248), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n356), .A2(new_n227), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n407), .A2(new_n408), .A3(G227gat), .A4(G233gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT32), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G15gat), .B(G43gat), .Z(new_n413));
  XNOR2_X1  g212(.A(G71gat), .B(G99gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n410), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n415), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n409), .B(KEYINPUT32), .C1(new_n411), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n407), .A2(new_n408), .B1(G227gat), .B2(G233gat), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT34), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(KEYINPUT72), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n424));
  OAI21_X1  g223(.A(new_n423), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n397), .A2(new_n404), .A3(new_n400), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(new_n416), .A3(new_n418), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n406), .A2(new_n427), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n314), .A2(new_n386), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT35), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n430), .A2(KEYINPUT35), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n301), .A2(new_n313), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(new_n386), .ZN(new_n437));
  AOI211_X1 g236(.A(KEYINPUT85), .B(new_n385), .C1(new_n301), .C2(new_n313), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n314), .A2(new_n386), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n406), .A2(new_n428), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT73), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT36), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n425), .A2(new_n416), .A3(new_n418), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n425), .B1(new_n416), .B2(new_n418), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n445), .B(new_n446), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n427), .A2(new_n443), .A3(new_n444), .A4(new_n429), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT40), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n267), .A2(new_n268), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n259), .B1(new_n257), .B2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n254), .A2(new_n255), .A3(new_n259), .A4(new_n280), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT39), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(KEYINPUT83), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n455), .B2(KEYINPUT39), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n454), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n257), .A2(new_n453), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT39), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n260), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n290), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n452), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n454), .ZN(new_n466));
  INV_X1    g265(.A(new_n457), .ZN(new_n467));
  INV_X1    g266(.A(new_n459), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n469), .A2(KEYINPUT40), .A3(new_n290), .A4(new_n463), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n292), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n441), .B1(new_n472), .B2(new_n385), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT37), .B1(new_n371), .B2(new_n377), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT37), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n379), .A2(new_n380), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n318), .A3(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT84), .B(KEYINPUT38), .Z(new_n478));
  OR2_X1    g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n381), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n477), .B2(new_n478), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n301), .A2(new_n313), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n451), .B1(new_n473), .B2(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n433), .A2(new_n439), .B1(new_n442), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT91), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n391), .A2(G15gat), .ZN(new_n486));
  INV_X1    g285(.A(G15gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(G22gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT16), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n486), .B(new_n488), .C1(new_n489), .C2(G1gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(G1gat), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G8gat), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT89), .B1(new_n491), .B2(G1gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI221_X1 g294(.A(new_n490), .B1(KEYINPUT89), .B2(G8gat), .C1(G1gat), .C2(new_n491), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT88), .ZN(new_n498));
  INV_X1    g297(.A(G29gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT14), .B(G29gat), .ZN(new_n502));
  INV_X1    g301(.A(G36gat), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g303(.A1(G43gat), .A2(G50gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(G43gat), .A2(G50gat), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT15), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G43gat), .ZN(new_n508));
  INV_X1    g307(.A(G50gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT15), .ZN(new_n511));
  NAND2_X1  g310(.A1(G43gat), .A2(G50gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n498), .B1(new_n504), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n507), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n504), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g316(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n518));
  NOR2_X1   g317(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n503), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n500), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n521), .A2(KEYINPUT88), .A3(new_n507), .A4(new_n513), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(new_n517), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n485), .B1(new_n497), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n522), .A2(new_n517), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n495), .A2(new_n496), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT91), .A4(new_n515), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n497), .A2(new_n523), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n497), .A2(KEYINPUT90), .A3(new_n523), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n534), .B(KEYINPUT13), .Z(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n523), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n515), .A2(KEYINPUT17), .A3(new_n522), .A4(new_n517), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n526), .A3(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n540), .A2(KEYINPUT18), .A3(new_n534), .A4(new_n529), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n529), .ZN(new_n543));
  INV_X1    g342(.A(new_n534), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n536), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT87), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G197gat), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT11), .B(G169gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n546), .A2(new_n547), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n484), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n314), .ZN(new_n561));
  XNOR2_X1  g360(.A(G120gat), .B(G148gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(KEYINPUT92), .A2(G57gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(KEYINPUT92), .A2(G57gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(G64gat), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G64gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(G57gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  INV_X1    g370(.A(G71gat), .ZN(new_n572));
  INV_X1    g371(.A(G78gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT9), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n568), .A2(new_n570), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n571), .ZN(new_n577));
  INV_X1    g376(.A(G57gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(G64gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n570), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n577), .B1(new_n580), .B2(KEYINPUT9), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT93), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n574), .A2(new_n571), .ZN(new_n583));
  AND2_X1   g382(.A1(KEYINPUT92), .A2(G57gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(KEYINPUT92), .A2(G57gat), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n584), .A2(new_n585), .A3(new_n569), .ZN(new_n586));
  INV_X1    g385(.A(new_n570), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n580), .A2(KEYINPUT9), .ZN(new_n589));
  INV_X1    g388(.A(new_n577), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT93), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n582), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT7), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  INV_X1    g396(.A(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(KEYINPUT8), .A2(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G99gat), .B(G106gat), .Z(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(new_n596), .A3(new_n600), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n594), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n603), .B(new_n605), .C1(new_n575), .C2(new_n581), .ZN(new_n608));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT10), .B1(new_n607), .B2(new_n608), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n606), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n618), .A2(new_n594), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n609), .B(KEYINPUT100), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n565), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT101), .ZN(new_n624));
  AND2_X1   g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625));
  OR3_X1    g424(.A1(new_n594), .A2(KEYINPUT21), .A3(new_n625), .ZN(new_n626));
  OAI211_X1 g425(.A(G231gat), .B(G233gat), .C1(new_n594), .C2(KEYINPUT21), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n626), .A2(new_n627), .A3(new_n208), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n208), .B1(new_n626), .B2(new_n627), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n497), .B1(new_n594), .B2(KEYINPUT21), .ZN(new_n630));
  OR3_X1    g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n630), .B1(new_n628), .B2(new_n629), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT94), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G155gat), .ZN(new_n636));
  XOR2_X1   g435(.A(G183gat), .B(G211gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n631), .A2(new_n632), .A3(new_n638), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(G232gat), .A2(G233gat), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n643), .A2(KEYINPUT41), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G190gat), .B(G218gat), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n647), .A2(KEYINPUT96), .B1(KEYINPUT41), .B2(new_n643), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n603), .A2(new_n605), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n523), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n538), .A2(new_n539), .A3(new_n606), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT95), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n650), .B1(new_n537), .B2(new_n523), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT95), .B1(new_n655), .B2(new_n539), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n651), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n647), .A2(KEYINPUT96), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n652), .A2(new_n653), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(KEYINPUT95), .A3(new_n539), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n658), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n663), .A3(new_n651), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n646), .B1(new_n659), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n659), .A2(new_n646), .A3(new_n664), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n615), .A2(new_n565), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n582), .A2(new_n593), .B1(new_n605), .B2(new_n603), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n575), .A2(new_n581), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n606), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n617), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n618), .A2(new_n594), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n610), .B1(new_n676), .B2(KEYINPUT97), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT97), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n674), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n670), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT97), .B1(new_n616), .B2(new_n619), .ZN(new_n681));
  AND4_X1   g480(.A1(new_n670), .A2(new_n681), .A3(new_n679), .A4(new_n609), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n669), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n624), .A2(new_n642), .A3(new_n668), .A4(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n560), .A2(new_n561), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g486(.A1(new_n292), .A2(new_n298), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n301), .B2(KEYINPUT81), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n385), .B1(new_n689), .B2(new_n306), .ZN(new_n690));
  INV_X1    g489(.A(new_n441), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n483), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT35), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n693), .B1(new_n690), .B2(new_n431), .ZN(new_n694));
  INV_X1    g493(.A(new_n434), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n303), .A2(new_n304), .B1(new_n312), .B2(KEYINPUT6), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT85), .B1(new_n696), .B2(new_n385), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n436), .A2(new_n435), .A3(new_n386), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n692), .B1(new_n694), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n558), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n684), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n493), .B1(new_n702), .B2(new_n385), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT16), .B(G8gat), .ZN(new_n704));
  NOR4_X1   g503(.A1(new_n701), .A2(new_n386), .A3(new_n684), .A4(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT42), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(KEYINPUT42), .B2(new_n705), .ZN(G1325gat));
  NOR2_X1   g506(.A1(new_n447), .A2(new_n448), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n702), .A2(new_n487), .A3(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n702), .A2(new_n451), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(new_n487), .ZN(G1326gat));
  NAND2_X1  g510(.A1(new_n702), .A2(new_n441), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT43), .B(G22gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n715));
  INV_X1    g514(.A(new_n642), .ZN(new_n716));
  INV_X1    g515(.A(new_n667), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n665), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n624), .A2(new_n683), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n560), .A2(new_n499), .A3(new_n561), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n715), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(KEYINPUT45), .A3(new_n723), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n642), .B(KEYINPUT103), .ZN(new_n729));
  INV_X1    g528(.A(new_n720), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(new_n558), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n484), .B2(new_n668), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n700), .A2(new_n718), .A3(new_n732), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n731), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n561), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G29gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n728), .A3(new_n741), .ZN(G1328gat));
  NAND4_X1  g541(.A1(new_n560), .A2(new_n503), .A3(new_n385), .A4(new_n721), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT46), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n743), .A2(KEYINPUT46), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n739), .A2(new_n385), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n503), .ZN(G1329gat));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n508), .B1(new_n739), .B2(new_n451), .ZN(new_n749));
  INV_X1    g548(.A(new_n708), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(G43gat), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n700), .A2(new_n558), .A3(new_n721), .A4(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n748), .B1(new_n749), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n731), .ZN(new_n756));
  AOI211_X1 g555(.A(new_n385), .B(new_n430), .C1(new_n689), .C2(new_n306), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n439), .B1(new_n757), .B2(new_n693), .ZN(new_n758));
  AOI211_X1 g557(.A(new_n668), .B(new_n733), .C1(new_n758), .C2(new_n692), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n735), .B1(new_n700), .B2(new_n718), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n451), .B(new_n756), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G43gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n752), .A2(KEYINPUT47), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT106), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n766), .B(new_n763), .C1(new_n761), .C2(G43gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n755), .B1(new_n765), .B2(new_n767), .ZN(G1330gat));
  NAND2_X1  g567(.A1(new_n441), .A2(new_n509), .ZN(new_n769));
  NOR4_X1   g568(.A1(new_n701), .A2(new_n720), .A3(new_n719), .A4(new_n769), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n441), .B(new_n756), .C1(new_n759), .C2(new_n760), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(G50gat), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g572(.A1(new_n642), .A2(new_n668), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n559), .A3(new_n720), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n484), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n561), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n777), .A2(KEYINPUT107), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n584), .A2(new_n585), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(KEYINPUT107), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(G1332gat));
  NAND2_X1  g582(.A1(new_n776), .A2(new_n385), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT49), .B(G64gat), .Z(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(G1333gat));
  AOI21_X1  g586(.A(new_n572), .B1(new_n776), .B2(new_n451), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n750), .A2(G71gat), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n776), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n441), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT108), .B(G78gat), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(G1335gat));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n642), .A2(new_n558), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n700), .A2(new_n718), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n668), .B1(new_n758), .B2(new_n692), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n801), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n796), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n314), .A2(G85gat), .A3(new_n730), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT110), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n720), .A2(new_n559), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n642), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n737), .B2(new_n738), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n561), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n806), .B1(new_n811), .B2(new_n598), .ZN(G1336gat));
  NOR3_X1   g611(.A1(new_n730), .A2(G92gat), .A3(new_n386), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n803), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n385), .B(new_n808), .C1(new_n759), .C2(new_n760), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT52), .B1(new_n815), .B2(G92gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n797), .A2(new_n818), .A3(KEYINPUT51), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT51), .B1(new_n797), .B2(new_n818), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n813), .B(KEYINPUT111), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n821), .A2(new_n822), .B1(G92gat), .B2(new_n815), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n817), .B1(new_n823), .B2(new_n824), .ZN(G1337gat));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n451), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n810), .A2(KEYINPUT113), .A3(new_n451), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(G99gat), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n750), .A2(G99gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n803), .A2(new_n720), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1338gat));
  NOR2_X1   g632(.A1(new_n691), .A2(G106gat), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n720), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n819), .A2(new_n820), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(G106gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n810), .B2(new_n441), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT53), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n803), .A2(new_n720), .A3(new_n834), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n441), .B(new_n808), .C1(new_n759), .C2(new_n760), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT53), .B1(new_n841), .B2(G106gat), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n843), .ZN(G1339gat));
  NAND2_X1  g643(.A1(new_n561), .A2(new_n386), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n536), .A2(new_n541), .A3(new_n545), .A4(new_n554), .ZN(new_n846));
  INV_X1    g645(.A(new_n535), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n528), .A2(new_n847), .A3(new_n531), .A4(new_n532), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n543), .A2(new_n544), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n552), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n717), .A2(new_n852), .A3(new_n665), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n620), .B2(new_n621), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n681), .A2(new_n679), .A3(new_n609), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT98), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n677), .A2(new_n670), .A3(new_n679), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n564), .B1(new_n622), .B2(new_n855), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n854), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n856), .B1(new_n680), .B2(new_n682), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(KEYINPUT55), .A3(new_n862), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n853), .A2(new_n864), .A3(new_n866), .A4(new_n683), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI211_X1 g668(.A(new_n565), .B(new_n615), .C1(new_n859), .C2(new_n860), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n861), .A2(new_n863), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(KEYINPUT55), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n872), .A2(KEYINPUT115), .A3(new_n864), .A4(new_n853), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n852), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n720), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n558), .A2(new_n864), .A3(new_n866), .A4(new_n683), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n718), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n729), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n730), .A2(new_n774), .A3(new_n880), .A4(new_n559), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT114), .B1(new_n684), .B2(new_n558), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI211_X1 g682(.A(new_n430), .B(new_n845), .C1(new_n879), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n558), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n720), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(G120gat), .ZN(G1341gat));
  NAND3_X1  g687(.A1(new_n884), .A2(new_n208), .A3(new_n642), .ZN(new_n889));
  INV_X1    g688(.A(new_n729), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n889), .B1(new_n891), .B2(new_n208), .ZN(G1342gat));
  NAND2_X1  g691(.A1(new_n884), .A2(new_n718), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n211), .A2(new_n212), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT116), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT116), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n899), .A3(new_n896), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n893), .B2(G134gat), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n898), .B(new_n900), .C1(new_n895), .C2(new_n901), .ZN(G1343gat));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n879), .A2(new_n883), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(KEYINPUT118), .A3(new_n561), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n451), .A2(new_n691), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT118), .B1(new_n904), .B2(new_n561), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n904), .A2(new_n561), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n912), .A2(KEYINPUT119), .A3(new_n905), .A4(new_n906), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n559), .A2(G141gat), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n909), .A2(new_n913), .A3(new_n386), .A4(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  INV_X1    g715(.A(new_n883), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n558), .A2(new_n866), .A3(new_n683), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT117), .B1(new_n861), .B2(new_n863), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n865), .A2(new_n920), .A3(new_n862), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n921), .A3(new_n854), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n918), .A2(new_n922), .B1(new_n720), .B2(new_n875), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n869), .B(new_n873), .C1(new_n923), .C2(new_n718), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n917), .B1(new_n924), .B2(new_n716), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT57), .B1(new_n925), .B2(new_n691), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n904), .A2(new_n927), .A3(new_n441), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n845), .A2(new_n451), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n926), .A2(new_n558), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(G141gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n916), .A3(new_n931), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n559), .A2(G141gat), .A3(new_n385), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n912), .A2(new_n905), .A3(new_n906), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT58), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n932), .A2(new_n936), .ZN(G1344gat));
  NAND3_X1  g736(.A1(new_n912), .A2(new_n905), .A3(new_n906), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n385), .B1(new_n938), .B2(new_n903), .ZN(new_n939));
  INV_X1    g738(.A(G148gat), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n720), .A4(new_n913), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n927), .B1(new_n904), .B2(new_n441), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n441), .A2(new_n927), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n918), .A2(new_n922), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n718), .B1(new_n945), .B2(new_n876), .ZN(new_n946));
  INV_X1    g745(.A(new_n867), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n716), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n685), .A2(new_n559), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n929), .A2(new_n720), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n943), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n940), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n904), .A2(new_n441), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT57), .ZN(new_n956));
  INV_X1    g755(.A(new_n950), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT120), .B1(new_n958), .B2(new_n951), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n942), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n961), .A2(new_n730), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n942), .A2(G148gat), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n941), .B1(new_n960), .B2(new_n964), .ZN(G1345gat));
  OAI21_X1  g764(.A(G155gat), .B1(new_n961), .B2(new_n729), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n939), .A2(new_n913), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n642), .A2(new_n235), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(G1346gat));
  OR2_X1    g768(.A1(new_n668), .A2(new_n250), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n926), .A2(new_n718), .A3(new_n928), .A4(new_n929), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT121), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n250), .B1(new_n971), .B2(new_n972), .ZN(new_n974));
  OAI22_X1  g773(.A1(new_n967), .A2(new_n970), .B1(new_n973), .B2(new_n974), .ZN(G1347gat));
  NAND2_X1  g774(.A1(new_n314), .A2(new_n385), .ZN(new_n976));
  AOI211_X1 g775(.A(new_n430), .B(new_n976), .C1(new_n879), .C2(new_n883), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(new_n558), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(G169gat), .ZN(G1348gat));
  INV_X1    g778(.A(G176gat), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n730), .B1(KEYINPUT122), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n980), .A2(KEYINPUT122), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n982), .B(new_n983), .ZN(G1349gat));
  NAND2_X1  g783(.A1(new_n977), .A2(new_n890), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n977), .A2(KEYINPUT124), .A3(new_n890), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n987), .A2(G183gat), .A3(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT123), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n642), .A2(new_n322), .A3(new_n324), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n977), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n991), .B1(new_n977), .B2(new_n992), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n990), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g795(.A(KEYINPUT60), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(new_n995), .ZN(new_n998));
  AOI21_X1  g797(.A(KEYINPUT125), .B1(new_n998), .B2(new_n993), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT60), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n987), .A2(G183gat), .A3(new_n988), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n997), .A2(new_n1002), .ZN(G1350gat));
  NOR2_X1   g802(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1004), .B1(new_n977), .B2(new_n718), .ZN(new_n1005));
  NAND2_X1  g804(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n1006));
  XOR2_X1   g805(.A(new_n1005), .B(new_n1006), .Z(G1351gat));
  INV_X1    g806(.A(G197gat), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n976), .A2(new_n451), .ZN(new_n1009));
  NAND4_X1  g808(.A1(new_n956), .A2(new_n957), .A3(new_n558), .A4(new_n1009), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT126), .ZN(new_n1011));
  AOI21_X1  g810(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1012), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n904), .A2(new_n441), .A3(new_n1009), .ZN(new_n1014));
  INV_X1    g813(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1015), .A2(new_n1008), .A3(new_n558), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1013), .A2(new_n1016), .ZN(G1352gat));
  NOR3_X1   g816(.A1(new_n1014), .A2(G204gat), .A3(new_n730), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(KEYINPUT62), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n956), .A2(new_n957), .A3(new_n1009), .ZN(new_n1020));
  OAI21_X1  g819(.A(G204gat), .B1(new_n1020), .B2(new_n730), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1019), .A2(new_n1021), .ZN(G1353gat));
  INV_X1    g821(.A(KEYINPUT63), .ZN(new_n1023));
  INV_X1    g822(.A(new_n1009), .ZN(new_n1024));
  NOR4_X1   g823(.A1(new_n943), .A2(new_n950), .A3(new_n716), .A4(new_n1024), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1023), .B1(new_n1025), .B2(new_n360), .ZN(new_n1026));
  NAND4_X1  g825(.A1(new_n956), .A2(new_n957), .A3(new_n642), .A4(new_n1009), .ZN(new_n1027));
  NAND3_X1  g826(.A1(new_n1027), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n1026), .A2(KEYINPUT127), .A3(new_n1028), .ZN(new_n1029));
  NOR3_X1   g828(.A1(new_n1014), .A2(G211gat), .A3(new_n716), .ZN(new_n1030));
  AOI21_X1  g829(.A(KEYINPUT63), .B1(new_n1027), .B2(G211gat), .ZN(new_n1031));
  INV_X1    g830(.A(KEYINPUT127), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g832(.A1(new_n1029), .A2(new_n1033), .ZN(G1354gat));
  OAI21_X1  g833(.A(G218gat), .B1(new_n1020), .B2(new_n668), .ZN(new_n1035));
  NAND3_X1  g834(.A1(new_n1015), .A2(new_n361), .A3(new_n718), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n1035), .A2(new_n1036), .ZN(G1355gat));
endmodule


