//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n217), .A2(KEYINPUT66), .A3(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n220), .B1(new_n201), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(KEYINPUT64), .B(G238), .Z(new_n223));
  AOI21_X1  g0023(.A(new_n222), .B1(G68), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(KEYINPUT66), .B1(new_n217), .B2(new_n218), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n212), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n211), .B(new_n215), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT67), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(G20), .ZN(new_n248));
  INV_X1    g0048(.A(G68), .ZN(new_n249));
  AOI22_X1  g0049(.A1(new_n248), .A2(G77), .B1(G20), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n250), .B1(new_n201), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n208), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT11), .ZN(new_n257));
  OR2_X1    g0057(.A1(KEYINPUT69), .A2(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT69), .A2(G1), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n258), .A2(G13), .A3(G20), .A4(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G68), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n261), .B(KEYINPUT12), .Z(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT69), .A2(G1), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT69), .A2(G1), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n263), .A2(new_n264), .A3(new_n209), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n255), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G68), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n257), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT14), .ZN(new_n269));
  AND2_X1   g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n208), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G97), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n272), .B1(new_n275), .B2(new_n221), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(G232), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(new_n274), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n271), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(G274), .B1(new_n270), .B2(new_n208), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G41), .A2(G45), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n280), .A2(G1), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n281), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n263), .A2(new_n264), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n271), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n282), .B1(G238), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT13), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n279), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(new_n279), .B2(new_n286), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n269), .B(G169), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n289), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n279), .A2(new_n286), .A3(new_n287), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n290), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n269), .B1(new_n293), .B2(G169), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n268), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n293), .A2(G200), .ZN(new_n298));
  INV_X1    g0098(.A(new_n268), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n298), .B(new_n299), .C1(new_n300), .C2(new_n293), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n273), .A2(G223), .A3(new_n274), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G87), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n273), .A2(G1698), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n303), .B(new_n304), .C1(new_n305), .C2(new_n221), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n271), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n282), .B1(G232), .B2(new_n285), .ZN(new_n308));
  AOI21_X1  g0108(.A(G169), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n307), .A2(new_n308), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n309), .B1(new_n294), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT7), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n273), .A2(new_n312), .A3(G20), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT7), .B1(new_n317), .B2(new_n209), .ZN(new_n318));
  OAI21_X1  g0118(.A(G68), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n251), .A2(G159), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n202), .A2(new_n249), .ZN(new_n321));
  NOR2_X1   g0121(.A1(G58), .A2(G68), .ZN(new_n322));
  OAI21_X1  g0122(.A(G20), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n319), .A2(KEYINPUT16), .A3(new_n320), .A4(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT16), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n312), .B1(new_n273), .B2(G20), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n317), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n249), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n323), .A2(new_n320), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n324), .A2(new_n330), .A3(new_n255), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT8), .B(G58), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(new_n260), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n333), .B2(new_n266), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n311), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT18), .ZN(new_n338));
  INV_X1    g0138(.A(new_n336), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n307), .A2(new_n308), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G200), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n300), .A2(KEYINPUT74), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n300), .A2(KEYINPUT74), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n307), .A2(new_n308), .A3(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n339), .A2(new_n347), .A3(KEYINPUT17), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT18), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n311), .A2(new_n336), .A3(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n331), .A2(new_n341), .A3(new_n335), .A4(new_n346), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT17), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n338), .A2(new_n348), .A3(new_n350), .A4(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  INV_X1    g0156(.A(new_n271), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n223), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G107), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n277), .A2(G1698), .B1(new_n362), .B2(new_n273), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n357), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n282), .B1(G244), .B2(new_n285), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n356), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n358), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n363), .B1(new_n370), .B2(new_n223), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n294), .B(new_n366), .C1(new_n371), .C2(new_n357), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n266), .A2(G77), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G77), .B2(new_n260), .ZN(new_n374));
  INV_X1    g0174(.A(new_n255), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n333), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n376));
  XOR2_X1   g0176(.A(KEYINPUT15), .B(G87), .Z(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n248), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n375), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n368), .A2(new_n372), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(G200), .B1(new_n365), .B2(new_n367), .ZN(new_n383));
  OAI211_X1 g0183(.A(G190), .B(new_n366), .C1(new_n371), .C2(new_n357), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n384), .A3(new_n380), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n302), .A2(new_n355), .A3(new_n382), .A4(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(G223), .B1(new_n359), .B2(new_n360), .ZN(new_n387));
  INV_X1    g0187(.A(G222), .ZN(new_n388));
  INV_X1    g0188(.A(G77), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n275), .A2(new_n388), .B1(new_n389), .B2(new_n273), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n357), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n282), .B1(G226), .B2(new_n285), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(G200), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT73), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT73), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n397), .B(G200), .C1(new_n392), .C2(new_n394), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n392), .A2(new_n394), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G190), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n260), .A2(new_n201), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n266), .B2(new_n201), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT71), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n403), .B(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n333), .A2(new_n248), .B1(G150), .B2(new_n251), .ZN(new_n406));
  OAI21_X1  g0206(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n255), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n405), .A2(KEYINPUT9), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT9), .B1(new_n405), .B2(new_n409), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n401), .B(new_n412), .C1(KEYINPUT72), .C2(KEYINPUT10), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n395), .A2(KEYINPUT73), .B1(new_n399), .B2(G190), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(new_n414), .A3(new_n398), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(KEYINPUT72), .A3(new_n398), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT10), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n399), .A2(new_n294), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n405), .A2(new_n409), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n419), .B(new_n420), .C1(G169), .C2(new_n399), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n413), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n386), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT85), .ZN(new_n425));
  INV_X1    g0225(.A(G116), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n254), .A2(new_n208), .B1(G20), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G283), .ZN(new_n428));
  INV_X1    g0228(.A(G97), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n428), .B(new_n209), .C1(G33), .C2(new_n429), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n427), .A2(KEYINPUT20), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT20), .B1(new_n427), .B2(new_n430), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n258), .A2(G33), .A3(new_n259), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n260), .A2(new_n375), .A3(new_n434), .A4(G116), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n265), .A2(G13), .A3(new_n426), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n425), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n427), .A2(new_n430), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT20), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n427), .A2(KEYINPUT20), .A3(new_n430), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n443), .A2(KEYINPUT85), .A3(new_n436), .A4(new_n435), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n438), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT5), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT76), .B1(new_n446), .B2(G41), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT76), .ZN(new_n448));
  INV_X1    g0248(.A(G41), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(new_n280), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n446), .A2(G41), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n258), .A2(new_n453), .A3(G45), .A4(new_n259), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT75), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT75), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n284), .A2(new_n456), .A3(G45), .A4(new_n453), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n357), .B(G270), .C1(new_n454), .C2(new_n451), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n315), .A2(G33), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n462));
  OAI21_X1  g0262(.A(G303), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n314), .A2(new_n316), .A3(G264), .A4(G1698), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n314), .A2(new_n316), .A3(G257), .A4(new_n274), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT84), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT84), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n463), .A2(new_n464), .A3(new_n465), .A4(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n271), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n460), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n445), .A2(KEYINPUT21), .A3(new_n471), .A4(G169), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n458), .A2(new_n459), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n357), .B1(new_n466), .B2(KEYINPUT84), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n445), .A2(new_n475), .A3(G179), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n314), .A2(new_n316), .A3(new_n209), .A4(G87), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT22), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT22), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n273), .A2(new_n480), .A3(new_n209), .A4(G87), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT23), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n209), .B2(G107), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n362), .A2(KEYINPUT23), .A3(G20), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n248), .A2(G116), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT24), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n375), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n488), .B1(new_n479), .B2(new_n481), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT24), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT25), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n265), .A2(new_n495), .A3(G13), .A4(new_n362), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n260), .A2(new_n375), .A3(new_n434), .A4(G107), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT25), .B1(new_n260), .B2(G107), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT86), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(KEYINPUT86), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n492), .A2(new_n494), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n314), .A2(new_n316), .A3(G257), .A4(G1698), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n314), .A2(new_n316), .A3(G250), .A4(new_n274), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G294), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n271), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n357), .B(G264), .C1(new_n454), .C2(new_n451), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n458), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n356), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n458), .A2(new_n508), .A3(new_n294), .A4(new_n509), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n356), .B1(new_n438), .B2(new_n444), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT21), .B1(new_n515), .B2(new_n471), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n477), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n460), .A2(new_n470), .A3(new_n345), .ZN(new_n518));
  INV_X1    g0318(.A(G200), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n460), .B2(new_n470), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n518), .A2(new_n520), .A3(new_n445), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n501), .A2(new_n502), .ZN(new_n522));
  INV_X1    g0322(.A(new_n494), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n255), .B1(new_n493), .B2(KEYINPUT24), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n510), .A2(G200), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n458), .A2(new_n508), .A3(G190), .A4(new_n509), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT87), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT87), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n503), .A2(new_n530), .A3(new_n527), .A4(new_n526), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n521), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n517), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n362), .A2(KEYINPUT6), .A3(G97), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n429), .A2(new_n362), .ZN(new_n535));
  NOR2_X1   g0335(.A1(G97), .A2(G107), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n534), .B1(new_n537), .B2(KEYINPUT6), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(G20), .B1(G77), .B2(new_n251), .ZN(new_n539));
  OAI21_X1  g0339(.A(G107), .B1(new_n313), .B2(new_n318), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n375), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n260), .A2(new_n375), .A3(new_n434), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G97), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(G97), .B2(new_n260), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n314), .A2(new_n316), .A3(G244), .A4(new_n274), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT4), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n273), .A2(KEYINPUT4), .A3(G244), .A4(new_n274), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n273), .A2(G250), .A3(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n428), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n271), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n357), .B(G257), .C1(new_n454), .C2(new_n451), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n458), .A2(KEYINPUT77), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT77), .B1(new_n458), .B2(new_n555), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n294), .B(new_n554), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(new_n458), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n356), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n547), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n458), .A2(new_n555), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT77), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n458), .A2(KEYINPUT77), .A3(new_n555), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n519), .B1(new_n566), .B2(new_n554), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n458), .A2(new_n555), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(G190), .A3(new_n554), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n546), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT78), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n554), .B1(new_n556), .B2(new_n557), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G200), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT78), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n573), .A2(new_n574), .A3(new_n546), .A4(new_n569), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n561), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n260), .A2(new_n377), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n314), .A2(new_n316), .A3(new_n209), .A4(G68), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT79), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n273), .A2(KEYINPUT79), .A3(new_n209), .A4(G68), .ZN(new_n581));
  NOR3_X1   g0381(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n582));
  AOI21_X1  g0382(.A(G20), .B1(G33), .B2(G97), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT19), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n248), .A2(new_n585), .A3(G97), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n580), .A2(new_n581), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT80), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n255), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n580), .A2(new_n581), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n586), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n590), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n577), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT81), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(KEYINPUT81), .B(new_n577), .C1(new_n589), .C2(new_n592), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n595), .A2(new_n596), .B1(G87), .B2(new_n543), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n314), .A2(new_n316), .A3(G244), .A4(G1698), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n314), .A2(new_n316), .A3(G238), .A4(new_n274), .ZN(new_n599));
  NAND2_X1  g0399(.A1(G33), .A2(G116), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n258), .A2(G45), .A3(new_n259), .ZN(new_n602));
  INV_X1    g0402(.A(G250), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n271), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(G274), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n284), .A2(G45), .A3(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n271), .A2(new_n601), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n519), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(G190), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n609), .A2(KEYINPUT83), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(KEYINPUT83), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n597), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n601), .A2(new_n271), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n604), .A2(new_n606), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G169), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n607), .A2(G179), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n595), .A2(new_n596), .B1(new_n377), .B2(new_n543), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(KEYINPUT82), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n590), .A2(new_n591), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT80), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n587), .A2(new_n588), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n255), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT81), .B1(new_n625), .B2(new_n577), .ZN(new_n626));
  INV_X1    g0426(.A(new_n596), .ZN(new_n627));
  INV_X1    g0427(.A(new_n377), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n626), .A2(new_n627), .B1(new_n628), .B2(new_n542), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT82), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n576), .B(new_n613), .C1(new_n621), .C2(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n424), .A2(new_n533), .A3(new_n632), .ZN(G372));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n595), .A2(new_n596), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n543), .A2(G87), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n635), .A2(new_n612), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n619), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n629), .B2(new_n630), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n620), .A2(KEYINPUT82), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n634), .B1(new_n641), .B2(new_n561), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n629), .A2(new_n619), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n608), .B1(G190), .B2(new_n607), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n597), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n643), .A2(new_n645), .A3(new_n634), .A4(new_n561), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n571), .A2(new_n575), .ZN(new_n647));
  INV_X1    g0447(.A(new_n561), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n647), .A2(new_n643), .A3(new_n648), .A4(new_n645), .ZN(new_n649));
  INV_X1    g0449(.A(new_n514), .ZN(new_n650));
  INV_X1    g0450(.A(new_n516), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(new_n476), .A4(new_n472), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n529), .A2(new_n531), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n643), .B(new_n646), .C1(new_n649), .C2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n423), .B1(new_n642), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n349), .B1(new_n311), .B2(new_n336), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n311), .A2(new_n336), .A3(new_n349), .ZN(new_n658));
  INV_X1    g0458(.A(new_n382), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n301), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n297), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n351), .B(KEYINPUT17), .ZN(new_n662));
  AOI211_X1 g0462(.A(new_n657), .B(new_n658), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n413), .A2(new_n418), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n421), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n656), .A2(new_n666), .ZN(G369));
  NOR2_X1   g0467(.A1(new_n477), .A2(new_n516), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n209), .A2(G13), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n284), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G343), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n445), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n668), .B(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n521), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G330), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n503), .A2(new_n675), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT88), .ZN(new_n684));
  INV_X1    g0484(.A(new_n653), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n650), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n650), .A2(new_n676), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n682), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n668), .A2(new_n676), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n687), .B1(new_n686), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n213), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n582), .A2(new_n426), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n697), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n206), .B2(new_n697), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n703), .B(new_n675), .C1(new_n642), .C2(new_n655), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n639), .A2(new_n640), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n634), .A3(new_n561), .A4(new_n613), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n643), .A2(new_n645), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT26), .B1(new_n708), .B2(new_n648), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n629), .A2(new_n619), .B1(new_n597), .B2(new_n644), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n576), .A3(new_n652), .A4(new_n653), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n707), .A2(new_n709), .A3(new_n643), .A4(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n703), .B1(new_n712), .B2(new_n675), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n517), .A2(new_n532), .A3(new_n675), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n641), .A2(new_n715), .A3(new_n576), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n510), .A2(new_n294), .A3(new_n616), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n572), .A2(new_n717), .A3(new_n471), .ZN(new_n718));
  XNOR2_X1  g0518(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n719));
  INV_X1    g0519(.A(new_n454), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n447), .A2(new_n450), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n271), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n722), .A2(G264), .B1(new_n271), .B2(new_n507), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n568), .A2(new_n723), .A3(new_n554), .A4(new_n607), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n460), .A2(new_n470), .A3(G179), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n719), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n718), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT90), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n607), .A2(new_n509), .A3(new_n508), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n559), .A2(new_n730), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n460), .A2(new_n470), .A3(G179), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(KEYINPUT30), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n718), .A2(new_n726), .A3(KEYINPUT90), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n729), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n675), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n733), .A2(new_n718), .A3(new_n726), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n676), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n735), .A2(new_n737), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n681), .B1(new_n716), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n714), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n702), .B1(new_n744), .B2(G1), .ZN(G364));
  INV_X1    g0545(.A(G1), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n669), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n696), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n682), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(G330), .B1(new_n678), .B2(new_n679), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n680), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n695), .A2(new_n317), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G355), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G116), .B2(new_n213), .ZN(new_n759));
  INV_X1    g0559(.A(G45), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n242), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n695), .A2(new_n273), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n760), .B2(new_n207), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n759), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n208), .B1(G20), .B2(new_n356), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n755), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n749), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n766), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G179), .A2(G200), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n209), .B1(new_n771), .B2(G190), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n429), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n209), .A2(new_n294), .A3(new_n519), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G190), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n773), .B1(new_n776), .B2(G68), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n209), .A2(new_n294), .A3(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n345), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n777), .B1(new_n202), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n209), .A2(G190), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n771), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT32), .Z(new_n785));
  NOR2_X1   g0585(.A1(new_n775), .A2(new_n344), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n778), .A2(new_n300), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n787), .A2(new_n201), .B1(new_n389), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n519), .A2(G179), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n781), .ZN(new_n791));
  INV_X1    g0591(.A(G87), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n790), .A2(G20), .A3(G190), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n273), .B1(new_n791), .B2(new_n362), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  OR4_X1    g0594(.A1(new_n780), .A2(new_n785), .A3(new_n789), .A4(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n772), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n786), .A2(G326), .B1(G294), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT91), .ZN(new_n798));
  INV_X1    g0598(.A(new_n779), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G322), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT33), .B(G317), .ZN(new_n801));
  INV_X1    g0601(.A(new_n788), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n776), .A2(new_n801), .B1(new_n802), .B2(G311), .ZN(new_n803));
  INV_X1    g0603(.A(new_n782), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n273), .B1(new_n804), .B2(G329), .ZN(new_n805));
  INV_X1    g0605(.A(G283), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n806), .B2(new_n791), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n793), .B(KEYINPUT92), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(G303), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n798), .A2(new_n800), .A3(new_n803), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n770), .B1(new_n795), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n769), .A2(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n750), .A2(new_n752), .B1(new_n756), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  OAI21_X1  g0614(.A(new_n675), .B1(new_n642), .B2(new_n655), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n676), .A2(new_n381), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n382), .A2(new_n385), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT96), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n659), .A2(new_n676), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n382), .A2(new_n385), .A3(KEYINPUT96), .A4(new_n816), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n815), .A2(new_n823), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n824), .A2(KEYINPUT97), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(KEYINPUT97), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n819), .A2(new_n821), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n675), .B(new_n827), .C1(new_n642), .C2(new_n655), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n749), .B1(new_n829), .B2(new_n742), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n742), .B2(new_n829), .ZN(new_n831));
  INV_X1    g0631(.A(new_n749), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n766), .A2(new_n753), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n389), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n273), .B1(new_n808), .B2(G107), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT93), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n791), .A2(new_n792), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n773), .B(new_n837), .C1(G311), .C2(new_n804), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n776), .A2(G283), .B1(new_n802), .B2(G116), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n799), .A2(G294), .B1(G303), .B2(new_n786), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n836), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n786), .A2(G137), .B1(new_n802), .B2(G159), .ZN(new_n842));
  INV_X1    g0642(.A(G143), .ZN(new_n843));
  INV_X1    g0643(.A(G150), .ZN(new_n844));
  INV_X1    g0644(.A(new_n776), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n842), .B1(new_n843), .B2(new_n779), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT34), .Z(new_n847));
  NOR2_X1   g0647(.A1(new_n791), .A2(new_n249), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(new_n808), .B2(G50), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n849), .A2(KEYINPUT94), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(KEYINPUT94), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n273), .B1(new_n772), .B2(new_n202), .C1(new_n852), .C2(new_n782), .ZN(new_n853));
  OR3_X1    g0653(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n841), .B1(new_n847), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT95), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n766), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n855), .A2(KEYINPUT95), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n834), .B1(new_n822), .B2(new_n754), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n831), .A2(new_n859), .ZN(G384));
  OAI21_X1  g0660(.A(new_n423), .B1(new_n705), .B2(new_n713), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n666), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT99), .Z(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n336), .A2(new_n674), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n658), .A2(new_n657), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n865), .B1(new_n866), .B2(new_n662), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n337), .A2(new_n865), .A3(new_n351), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n337), .A2(new_n865), .A3(KEYINPUT37), .A4(new_n351), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n864), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n865), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n354), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n875), .A2(KEYINPUT38), .A3(new_n871), .A4(new_n870), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n297), .A2(new_n676), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n873), .A2(new_n876), .A3(KEYINPUT39), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n866), .A2(new_n674), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n659), .A2(new_n675), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n828), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT98), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n268), .A2(new_n889), .A3(new_n676), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n268), .B2(new_n676), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n297), .A2(new_n301), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n892), .B1(new_n297), .B2(new_n301), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n888), .A2(new_n895), .A3(new_n877), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n886), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n863), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n822), .B1(new_n893), .B2(new_n894), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n873), .B2(new_n876), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT100), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n739), .A2(new_n736), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT100), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n738), .A2(new_n904), .A3(KEYINPUT31), .A4(new_n676), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n716), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT101), .B1(new_n873), .B2(new_n876), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n900), .B(new_n907), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  INV_X1    g0711(.A(new_n899), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n907), .A3(new_n877), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n423), .A2(new_n907), .ZN(new_n917));
  OAI21_X1  g0717(.A(G330), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n917), .B2(new_n916), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n898), .A2(new_n919), .B1(new_n284), .B2(new_n669), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n898), .B2(new_n919), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n922), .A2(G116), .A3(new_n210), .A4(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT36), .Z(new_n925));
  OAI211_X1 g0725(.A(new_n207), .B(G77), .C1(new_n202), .C2(new_n249), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n201), .A2(G68), .ZN(new_n927));
  AOI211_X1 g0727(.A(G13), .B(new_n284), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n921), .A2(new_n925), .A3(new_n928), .ZN(G367));
  OR2_X1    g0729(.A1(new_n597), .A2(new_n675), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n710), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT102), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n643), .B2(new_n930), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n931), .A2(KEYINPUT102), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n755), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n767), .B1(new_n213), .B2(new_n628), .C1(new_n237), .C2(new_n763), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n749), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n787), .A2(new_n843), .B1(new_n845), .B2(new_n783), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n273), .B1(new_n791), .B2(new_n389), .ZN(new_n940));
  XOR2_X1   g0740(.A(KEYINPUT105), .B(G137), .Z(new_n941));
  OAI22_X1  g0741(.A1(new_n782), .A2(new_n941), .B1(new_n793), .B2(new_n202), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n939), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n799), .A2(G150), .B1(G68), .B2(new_n796), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(new_n201), .C2(new_n788), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n799), .A2(G303), .B1(G283), .B2(new_n802), .ZN(new_n946));
  INV_X1    g0746(.A(new_n793), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT46), .B1(new_n947), .B2(G116), .ZN(new_n948));
  XNOR2_X1  g0748(.A(KEYINPUT104), .B(G311), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n948), .B1(new_n786), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n808), .A2(KEYINPUT46), .A3(G116), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n804), .A2(G317), .ZN(new_n953));
  INV_X1    g0753(.A(new_n791), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n273), .B1(new_n954), .B2(G97), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n776), .A2(G294), .B1(G107), .B2(new_n796), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n952), .A2(new_n953), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n945), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT47), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n938), .B1(new_n959), .B2(new_n766), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n936), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n692), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n689), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n692), .B1(new_n686), .B2(new_n688), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n682), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n682), .B1(new_n963), .B2(new_n964), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n714), .A2(new_n969), .A3(new_n742), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n547), .A2(new_n676), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n576), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT103), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n561), .A2(new_n676), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT103), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n576), .A2(new_n975), .A3(new_n971), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  OR3_X1    g0778(.A1(new_n977), .A2(new_n693), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n978), .B1(new_n977), .B2(new_n693), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n977), .A2(new_n693), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n977), .A2(KEYINPUT45), .A3(new_n693), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n691), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n981), .A2(new_n986), .A3(new_n691), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n970), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n744), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n696), .B(KEYINPUT41), .Z(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n748), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n973), .A2(new_n976), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n648), .B1(new_n996), .B2(new_n650), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n963), .A2(new_n977), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n997), .A2(new_n675), .B1(new_n998), .B2(KEYINPUT42), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(KEYINPUT42), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n935), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(KEYINPUT43), .B1(new_n933), .B2(new_n934), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .A4(new_n935), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n988), .A2(new_n977), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1005), .A2(new_n988), .A3(new_n977), .A4(new_n1006), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n961), .B1(new_n995), .B2(new_n1011), .ZN(G387));
  NAND3_X1  g0812(.A1(new_n743), .A2(new_n968), .A3(new_n967), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n714), .A2(new_n969), .A3(new_n742), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(new_n696), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n947), .A2(G77), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n844), .B2(new_n782), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n317), .B(new_n1017), .C1(G97), .C2(new_n954), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n802), .A2(G68), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n799), .A2(G50), .B1(new_n333), .B2(new_n776), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n786), .A2(G159), .B1(new_n377), .B2(new_n796), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n772), .A2(new_n806), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n799), .A2(G317), .B1(G322), .B2(new_n786), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n776), .A2(new_n949), .B1(new_n802), .B2(G303), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT48), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1023), .B(new_n1026), .C1(G294), .C2(new_n947), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(KEYINPUT48), .A3(new_n1025), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(KEYINPUT49), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n273), .B1(new_n804), .B2(G326), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(new_n426), .C2(new_n791), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT49), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1022), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n766), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n757), .A2(new_n698), .B1(new_n362), .B2(new_n695), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n234), .A2(new_n760), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n333), .A2(new_n201), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT50), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n699), .B(new_n760), .C1(new_n249), .C2(new_n389), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n762), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1035), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n832), .B1(new_n1041), .B2(new_n767), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1034), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n689), .B2(new_n755), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n969), .B2(new_n748), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1015), .A2(new_n1045), .ZN(G393));
  NAND3_X1  g0846(.A1(new_n989), .A2(new_n748), .A3(new_n990), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n996), .A2(new_n755), .A3(new_n974), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n799), .A2(G159), .B1(G150), .B2(new_n786), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT51), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n837), .A2(new_n317), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n249), .B2(new_n793), .C1(new_n843), .C2(new_n782), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n772), .A2(new_n389), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n845), .A2(new_n201), .B1(new_n332), .B2(new_n788), .ZN(new_n1054));
  NOR4_X1   g0854(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT106), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n799), .A2(G311), .B1(G317), .B2(new_n786), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT52), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n947), .A2(G283), .B1(new_n804), .B2(G322), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1060), .B(new_n317), .C1(new_n362), .C2(new_n791), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n776), .A2(G303), .B1(new_n802), .B2(G294), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n426), .B2(new_n772), .ZN(new_n1063));
  OR3_X1    g0863(.A1(new_n1059), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1056), .A2(KEYINPUT106), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1057), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n766), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n767), .B1(new_n429), .B2(new_n213), .C1(new_n245), .C2(new_n763), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1048), .A2(new_n749), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1047), .A2(new_n1069), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n981), .A2(new_n691), .A3(new_n986), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n691), .B1(new_n981), .B2(new_n986), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1014), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n991), .A2(new_n1073), .A3(new_n696), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT107), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n991), .A2(new_n1073), .A3(KEYINPUT107), .A4(new_n696), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1070), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(G390));
  AOI21_X1  g0879(.A(new_n881), .B1(new_n873), .B2(new_n876), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n709), .A2(new_n711), .A3(new_n643), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n561), .B(new_n613), .C1(new_n621), .C2(new_n631), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(KEYINPUT26), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n675), .B(new_n827), .C1(new_n1081), .C2(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1084), .A2(new_n887), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n893), .A2(new_n894), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1080), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n879), .A2(new_n882), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1086), .B1(new_n828), .B2(new_n887), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(new_n881), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n681), .B1(new_n716), .B2(new_n906), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1092), .A2(new_n912), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n517), .A2(new_n532), .A3(new_n675), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n740), .B1(new_n632), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1096), .A2(new_n895), .A3(G330), .A4(new_n822), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1087), .A2(new_n1090), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n822), .B1(new_n1092), .B2(KEYINPUT109), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT109), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1101), .B(new_n681), .C1(new_n716), .C2(new_n906), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1086), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1097), .A2(new_n1084), .A3(new_n887), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n895), .B1(new_n741), .B2(new_n822), .ZN(new_n1106));
  OAI211_X1 g0906(.A(KEYINPUT108), .B(new_n888), .C1(new_n1093), .C2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT108), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n828), .A2(new_n887), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1096), .A2(G330), .A3(new_n822), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1110), .A2(new_n1086), .B1(new_n1092), .B2(new_n912), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1108), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1105), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1092), .A2(new_n423), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n861), .A2(new_n666), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n697), .B1(new_n1099), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1094), .A2(new_n1098), .A3(new_n1116), .A4(new_n1113), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n799), .A2(G116), .B1(G283), .B2(new_n786), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n362), .B2(new_n845), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n273), .B(new_n848), .C1(G294), .C2(new_n804), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1053), .B1(new_n802), .B2(G97), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n808), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1123), .B(new_n1124), .C1(new_n792), .C2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n802), .A2(new_n1128), .B1(G159), .B2(new_n796), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n852), .B2(new_n779), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n791), .A2(new_n201), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n317), .B(new_n1131), .C1(G125), .C2(new_n804), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n793), .A2(new_n844), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1133), .B(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n941), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(G128), .A2(new_n786), .B1(new_n776), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1132), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1122), .A2(new_n1126), .B1(new_n1130), .B2(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1139), .A2(new_n766), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n833), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n749), .B1(new_n333), .B2(new_n1141), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(new_n1088), .C2(new_n753), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n1099), .B2(new_n747), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1120), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(G378));
  INV_X1    g0947(.A(KEYINPUT57), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1119), .A2(new_n1116), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n896), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n883), .A2(new_n885), .ZN(new_n1151));
  OAI21_X1  g0951(.A(KEYINPUT116), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(KEYINPUT117), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n915), .A2(G330), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n420), .A2(new_n674), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n422), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n413), .A2(new_n418), .A3(new_n421), .A4(new_n1155), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1159), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1154), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1162), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n915), .A2(G330), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT117), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n897), .A2(KEYINPUT116), .A3(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1153), .A2(new_n1163), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1166), .B1(new_n897), .B2(KEYINPUT116), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT116), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1170), .B(KEYINPUT117), .C1(new_n886), .C2(new_n896), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1164), .B1(new_n915), .B2(G330), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n915), .A2(G330), .A3(new_n1164), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n1169), .A2(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1168), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1148), .B1(new_n1149), .B2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1163), .A2(new_n896), .A3(new_n886), .A4(new_n1165), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n897), .B1(new_n1173), .B2(new_n1172), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1148), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1119), .A2(new_n1116), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n697), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n247), .A2(new_n449), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT111), .ZN(new_n1184));
  AOI211_X1 g0984(.A(G50), .B(new_n1184), .C1(new_n449), .C2(new_n317), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n786), .A2(G116), .B1(new_n802), .B2(new_n377), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n362), .B2(new_n779), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n791), .A2(new_n202), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G283), .B2(new_n804), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1189), .A2(new_n449), .A3(new_n317), .A4(new_n1016), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n845), .A2(new_n429), .B1(new_n249), .B2(new_n772), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1187), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT112), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT58), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1185), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1194), .B2(new_n1193), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n799), .A2(G128), .B1(G137), .B2(new_n802), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n947), .A2(new_n1128), .B1(new_n796), .B2(G150), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G125), .A2(new_n786), .B1(new_n776), .B2(G132), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT113), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n804), .A2(G124), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1204), .B(new_n1184), .C1(new_n783), .C2(new_n791), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT114), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1202), .A2(new_n1203), .A3(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n766), .B1(new_n1196), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n749), .C1(G50), .C2(new_n1141), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1162), .B2(new_n753), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT115), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n1175), .B2(new_n747), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1182), .A2(new_n1213), .ZN(G375));
  NAND2_X1  g1014(.A1(new_n1113), .A2(new_n748), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n799), .A2(new_n1136), .B1(new_n776), .B2(new_n1128), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n317), .B(new_n1188), .C1(G128), .C2(new_n804), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n783), .C2(new_n1125), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n802), .A2(G150), .B1(G50), .B2(new_n796), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n852), .B2(new_n787), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n799), .A2(G283), .B1(G294), .B2(new_n786), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n426), .B2(new_n845), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n317), .B1(new_n791), .B2(new_n389), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G303), .B2(new_n804), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n802), .A2(G107), .B1(new_n377), .B2(new_n796), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n1125), .C2(new_n429), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1218), .A2(new_n1220), .B1(new_n1222), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n766), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n832), .B1(new_n249), .B2(new_n833), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(new_n895), .C2(new_n754), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1215), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1115), .A2(new_n1105), .A3(new_n1107), .A4(new_n1112), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1117), .A2(new_n994), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(G381));
  AOI21_X1  g1035(.A(new_n1212), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1146), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1071), .A2(new_n1014), .A3(new_n1072), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n994), .B1(new_n1239), .B2(new_n743), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n747), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1241), .A2(new_n1242), .B1(new_n936), .B2(new_n960), .ZN(new_n1243));
  INV_X1    g1043(.A(G384), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(G393), .A2(G396), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1246), .A2(G390), .A3(G381), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1238), .A2(new_n1247), .ZN(G407));
  INV_X1    g1048(.A(G213), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(G343), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1238), .A2(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT118), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1249), .B1(new_n1238), .B2(new_n1247), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(KEYINPUT119), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT119), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1252), .A2(new_n1256), .A3(new_n1253), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(G409));
  NAND3_X1  g1058(.A1(G390), .A2(new_n1243), .A3(KEYINPUT124), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(G393), .B(new_n813), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G387), .B2(new_n1078), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT124), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(G387), .B2(new_n1078), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1259), .A2(new_n1261), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT125), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1259), .A2(new_n1261), .A3(KEYINPUT125), .A4(new_n1263), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G387), .B(new_n1078), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1260), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1250), .A2(G2897), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1233), .A2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(new_n697), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1233), .A2(new_n1275), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1278), .A2(KEYINPUT122), .A3(new_n1117), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT122), .B1(new_n1278), .B2(new_n1117), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1277), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT123), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI211_X1 g1083(.A(KEYINPUT123), .B(new_n1277), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G384), .B1(new_n1285), .B2(new_n1232), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n1244), .B(new_n1231), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1274), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1278), .A2(new_n1117), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT122), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1278), .A2(KEYINPUT122), .A3(new_n1117), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT123), .B1(new_n1293), .B2(new_n1277), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1284), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1232), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1244), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1285), .A2(G384), .A3(new_n1232), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1273), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1250), .B1(G375), .B2(G378), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1180), .A2(new_n994), .A3(new_n1168), .A4(new_n1174), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT120), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n747), .B1(new_n1303), .B2(KEYINPUT121), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT121), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1177), .A2(new_n1178), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1210), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1168), .A2(new_n1174), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT120), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1308), .A2(new_n1309), .A3(new_n994), .A4(new_n1180), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1146), .A2(new_n1302), .A3(new_n1307), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1300), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1288), .A2(new_n1299), .A3(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT126), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1316));
  OAI21_X1  g1116(.A(KEYINPUT62), .B1(new_n1312), .B2(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1250), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1319), .B1(new_n1236), .B2(new_n1146), .ZN(new_n1320));
  AND4_X1   g1120(.A1(new_n1146), .A2(new_n1302), .A3(new_n1307), .A4(new_n1310), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1318), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1317), .A2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1272), .B1(new_n1315), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT126), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1268), .A2(new_n1327), .A3(new_n1270), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1313), .A2(new_n1314), .A3(new_n1328), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1318), .A2(new_n1322), .A3(KEYINPUT63), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT63), .B1(new_n1318), .B2(new_n1322), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1271), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1329), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1326), .A2(new_n1333), .ZN(G405));
  NOR2_X1   g1134(.A1(new_n1236), .A2(new_n1146), .ZN(new_n1335));
  OR3_X1    g1135(.A1(new_n1318), .A2(new_n1238), .A3(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1318), .B1(new_n1238), .B2(new_n1335), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT127), .ZN(new_n1338));
  AOI22_X1  g1138(.A1(new_n1336), .A2(new_n1337), .B1(new_n1271), .B2(new_n1338), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(new_n1271), .B(new_n1338), .ZN(new_n1340));
  AND2_X1   g1140(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1339), .B1(new_n1340), .B2(new_n1341), .ZN(G402));
endmodule


