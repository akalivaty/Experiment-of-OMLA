

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593;

  XNOR2_X1 U324 ( .A(n524), .B(n523), .ZN(n555) );
  INV_X1 U325 ( .A(n580), .ZN(n540) );
  XOR2_X1 U326 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n292) );
  XOR2_X1 U327 ( .A(KEYINPUT87), .B(G176GAT), .Z(n293) );
  XNOR2_X1 U328 ( .A(n432), .B(n431), .ZN(n441) );
  XNOR2_X1 U329 ( .A(n522), .B(KEYINPUT48), .ZN(n523) );
  XNOR2_X1 U330 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U331 ( .A(n342), .B(n293), .ZN(n343) );
  XNOR2_X1 U332 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U333 ( .A(n366), .B(KEYINPUT26), .ZN(n580) );
  XOR2_X1 U334 ( .A(n445), .B(n444), .Z(n584) );
  INV_X1 U335 ( .A(KEYINPUT111), .ZN(n500) );
  XNOR2_X1 U336 ( .A(n349), .B(n348), .ZN(n350) );
  NOR2_X1 U337 ( .A1(n562), .A2(n561), .ZN(n572) );
  XNOR2_X1 U338 ( .A(n501), .B(n500), .ZN(n507) );
  XNOR2_X1 U339 ( .A(n351), .B(n350), .ZN(n562) );
  XOR2_X1 U340 ( .A(G155GAT), .B(G148GAT), .Z(n295) );
  XNOR2_X1 U341 ( .A(G1GAT), .B(G127GAT), .ZN(n294) );
  XNOR2_X1 U342 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U343 ( .A(G85GAT), .B(G162GAT), .Z(n297) );
  XNOR2_X1 U344 ( .A(G29GAT), .B(G120GAT), .ZN(n296) );
  XNOR2_X1 U345 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n316) );
  XOR2_X1 U347 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n301) );
  XNOR2_X1 U348 ( .A(G57GAT), .B(KEYINPUT97), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U350 ( .A(KEYINPUT96), .B(KEYINPUT1), .Z(n303) );
  XNOR2_X1 U351 ( .A(KEYINPUT6), .B(KEYINPUT98), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U353 ( .A(n305), .B(n304), .Z(n314) );
  XOR2_X1 U354 ( .A(KEYINPUT2), .B(KEYINPUT93), .Z(n307) );
  XNOR2_X1 U355 ( .A(KEYINPUT3), .B(KEYINPUT92), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U357 ( .A(G141GAT), .B(n308), .Z(n335) );
  XOR2_X1 U358 ( .A(G134GAT), .B(KEYINPUT80), .Z(n413) );
  XNOR2_X1 U359 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n309), .B(KEYINPUT86), .ZN(n342) );
  XOR2_X1 U361 ( .A(n413), .B(n342), .Z(n311) );
  NAND2_X1 U362 ( .A1(G225GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n335), .B(n312), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n557) );
  XOR2_X1 U367 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n318) );
  XNOR2_X1 U368 ( .A(G197GAT), .B(G211GAT), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n320) );
  XNOR2_X1 U370 ( .A(G218GAT), .B(KEYINPUT91), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n352) );
  XOR2_X1 U372 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n322) );
  XNOR2_X1 U373 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U375 ( .A(n323), .B(KEYINPUT24), .Z(n325) );
  XOR2_X1 U376 ( .A(G22GAT), .B(G155GAT), .Z(n385) );
  XNOR2_X1 U377 ( .A(n385), .B(KEYINPUT94), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n330) );
  XNOR2_X1 U379 ( .A(G50GAT), .B(KEYINPUT77), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n326), .B(G162GAT), .ZN(n418) );
  XOR2_X1 U381 ( .A(n418), .B(KEYINPUT95), .Z(n328) );
  NAND2_X1 U382 ( .A1(G228GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U384 ( .A(n330), .B(n329), .Z(n337) );
  XNOR2_X1 U385 ( .A(G148GAT), .B(KEYINPUT72), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n331), .B(KEYINPUT73), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n332), .B(G204GAT), .ZN(n334) );
  XOR2_X1 U388 ( .A(G78GAT), .B(G106GAT), .Z(n333) );
  XOR2_X1 U389 ( .A(n334), .B(n333), .Z(n444) );
  XOR2_X1 U390 ( .A(n444), .B(n335), .Z(n336) );
  XNOR2_X1 U391 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U392 ( .A(n352), .B(n338), .Z(n559) );
  XOR2_X1 U393 ( .A(G120GAT), .B(G71GAT), .Z(n431) );
  XNOR2_X1 U394 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n292), .B(n339), .ZN(n358) );
  XOR2_X1 U396 ( .A(n431), .B(n358), .Z(n341) );
  NAND2_X1 U397 ( .A1(G227GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n344) );
  XOR2_X1 U399 ( .A(G15GAT), .B(G127GAT), .Z(n395) );
  XOR2_X1 U400 ( .A(n345), .B(n395), .Z(n351) );
  XOR2_X1 U401 ( .A(G183GAT), .B(KEYINPUT20), .Z(n347) );
  XNOR2_X1 U402 ( .A(G99GAT), .B(G190GAT), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n349) );
  XNOR2_X1 U404 ( .A(G43GAT), .B(G134GAT), .ZN(n348) );
  XOR2_X1 U405 ( .A(G36GAT), .B(G190GAT), .Z(n406) );
  XOR2_X1 U406 ( .A(G8GAT), .B(G183GAT), .Z(n386) );
  XOR2_X1 U407 ( .A(KEYINPUT99), .B(n386), .Z(n354) );
  XNOR2_X1 U408 ( .A(n352), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n406), .B(n355), .ZN(n357) );
  AND2_X1 U411 ( .A1(G226GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n359) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n361) );
  XNOR2_X1 U414 ( .A(G176GAT), .B(G92GAT), .ZN(n360) );
  XOR2_X1 U415 ( .A(n360), .B(G64GAT), .Z(n430) );
  XNOR2_X1 U416 ( .A(n361), .B(n430), .ZN(n365) );
  INV_X1 U417 ( .A(n365), .ZN(n362) );
  INV_X1 U418 ( .A(n362), .ZN(n554) );
  NOR2_X1 U419 ( .A1(n562), .A2(n554), .ZN(n363) );
  NOR2_X1 U420 ( .A1(n559), .A2(n363), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n364), .B(KEYINPUT25), .ZN(n368) );
  XNOR2_X1 U422 ( .A(KEYINPUT27), .B(n365), .ZN(n371) );
  NAND2_X1 U423 ( .A1(n562), .A2(n559), .ZN(n366) );
  OR2_X1 U424 ( .A1(n371), .A2(n580), .ZN(n367) );
  NAND2_X1 U425 ( .A1(n368), .A2(n367), .ZN(n369) );
  NAND2_X1 U426 ( .A1(n369), .A2(n557), .ZN(n377) );
  XNOR2_X1 U427 ( .A(n559), .B(KEYINPUT67), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n370), .B(KEYINPUT28), .ZN(n528) );
  NOR2_X1 U429 ( .A1(n371), .A2(n557), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n372), .B(KEYINPUT100), .ZN(n525) );
  NAND2_X1 U431 ( .A1(n528), .A2(n525), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n373), .B(KEYINPUT101), .ZN(n374) );
  NAND2_X1 U433 ( .A1(n374), .A2(n562), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n375), .B(KEYINPUT102), .ZN(n376) );
  NAND2_X1 U435 ( .A1(n377), .A2(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n378), .B(KEYINPUT103), .ZN(n472) );
  XOR2_X1 U437 ( .A(KEYINPUT15), .B(KEYINPUT84), .Z(n380) );
  XNOR2_X1 U438 ( .A(G64GAT), .B(KEYINPUT85), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U440 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n382) );
  XNOR2_X1 U441 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n403) );
  XOR2_X1 U444 ( .A(n386), .B(n385), .Z(n388) );
  XNOR2_X1 U445 ( .A(G71GAT), .B(G78GAT), .ZN(n387) );
  XNOR2_X1 U446 ( .A(n388), .B(n387), .ZN(n399) );
  INV_X1 U447 ( .A(KEYINPUT70), .ZN(n389) );
  NAND2_X1 U448 ( .A1(KEYINPUT13), .A2(n389), .ZN(n392) );
  INV_X1 U449 ( .A(KEYINPUT13), .ZN(n390) );
  NAND2_X1 U450 ( .A1(n390), .A2(KEYINPUT70), .ZN(n391) );
  NAND2_X1 U451 ( .A1(n392), .A2(n391), .ZN(n394) );
  XNOR2_X1 U452 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n433) );
  XOR2_X1 U454 ( .A(n433), .B(n395), .Z(n397) );
  NAND2_X1 U455 ( .A1(G231GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U457 ( .A(n399), .B(n398), .Z(n401) );
  XNOR2_X1 U458 ( .A(G1GAT), .B(G211GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n548) );
  XOR2_X1 U461 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n405) );
  XNOR2_X1 U462 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U464 ( .A(n407), .B(n406), .Z(n409) );
  XNOR2_X1 U465 ( .A(G218GAT), .B(G106GAT), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U467 ( .A(G99GAT), .B(G85GAT), .Z(n429) );
  XOR2_X1 U468 ( .A(n410), .B(n429), .Z(n415) );
  XOR2_X1 U469 ( .A(G29GAT), .B(G43GAT), .Z(n412) );
  XNOR2_X1 U470 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n450) );
  XNOR2_X1 U472 ( .A(n450), .B(n413), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n424) );
  XOR2_X1 U474 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n417) );
  XNOR2_X1 U475 ( .A(KEYINPUT78), .B(KEYINPUT11), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n422) );
  XOR2_X1 U477 ( .A(KEYINPUT9), .B(n418), .Z(n420) );
  NAND2_X1 U478 ( .A1(G232GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U480 ( .A(n422), .B(n421), .Z(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n571) );
  NOR2_X1 U482 ( .A1(n548), .A2(n571), .ZN(n425) );
  XOR2_X1 U483 ( .A(KEYINPUT16), .B(n425), .Z(n426) );
  NOR2_X1 U484 ( .A1(n472), .A2(n426), .ZN(n485) );
  XOR2_X1 U485 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n428) );
  XNOR2_X1 U486 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n427) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n443) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n432) );
  NAND2_X1 U489 ( .A1(n433), .A2(KEYINPUT31), .ZN(n437) );
  INV_X1 U490 ( .A(n433), .ZN(n435) );
  INV_X1 U491 ( .A(KEYINPUT31), .ZN(n434) );
  NAND2_X1 U492 ( .A1(n435), .A2(n434), .ZN(n436) );
  NAND2_X1 U493 ( .A1(n437), .A2(n436), .ZN(n439) );
  AND2_X1 U494 ( .A1(G230GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U497 ( .A(G141GAT), .B(G113GAT), .Z(n447) );
  XNOR2_X1 U498 ( .A(G169GAT), .B(G15GAT), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n461) );
  XOR2_X1 U500 ( .A(G50GAT), .B(G36GAT), .Z(n449) );
  NAND2_X1 U501 ( .A1(G229GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n451) );
  XOR2_X1 U503 ( .A(n451), .B(n450), .Z(n459) );
  XOR2_X1 U504 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n453) );
  XNOR2_X1 U505 ( .A(G22GAT), .B(G197GAT), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n457) );
  XOR2_X1 U507 ( .A(G1GAT), .B(KEYINPUT29), .Z(n455) );
  XNOR2_X1 U508 ( .A(KEYINPUT69), .B(G8GAT), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U511 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n461), .B(n460), .ZN(n581) );
  INV_X1 U513 ( .A(n581), .ZN(n541) );
  NOR2_X1 U514 ( .A1(n584), .A2(n541), .ZN(n462) );
  XNOR2_X1 U515 ( .A(n462), .B(KEYINPUT76), .ZN(n474) );
  NAND2_X1 U516 ( .A1(n485), .A2(n474), .ZN(n468) );
  NOR2_X1 U517 ( .A1(n557), .A2(n468), .ZN(n463) );
  XOR2_X1 U518 ( .A(KEYINPUT34), .B(n463), .Z(n464) );
  XNOR2_X1 U519 ( .A(G1GAT), .B(n464), .ZN(G1324GAT) );
  NOR2_X1 U520 ( .A1(n554), .A2(n468), .ZN(n465) );
  XOR2_X1 U521 ( .A(G8GAT), .B(n465), .Z(G1325GAT) );
  NOR2_X1 U522 ( .A1(n562), .A2(n468), .ZN(n467) );
  XNOR2_X1 U523 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n467), .B(n466), .ZN(G1326GAT) );
  NOR2_X1 U525 ( .A1(n528), .A2(n468), .ZN(n469) );
  XOR2_X1 U526 ( .A(G22GAT), .B(n469), .Z(G1327GAT) );
  INV_X1 U527 ( .A(n548), .ZN(n588) );
  XNOR2_X1 U528 ( .A(KEYINPUT36), .B(n571), .ZN(n590) );
  INV_X1 U529 ( .A(n590), .ZN(n470) );
  OR2_X1 U530 ( .A1(n588), .A2(n470), .ZN(n471) );
  OR2_X1 U531 ( .A1(n472), .A2(n471), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(KEYINPUT37), .ZN(n499) );
  NAND2_X1 U533 ( .A1(n474), .A2(n499), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT38), .ZN(n482) );
  NOR2_X1 U535 ( .A1(n557), .A2(n482), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n476), .B(KEYINPUT39), .ZN(n477) );
  XNOR2_X1 U537 ( .A(G29GAT), .B(n477), .ZN(G1328GAT) );
  NOR2_X1 U538 ( .A1(n482), .A2(n554), .ZN(n478) );
  XOR2_X1 U539 ( .A(G36GAT), .B(n478), .Z(G1329GAT) );
  NOR2_X1 U540 ( .A1(n482), .A2(n562), .ZN(n480) );
  XNOR2_X1 U541 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U543 ( .A(G43GAT), .B(n481), .Z(G1330GAT) );
  NOR2_X1 U544 ( .A1(n528), .A2(n482), .ZN(n483) );
  XOR2_X1 U545 ( .A(G50GAT), .B(n483), .Z(G1331GAT) );
  XNOR2_X1 U546 ( .A(KEYINPUT41), .B(n584), .ZN(n545) );
  INV_X1 U547 ( .A(n545), .ZN(n567) );
  NAND2_X1 U548 ( .A1(n567), .A2(n541), .ZN(n484) );
  XOR2_X1 U549 ( .A(KEYINPUT106), .B(n484), .Z(n498) );
  NAND2_X1 U550 ( .A1(n485), .A2(n498), .ZN(n493) );
  NOR2_X1 U551 ( .A1(n493), .A2(n557), .ZN(n489) );
  XOR2_X1 U552 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n487) );
  XNOR2_X1 U553 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n486) );
  XNOR2_X1 U554 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U555 ( .A(n489), .B(n488), .ZN(G1332GAT) );
  NOR2_X1 U556 ( .A1(n554), .A2(n493), .ZN(n490) );
  XOR2_X1 U557 ( .A(KEYINPUT108), .B(n490), .Z(n491) );
  XNOR2_X1 U558 ( .A(G64GAT), .B(n491), .ZN(G1333GAT) );
  NOR2_X1 U559 ( .A1(n562), .A2(n493), .ZN(n492) );
  XOR2_X1 U560 ( .A(G71GAT), .B(n492), .Z(G1334GAT) );
  NOR2_X1 U561 ( .A1(n493), .A2(n528), .ZN(n497) );
  XOR2_X1 U562 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n495) );
  XNOR2_X1 U563 ( .A(G78GAT), .B(KEYINPUT110), .ZN(n494) );
  XNOR2_X1 U564 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U565 ( .A(n497), .B(n496), .ZN(G1335GAT) );
  NAND2_X1 U566 ( .A1(n499), .A2(n498), .ZN(n501) );
  NOR2_X1 U567 ( .A1(n557), .A2(n507), .ZN(n502) );
  XOR2_X1 U568 ( .A(G85GAT), .B(n502), .Z(G1336GAT) );
  NOR2_X1 U569 ( .A1(n554), .A2(n507), .ZN(n503) );
  XOR2_X1 U570 ( .A(G92GAT), .B(n503), .Z(G1337GAT) );
  NOR2_X1 U571 ( .A1(n562), .A2(n507), .ZN(n505) );
  XNOR2_X1 U572 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U574 ( .A(G99GAT), .B(n506), .ZN(G1338GAT) );
  NOR2_X1 U575 ( .A1(n507), .A2(n528), .ZN(n509) );
  XNOR2_X1 U576 ( .A(KEYINPUT44), .B(KEYINPUT114), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U578 ( .A(n510), .B(G106GAT), .Z(G1339GAT) );
  NAND2_X1 U579 ( .A1(n567), .A2(n581), .ZN(n511) );
  XNOR2_X1 U580 ( .A(KEYINPUT46), .B(n511), .ZN(n513) );
  NOR2_X1 U581 ( .A1(n571), .A2(n588), .ZN(n512) );
  AND2_X1 U582 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U583 ( .A(KEYINPUT47), .B(n514), .ZN(n521) );
  XOR2_X1 U584 ( .A(KEYINPUT45), .B(KEYINPUT115), .Z(n516) );
  NAND2_X1 U585 ( .A1(n590), .A2(n588), .ZN(n515) );
  XNOR2_X1 U586 ( .A(n516), .B(n515), .ZN(n517) );
  NOR2_X1 U587 ( .A1(n584), .A2(n517), .ZN(n518) );
  XNOR2_X1 U588 ( .A(KEYINPUT116), .B(n518), .ZN(n519) );
  NAND2_X1 U589 ( .A1(n519), .A2(n541), .ZN(n520) );
  NAND2_X1 U590 ( .A1(n521), .A2(n520), .ZN(n524) );
  XNOR2_X1 U591 ( .A(KEYINPUT64), .B(KEYINPUT117), .ZN(n522) );
  INV_X1 U592 ( .A(n525), .ZN(n526) );
  NOR2_X1 U593 ( .A1(n555), .A2(n526), .ZN(n527) );
  XNOR2_X1 U594 ( .A(KEYINPUT118), .B(n527), .ZN(n539) );
  NAND2_X1 U595 ( .A1(n528), .A2(n539), .ZN(n529) );
  NOR2_X1 U596 ( .A1(n562), .A2(n529), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n536), .A2(n581), .ZN(n530) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U600 ( .A1(n536), .A2(n567), .ZN(n531) );
  XNOR2_X1 U601 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n534) );
  NAND2_X1 U603 ( .A1(n536), .A2(n588), .ZN(n533) );
  XNOR2_X1 U604 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U607 ( .A1(n536), .A2(n571), .ZN(n537) );
  XNOR2_X1 U608 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n540), .A2(n539), .ZN(n551) );
  NOR2_X1 U610 ( .A1(n541), .A2(n551), .ZN(n542) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n542), .Z(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n544) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n544), .B(n543), .ZN(n547) );
  NOR2_X1 U615 ( .A1(n545), .A2(n551), .ZN(n546) );
  XOR2_X1 U616 ( .A(n547), .B(n546), .Z(G1345GAT) );
  NOR2_X1 U617 ( .A1(n548), .A2(n551), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(G1346GAT) );
  INV_X1 U620 ( .A(n571), .ZN(n552) );
  NOR2_X1 U621 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n553), .Z(G1347GAT) );
  NOR2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(KEYINPUT54), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n579) );
  NOR2_X1 U626 ( .A1(n559), .A2(n579), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT55), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n572), .A2(n581), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n565) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(n566), .Z(n569) );
  NAND2_X1 U634 ( .A1(n572), .A2(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NAND2_X1 U636 ( .A1(n588), .A2(n572), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U638 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1351GAT) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n577), .B(KEYINPUT60), .ZN(n578) );
  XOR2_X1 U645 ( .A(KEYINPUT59), .B(n578), .Z(n583) );
  NOR2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n591) );
  NAND2_X1 U647 ( .A1(n591), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n586) );
  NAND2_X1 U650 ( .A1(n591), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U652 ( .A(G204GAT), .B(n587), .Z(G1353GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n591), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(n592), .B(KEYINPUT62), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

