

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821;

  NOR2_X1 U372 ( .A1(n796), .A2(n701), .ZN(n783) );
  NOR2_X1 U373 ( .A1(n679), .A2(n680), .ZN(n474) );
  BUF_X1 U374 ( .A(n388), .Z(n385) );
  AND2_X1 U375 ( .A1(n475), .A2(n420), .ZN(n662) );
  XNOR2_X2 U376 ( .A(n700), .B(n694), .ZN(n696) );
  XNOR2_X2 U377 ( .A(n683), .B(n682), .ZN(n487) );
  NAND2_X2 U378 ( .A1(n350), .A2(n533), .ZN(n535) );
  XNOR2_X2 U379 ( .A(n659), .B(KEYINPUT19), .ZN(n350) );
  NOR2_X1 U380 ( .A1(G953), .A2(G237), .ZN(n577) );
  XOR2_X1 U381 ( .A(G113), .B(G104), .Z(n404) );
  XNOR2_X1 U382 ( .A(n662), .B(KEYINPUT88), .ZN(n741) );
  BUF_X1 U383 ( .A(G104), .Z(n424) );
  XNOR2_X1 U384 ( .A(n465), .B(KEYINPUT62), .ZN(n351) );
  XNOR2_X2 U385 ( .A(G134), .B(KEYINPUT72), .ZN(n464) );
  NAND2_X2 U386 ( .A1(n481), .A2(n479), .ZN(n700) );
  XNOR2_X2 U387 ( .A(n383), .B(n536), .ZN(n620) );
  XNOR2_X2 U388 ( .A(n576), .B(n575), .ZN(n750) );
  AND2_X2 U389 ( .A1(n573), .A2(n388), .ZN(n576) );
  NAND2_X2 U390 ( .A1(n465), .A2(n548), .ZN(n558) );
  INV_X2 U391 ( .A(G953), .ZN(n812) );
  AND2_X1 U392 ( .A1(n354), .A2(n396), .ZN(n353) );
  INV_X1 U393 ( .A(n362), .ZN(n356) );
  XNOR2_X1 U394 ( .A(n684), .B(n473), .ZN(n362) );
  AND2_X1 U395 ( .A1(n628), .A2(n627), .ZN(n655) );
  XNOR2_X2 U396 ( .A(G110), .B(KEYINPUT77), .ZN(n512) );
  XNOR2_X1 U397 ( .A(n352), .B(n351), .ZN(n511) );
  NAND2_X1 U398 ( .A1(n364), .A2(n365), .ZN(n352) );
  NAND2_X1 U399 ( .A1(n444), .A2(n353), .ZN(n392) );
  AND2_X1 U400 ( .A1(G472), .A2(n702), .ZN(n365) );
  NAND2_X1 U401 ( .A1(n419), .A2(KEYINPUT91), .ZN(n354) );
  NAND2_X1 U402 ( .A1(n449), .A2(n448), .ZN(n447) );
  AND2_X1 U403 ( .A1(n485), .A2(n482), .ZN(n481) );
  XNOR2_X1 U404 ( .A(n644), .B(KEYINPUT40), .ZN(n709) );
  NAND2_X1 U405 ( .A1(n357), .A2(n355), .ZN(n708) );
  NAND2_X1 U406 ( .A1(n643), .A2(n655), .ZN(n644) );
  AND2_X1 U407 ( .A1(n360), .A2(n358), .ZN(n357) );
  NAND2_X1 U408 ( .A1(n356), .A2(KEYINPUT36), .ZN(n355) );
  NAND2_X1 U409 ( .A1(n362), .A2(n361), .ZN(n360) );
  AND2_X1 U410 ( .A1(n385), .A2(n359), .ZN(n358) );
  AND2_X1 U411 ( .A1(n493), .A2(n492), .ZN(n491) );
  OR2_X1 U412 ( .A1(n472), .A2(n660), .ZN(n359) );
  BUF_X1 U413 ( .A(n725), .Z(n366) );
  XNOR2_X1 U414 ( .A(n591), .B(n590), .ZN(n628) );
  XNOR2_X1 U415 ( .A(n512), .B(KEYINPUT76), .ZN(n537) );
  XOR2_X1 U416 ( .A(G122), .B(G107), .Z(n592) );
  XNOR2_X1 U417 ( .A(n441), .B(n507), .ZN(n606) );
  XNOR2_X2 U418 ( .A(n648), .B(KEYINPUT1), .ZN(n388) );
  NAND2_X1 U419 ( .A1(n354), .A2(n417), .ZN(n390) );
  AND2_X1 U420 ( .A1(n472), .A2(n660), .ZN(n361) );
  INV_X2 U421 ( .A(G125), .ZN(n398) );
  BUF_X1 U422 ( .A(n393), .Z(n363) );
  AND2_X1 U423 ( .A1(n440), .A2(KEYINPUT66), .ZN(n391) );
  NAND2_X1 U424 ( .A1(n363), .A2(n392), .ZN(n364) );
  BUF_X1 U425 ( .A(n642), .Z(n691) );
  OR2_X2 U426 ( .A1(n642), .A2(n685), .ZN(n659) );
  XNOR2_X1 U427 ( .A(n525), .B(n524), .ZN(n642) );
  NAND2_X1 U428 ( .A1(n369), .A2(n427), .ZN(n426) );
  XNOR2_X1 U429 ( .A(n608), .B(KEYINPUT109), .ZN(n755) );
  XNOR2_X1 U430 ( .A(n569), .B(n568), .ZN(n766) );
  OR2_X1 U431 ( .A1(n741), .A2(n663), .ZN(n665) );
  INV_X1 U432 ( .A(n430), .ZN(n551) );
  AND2_X1 U433 ( .A1(n483), .A2(n748), .ZN(n482) );
  NAND2_X1 U434 ( .A1(n484), .A2(KEYINPUT94), .ZN(n483) );
  INV_X1 U435 ( .A(n705), .ZN(n484) );
  INV_X1 U436 ( .A(n729), .ZN(n503) );
  INV_X1 U437 ( .A(KEYINPUT79), .ZN(n498) );
  AND2_X1 U438 ( .A1(n379), .A2(n418), .ZN(n417) );
  XNOR2_X1 U439 ( .A(n531), .B(KEYINPUT101), .ZN(n634) );
  INV_X1 U440 ( .A(G146), .ZN(n382) );
  XNOR2_X1 U441 ( .A(G119), .B(G116), .ZN(n521) );
  XNOR2_X1 U442 ( .A(G101), .B(G107), .ZN(n539) );
  INV_X1 U443 ( .A(n424), .ZN(n541) );
  NAND2_X1 U444 ( .A1(n489), .A2(n368), .ZN(n488) );
  INV_X1 U445 ( .A(n691), .ZN(n469) );
  NOR2_X1 U446 ( .A1(n450), .A2(n437), .ZN(n638) );
  INV_X1 U447 ( .A(n645), .ZN(n437) );
  XNOR2_X1 U448 ( .A(n641), .B(n640), .ZN(n670) );
  INV_X1 U449 ( .A(KEYINPUT28), .ZN(n476) );
  NOR2_X1 U450 ( .A1(G902), .A2(n718), .ZN(n591) );
  NAND2_X1 U451 ( .A1(n471), .A2(n446), .ZN(n631) );
  INV_X1 U452 ( .A(n616), .ZN(n471) );
  XNOR2_X1 U453 ( .A(n783), .B(n506), .ZN(n505) );
  XNOR2_X1 U454 ( .A(KEYINPUT92), .B(KEYINPUT2), .ZN(n506) );
  XNOR2_X1 U455 ( .A(n708), .B(KEYINPUT95), .ZN(n680) );
  AND2_X1 U456 ( .A1(n457), .A2(n377), .ZN(n456) );
  INV_X1 U457 ( .A(n746), .ZN(n463) );
  INV_X1 U458 ( .A(KEYINPUT68), .ZN(n501) );
  XNOR2_X1 U459 ( .A(n593), .B(n401), .ZN(n384) );
  XNOR2_X1 U460 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n401) );
  AND2_X1 U461 ( .A1(n451), .A2(n438), .ZN(n573) );
  INV_X1 U462 ( .A(G237), .ZN(n523) );
  XOR2_X1 U463 ( .A(KEYINPUT103), .B(KEYINPUT20), .Z(n566) );
  XNOR2_X1 U464 ( .A(KEYINPUT83), .B(KEYINPUT5), .ZN(n553) );
  NAND2_X1 U465 ( .A1(n480), .A2(KEYINPUT94), .ZN(n479) );
  XNOR2_X1 U466 ( .A(KEYINPUT93), .B(KEYINPUT45), .ZN(n633) );
  AND2_X1 U467 ( .A1(n632), .A2(n375), .ZN(n502) );
  XNOR2_X1 U468 ( .A(n399), .B(n384), .ZN(n453) );
  XNOR2_X1 U469 ( .A(n439), .B(n400), .ZN(n399) );
  NAND2_X1 U470 ( .A1(n812), .A2(G224), .ZN(n400) );
  XNOR2_X1 U471 ( .A(KEYINPUT18), .B(KEYINPUT86), .ZN(n517) );
  AND2_X1 U472 ( .A1(n417), .A2(n397), .ZN(n396) );
  INV_X1 U473 ( .A(KEYINPUT66), .ZN(n397) );
  XNOR2_X1 U474 ( .A(n428), .B(n527), .ZN(n530) );
  XNOR2_X1 U475 ( .A(KEYINPUT82), .B(KEYINPUT14), .ZN(n428) );
  NAND2_X1 U476 ( .A1(n752), .A2(n496), .ZN(n495) );
  NAND2_X1 U477 ( .A1(n490), .A2(n752), .ZN(n489) );
  NOR2_X1 U478 ( .A1(n766), .A2(n646), .ZN(n656) );
  XNOR2_X1 U479 ( .A(G110), .B(KEYINPUT24), .ZN(n435) );
  XNOR2_X1 U480 ( .A(n433), .B(KEYINPUT23), .ZN(n432) );
  XNOR2_X1 U481 ( .A(G119), .B(G137), .ZN(n433) );
  XOR2_X1 U482 ( .A(KEYINPUT108), .B(KEYINPUT11), .Z(n579) );
  XNOR2_X1 U483 ( .A(G143), .B(G122), .ZN(n580) );
  XOR2_X1 U484 ( .A(KEYINPUT12), .B(G140), .Z(n581) );
  INV_X1 U485 ( .A(KEYINPUT114), .ZN(n473) );
  INV_X1 U486 ( .A(KEYINPUT35), .ZN(n507) );
  XNOR2_X1 U487 ( .A(n611), .B(KEYINPUT22), .ZN(n616) );
  INV_X1 U488 ( .A(n592), .ZN(n455) );
  XOR2_X1 U489 ( .A(G116), .B(KEYINPUT9), .Z(n598) );
  XNOR2_X1 U490 ( .A(n542), .B(n541), .ZN(n543) );
  NOR2_X1 U491 ( .A1(n776), .A2(n421), .ZN(n651) );
  NOR2_X1 U492 ( .A1(n631), .A2(n612), .ZN(n614) );
  BUF_X1 U493 ( .A(G113), .Z(n430) );
  AND2_X1 U494 ( .A1(n670), .A2(n468), .ZN(n672) );
  AND2_X1 U495 ( .A1(n671), .A2(n469), .ZN(n468) );
  NOR2_X1 U496 ( .A1(n661), .A2(n649), .ZN(n420) );
  NAND2_X1 U497 ( .A1(n387), .A2(n386), .ZN(n630) );
  INV_X1 U498 ( .A(n629), .ZN(n386) );
  AND2_X1 U499 ( .A1(n505), .A2(n371), .ZN(n784) );
  AND2_X1 U500 ( .A1(n376), .A2(n388), .ZN(n367) );
  XNOR2_X1 U501 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n368) );
  AND2_X1 U502 ( .A1(G953), .A2(n634), .ZN(n369) );
  XOR2_X1 U503 ( .A(n518), .B(n517), .Z(n370) );
  OR2_X1 U504 ( .A1(n782), .A2(n781), .ZN(n371) );
  NAND2_X1 U505 ( .A1(n766), .A2(n765), .ZN(n450) );
  OR2_X1 U506 ( .A1(n615), .A2(n388), .ZN(n372) );
  AND2_X1 U507 ( .A1(n820), .A2(n737), .ZN(n373) );
  OR2_X1 U508 ( .A1(n769), .A2(KEYINPUT106), .ZN(n374) );
  AND2_X1 U509 ( .A1(n504), .A2(n503), .ZN(n375) );
  AND2_X1 U510 ( .A1(n647), .A2(n438), .ZN(n376) );
  AND2_X1 U511 ( .A1(n463), .A2(n374), .ZN(n377) );
  INV_X1 U512 ( .A(G902), .ZN(n548) );
  OR2_X1 U513 ( .A1(KEYINPUT90), .A2(KEYINPUT47), .ZN(n378) );
  XOR2_X1 U514 ( .A(KEYINPUT67), .B(n698), .Z(n379) );
  INV_X1 U515 ( .A(KEYINPUT91), .ZN(n508) );
  AND2_X1 U516 ( .A1(n697), .A2(n508), .ZN(n380) );
  INV_X1 U517 ( .A(n406), .ZN(n381) );
  XNOR2_X1 U518 ( .A(n811), .B(n382), .ZN(n406) );
  NAND2_X1 U519 ( .A1(n381), .A2(n466), .ZN(n407) );
  XNOR2_X2 U520 ( .A(n381), .B(n547), .ZN(n725) );
  NAND2_X1 U521 ( .A1(n383), .A2(n367), .ZN(n625) );
  NAND2_X1 U522 ( .A1(n383), .A2(n610), .ZN(n611) );
  XNOR2_X2 U523 ( .A(n535), .B(n534), .ZN(n383) );
  XNOR2_X1 U524 ( .A(n546), .B(n384), .ZN(n811) );
  NOR2_X1 U525 ( .A1(n385), .A2(n685), .ZN(n686) );
  NAND2_X1 U526 ( .A1(n385), .A2(n629), .ZN(n612) );
  NOR2_X1 U527 ( .A1(n385), .A2(n438), .ZN(n764) );
  INV_X1 U528 ( .A(n385), .ZN(n387) );
  NAND2_X1 U529 ( .A1(n390), .A2(KEYINPUT66), .ZN(n394) );
  NAND2_X1 U530 ( .A1(n391), .A2(n447), .ZN(n395) );
  NAND2_X1 U531 ( .A1(n393), .A2(n392), .ZN(n445) );
  AND2_X2 U532 ( .A1(n395), .A2(n394), .ZN(n393) );
  XNOR2_X2 U533 ( .A(n398), .B(G146), .ZN(n439) );
  XNOR2_X2 U534 ( .A(G143), .B(G128), .ZN(n593) );
  AND2_X1 U535 ( .A1(n402), .A2(n378), .ZN(n675) );
  XNOR2_X1 U536 ( .A(n402), .B(G143), .ZN(G45) );
  NAND2_X1 U537 ( .A1(n674), .A2(n673), .ZN(n402) );
  OR2_X1 U538 ( .A1(n753), .A2(n496), .ZN(n492) );
  AND2_X1 U539 ( .A1(n671), .A2(n753), .ZN(n467) );
  XNOR2_X1 U540 ( .A(n718), .B(n717), .ZN(n719) );
  BUF_X1 U541 ( .A(n699), .Z(n796) );
  XNOR2_X1 U542 ( .A(n436), .B(n435), .ZN(n434) );
  XNOR2_X1 U543 ( .A(KEYINPUT85), .B(G128), .ZN(n436) );
  XNOR2_X1 U544 ( .A(n434), .B(n432), .ZN(n562) );
  BUF_X1 U545 ( .A(n556), .Z(n403) );
  XNOR2_X2 U546 ( .A(n422), .B(n455), .ZN(n454) );
  XNOR2_X2 U547 ( .A(n452), .B(n803), .ZN(n712) );
  XNOR2_X1 U548 ( .A(n639), .B(KEYINPUT6), .ZN(n405) );
  NAND2_X1 U549 ( .A1(n406), .A2(n557), .ZN(n408) );
  NAND2_X1 U550 ( .A1(n407), .A2(n408), .ZN(n465) );
  BUF_X1 U551 ( .A(n811), .Z(n409) );
  XNOR2_X1 U552 ( .A(n639), .B(KEYINPUT6), .ZN(n451) );
  NAND2_X1 U553 ( .A1(n453), .A2(n478), .ZN(n412) );
  NAND2_X1 U554 ( .A1(n410), .A2(n411), .ZN(n413) );
  NAND2_X1 U555 ( .A1(n412), .A2(n413), .ZN(n452) );
  INV_X1 U556 ( .A(n453), .ZN(n410) );
  INV_X1 U557 ( .A(n478), .ZN(n411) );
  XNOR2_X1 U558 ( .A(n370), .B(n537), .ZN(n478) );
  OR2_X1 U559 ( .A1(n639), .A2(n685), .ZN(n641) );
  XNOR2_X1 U560 ( .A(n659), .B(KEYINPUT19), .ZN(n414) );
  BUF_X1 U561 ( .A(n712), .Z(n415) );
  NAND2_X1 U562 ( .A1(n442), .A2(n604), .ZN(n441) );
  BUF_X1 U563 ( .A(n723), .Z(n791) );
  NAND2_X1 U564 ( .A1(n699), .A2(n508), .ZN(n416) );
  NAND2_X1 U565 ( .A1(n699), .A2(n508), .ZN(n440) );
  NAND2_X1 U566 ( .A1(n695), .A2(KEYINPUT91), .ZN(n418) );
  INV_X1 U567 ( .A(n696), .ZN(n419) );
  NAND2_X1 U568 ( .A1(n475), .A2(n648), .ZN(n421) );
  INV_X1 U569 ( .A(n795), .ZN(n510) );
  XNOR2_X2 U570 ( .A(G902), .B(KEYINPUT15), .ZN(n695) );
  XNOR2_X2 U571 ( .A(n585), .B(n519), .ZN(n422) );
  XNOR2_X1 U572 ( .A(n443), .B(KEYINPUT34), .ZN(n442) );
  NAND2_X1 U573 ( .A1(n647), .A2(n656), .ZN(n425) );
  XNOR2_X2 U574 ( .A(n423), .B(n521), .ZN(n556) );
  XNOR2_X2 U575 ( .A(n520), .B(n522), .ZN(n423) );
  XNOR2_X1 U576 ( .A(n425), .B(n476), .ZN(n475) );
  NAND2_X1 U577 ( .A1(n426), .A2(n635), .ZN(n637) );
  INV_X1 U578 ( .A(G900), .ZN(n427) );
  AND2_X2 U579 ( .A1(n445), .A2(n702), .ZN(n723) );
  INV_X2 U580 ( .A(n429), .ZN(n585) );
  XNOR2_X2 U581 ( .A(G113), .B(G104), .ZN(n429) );
  XNOR2_X2 U582 ( .A(n431), .B(n633), .ZN(n699) );
  NAND2_X1 U583 ( .A1(n497), .A2(n502), .ZN(n431) );
  NAND2_X1 U584 ( .A1(n643), .A2(n745), .ZN(n748) );
  XNOR2_X2 U585 ( .A(n470), .B(KEYINPUT39), .ZN(n643) );
  NAND2_X1 U586 ( .A1(n648), .A2(n438), .ZN(n619) );
  INV_X1 U587 ( .A(n450), .ZN(n438) );
  XNOR2_X1 U588 ( .A(n439), .B(KEYINPUT10), .ZN(n587) );
  NAND2_X1 U589 ( .A1(n447), .A2(n416), .ZN(n444) );
  NOR2_X2 U590 ( .A1(n620), .A2(n750), .ZN(n443) );
  NAND2_X1 U591 ( .A1(n606), .A2(n605), .ZN(n607) );
  INV_X1 U592 ( .A(n405), .ZN(n446) );
  NAND2_X1 U593 ( .A1(n696), .A2(n380), .ZN(n448) );
  INV_X1 U594 ( .A(n699), .ZN(n449) );
  NAND2_X1 U595 ( .A1(n658), .A2(n405), .ZN(n684) );
  NAND2_X1 U596 ( .A1(n712), .A2(n695), .ZN(n525) );
  XNOR2_X2 U597 ( .A(n454), .B(n556), .ZN(n803) );
  AND2_X1 U598 ( .A1(n457), .A2(n374), .ZN(n461) );
  NAND2_X1 U599 ( .A1(n456), .A2(n459), .ZN(n462) );
  NAND2_X1 U600 ( .A1(n622), .A2(n460), .ZN(n459) );
  NAND2_X1 U601 ( .A1(n458), .A2(n623), .ZN(n457) );
  INV_X1 U602 ( .A(n622), .ZN(n458) );
  NAND2_X1 U603 ( .A1(n461), .A2(n459), .ZN(n730) );
  AND2_X1 U604 ( .A1(n769), .A2(KEYINPUT106), .ZN(n460) );
  NAND2_X1 U605 ( .A1(n462), .A2(n664), .ZN(n504) );
  XNOR2_X1 U606 ( .A(n464), .B(G137), .ZN(n545) );
  INV_X1 U607 ( .A(n557), .ZN(n466) );
  NAND2_X1 U608 ( .A1(n670), .A2(n467), .ZN(n470) );
  XNOR2_X2 U609 ( .A(G101), .B(KEYINPUT74), .ZN(n520) );
  NOR2_X1 U610 ( .A1(n787), .A2(G902), .ZN(n602) );
  XNOR2_X1 U611 ( .A(n600), .B(n599), .ZN(n787) );
  NAND2_X1 U612 ( .A1(n709), .A2(n477), .ZN(n653) );
  INV_X1 U613 ( .A(n659), .ZN(n472) );
  NAND2_X1 U614 ( .A1(n681), .A2(n474), .ZN(n683) );
  XNOR2_X1 U615 ( .A(n607), .B(n501), .ZN(n500) );
  XNOR2_X2 U616 ( .A(n550), .B(n549), .ZN(n648) );
  XNOR2_X1 U617 ( .A(n477), .B(G137), .ZN(G39) );
  XNOR2_X1 U618 ( .A(n651), .B(n650), .ZN(n477) );
  NAND2_X1 U619 ( .A1(n487), .A2(n486), .ZN(n485) );
  INV_X1 U620 ( .A(n487), .ZN(n480) );
  AND2_X1 U621 ( .A1(n705), .A2(n693), .ZN(n486) );
  NAND2_X1 U622 ( .A1(n753), .A2(n752), .ZN(n756) );
  NAND2_X1 U623 ( .A1(n491), .A2(n488), .ZN(n776) );
  INV_X1 U624 ( .A(n755), .ZN(n490) );
  NAND2_X1 U625 ( .A1(n494), .A2(n753), .ZN(n493) );
  NOR2_X1 U626 ( .A1(n755), .A2(n495), .ZN(n494) );
  INV_X1 U627 ( .A(n368), .ZN(n496) );
  XNOR2_X2 U628 ( .A(n691), .B(KEYINPUT38), .ZN(n753) );
  XNOR2_X1 U629 ( .A(n499), .B(n498), .ZN(n497) );
  NAND2_X1 U630 ( .A1(n500), .A2(n373), .ZN(n499) );
  INV_X1 U631 ( .A(n606), .ZN(n706) );
  XNOR2_X1 U632 ( .A(n509), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U633 ( .A1(n511), .A2(n510), .ZN(n509) );
  BUF_X1 U634 ( .A(n639), .Z(n769) );
  INV_X1 U635 ( .A(KEYINPUT84), .ZN(n694) );
  XNOR2_X1 U636 ( .A(n404), .B(n584), .ZN(n586) );
  XNOR2_X1 U637 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U638 ( .A(n567), .B(KEYINPUT25), .ZN(n568) );
  XNOR2_X1 U639 ( .A(G475), .B(KEYINPUT13), .ZN(n590) );
  INV_X1 U640 ( .A(KEYINPUT98), .ZN(n513) );
  NAND2_X1 U641 ( .A1(KEYINPUT17), .A2(n513), .ZN(n516) );
  INV_X1 U642 ( .A(KEYINPUT17), .ZN(n514) );
  NAND2_X1 U643 ( .A1(n514), .A2(KEYINPUT98), .ZN(n515) );
  NAND2_X1 U644 ( .A1(n516), .A2(n515), .ZN(n518) );
  XNOR2_X2 U645 ( .A(KEYINPUT80), .B(KEYINPUT16), .ZN(n519) );
  XNOR2_X2 U646 ( .A(KEYINPUT75), .B(KEYINPUT3), .ZN(n522) );
  NAND2_X1 U647 ( .A1(n548), .A2(n523), .ZN(n526) );
  NAND2_X1 U648 ( .A1(n526), .A2(G210), .ZN(n524) );
  AND2_X1 U649 ( .A1(n526), .A2(G214), .ZN(n685) );
  NAND2_X1 U650 ( .A1(G234), .A2(G237), .ZN(n527) );
  NAND2_X1 U651 ( .A1(n530), .A2(G952), .ZN(n528) );
  XNOR2_X1 U652 ( .A(n528), .B(KEYINPUT100), .ZN(n782) );
  INV_X1 U653 ( .A(n782), .ZN(n529) );
  NAND2_X1 U654 ( .A1(n529), .A2(n812), .ZN(n635) );
  NAND2_X1 U655 ( .A1(n530), .A2(G902), .ZN(n531) );
  NOR2_X1 U656 ( .A1(G898), .A2(n812), .ZN(n804) );
  NAND2_X1 U657 ( .A1(n634), .A2(n804), .ZN(n532) );
  NAND2_X1 U658 ( .A1(n635), .A2(n532), .ZN(n533) );
  XNOR2_X1 U659 ( .A(KEYINPUT97), .B(KEYINPUT0), .ZN(n534) );
  INV_X1 U660 ( .A(KEYINPUT102), .ZN(n536) );
  XOR2_X1 U661 ( .A(G140), .B(KEYINPUT71), .Z(n563) );
  XNOR2_X1 U662 ( .A(n537), .B(n563), .ZN(n538) );
  INV_X1 U663 ( .A(n538), .ZN(n540) );
  XNOR2_X2 U664 ( .A(n540), .B(n539), .ZN(n544) );
  NAND2_X1 U665 ( .A1(G227), .A2(n812), .ZN(n542) );
  XNOR2_X2 U666 ( .A(n544), .B(n543), .ZN(n547) );
  XNOR2_X1 U667 ( .A(KEYINPUT70), .B(G131), .ZN(n584) );
  XNOR2_X1 U668 ( .A(n545), .B(n584), .ZN(n546) );
  NAND2_X1 U669 ( .A1(n725), .A2(n548), .ZN(n550) );
  XOR2_X1 U670 ( .A(KEYINPUT73), .B(G469), .Z(n549) );
  NAND2_X1 U671 ( .A1(n577), .A2(G210), .ZN(n552) );
  XNOR2_X1 U672 ( .A(n552), .B(n551), .ZN(n554) );
  XNOR2_X1 U673 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U674 ( .A(n403), .B(n555), .ZN(n557) );
  INV_X1 U675 ( .A(G472), .ZN(n703) );
  XNOR2_X2 U676 ( .A(n558), .B(n703), .ZN(n639) );
  NAND2_X1 U677 ( .A1(n812), .A2(G234), .ZN(n560) );
  XNOR2_X1 U678 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n559) );
  XNOR2_X1 U679 ( .A(n560), .B(n559), .ZN(n596) );
  NAND2_X1 U680 ( .A1(G221), .A2(n596), .ZN(n561) );
  XNOR2_X1 U681 ( .A(n562), .B(n561), .ZN(n564) );
  XNOR2_X1 U682 ( .A(n587), .B(n563), .ZN(n809) );
  XNOR2_X1 U683 ( .A(n564), .B(n809), .ZN(n792) );
  NOR2_X1 U684 ( .A1(n792), .A2(G902), .ZN(n569) );
  NAND2_X1 U685 ( .A1(G234), .A2(n695), .ZN(n565) );
  XNOR2_X1 U686 ( .A(n566), .B(n565), .ZN(n570) );
  NAND2_X1 U687 ( .A1(G217), .A2(n570), .ZN(n567) );
  NAND2_X1 U688 ( .A1(n570), .A2(G221), .ZN(n571) );
  XNOR2_X1 U689 ( .A(n571), .B(KEYINPUT21), .ZN(n572) );
  XOR2_X1 U690 ( .A(KEYINPUT104), .B(n572), .Z(n765) );
  INV_X1 U691 ( .A(KEYINPUT78), .ZN(n574) );
  XOR2_X1 U692 ( .A(n574), .B(KEYINPUT33), .Z(n575) );
  NAND2_X1 U693 ( .A1(G214), .A2(n577), .ZN(n578) );
  XNOR2_X1 U694 ( .A(n579), .B(n578), .ZN(n583) );
  XNOR2_X1 U695 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U696 ( .A(n583), .B(n582), .Z(n589) );
  XNOR2_X1 U697 ( .A(n589), .B(n588), .ZN(n718) );
  XOR2_X1 U698 ( .A(KEYINPUT7), .B(n592), .Z(n595) );
  XOR2_X1 U699 ( .A(n593), .B(G134), .Z(n594) );
  XNOR2_X1 U700 ( .A(n595), .B(n594), .ZN(n600) );
  NAND2_X1 U701 ( .A1(G217), .A2(n596), .ZN(n597) );
  XNOR2_X1 U702 ( .A(n598), .B(n597), .ZN(n599) );
  INV_X1 U703 ( .A(G478), .ZN(n601) );
  XNOR2_X1 U704 ( .A(n602), .B(n601), .ZN(n626) );
  AND2_X1 U705 ( .A1(n628), .A2(n626), .ZN(n673) );
  INV_X1 U706 ( .A(n673), .ZN(n603) );
  XNOR2_X1 U707 ( .A(n603), .B(KEYINPUT87), .ZN(n604) );
  INV_X1 U708 ( .A(KEYINPUT44), .ZN(n605) );
  NOR2_X1 U709 ( .A1(n626), .A2(n628), .ZN(n608) );
  INV_X1 U710 ( .A(n765), .ZN(n609) );
  NOR2_X1 U711 ( .A1(n755), .A2(n609), .ZN(n610) );
  INV_X1 U712 ( .A(n766), .ZN(n629) );
  INV_X1 U713 ( .A(KEYINPUT32), .ZN(n613) );
  XNOR2_X1 U714 ( .A(n614), .B(n613), .ZN(n820) );
  NAND2_X1 U715 ( .A1(n629), .A2(n769), .ZN(n615) );
  OR2_X1 U716 ( .A1(n616), .A2(n372), .ZN(n737) );
  INV_X1 U717 ( .A(n706), .ZN(n617) );
  NAND2_X1 U718 ( .A1(n373), .A2(n617), .ZN(n618) );
  NAND2_X1 U719 ( .A1(n618), .A2(KEYINPUT44), .ZN(n632) );
  OR2_X1 U720 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U721 ( .A(n621), .B(KEYINPUT105), .ZN(n622) );
  INV_X1 U722 ( .A(KEYINPUT106), .ZN(n623) );
  INV_X1 U723 ( .A(n639), .ZN(n647) );
  XOR2_X1 U724 ( .A(KEYINPUT107), .B(KEYINPUT31), .Z(n624) );
  XNOR2_X1 U725 ( .A(n625), .B(n624), .ZN(n746) );
  INV_X1 U726 ( .A(n626), .ZN(n627) );
  NOR2_X1 U727 ( .A1(n628), .A2(n627), .ZN(n745) );
  NOR2_X1 U728 ( .A1(n745), .A2(n655), .ZN(n757) );
  INV_X1 U729 ( .A(n757), .ZN(n664) );
  NOR2_X1 U730 ( .A1(n631), .A2(n630), .ZN(n729) );
  INV_X1 U731 ( .A(KEYINPUT89), .ZN(n636) );
  XNOR2_X1 U732 ( .A(n637), .B(n636), .ZN(n645) );
  AND2_X1 U733 ( .A1(n648), .A2(n638), .ZN(n671) );
  INV_X1 U734 ( .A(KEYINPUT30), .ZN(n640) );
  INV_X1 U735 ( .A(n685), .ZN(n752) );
  NAND2_X1 U736 ( .A1(n645), .A2(n765), .ZN(n646) );
  INV_X1 U737 ( .A(n648), .ZN(n649) );
  INV_X1 U738 ( .A(KEYINPUT42), .ZN(n650) );
  XOR2_X1 U739 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n652) );
  XNOR2_X1 U740 ( .A(n653), .B(n652), .ZN(n681) );
  INV_X1 U741 ( .A(KEYINPUT110), .ZN(n654) );
  XNOR2_X1 U742 ( .A(n655), .B(n654), .ZN(n731) );
  INV_X1 U743 ( .A(n656), .ZN(n657) );
  NOR2_X1 U744 ( .A1(n731), .A2(n657), .ZN(n658) );
  INV_X1 U745 ( .A(KEYINPUT36), .ZN(n660) );
  INV_X1 U746 ( .A(n414), .ZN(n661) );
  INV_X1 U747 ( .A(KEYINPUT90), .ZN(n663) );
  NAND2_X1 U748 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U749 ( .A1(n666), .A2(KEYINPUT47), .ZN(n678) );
  NOR2_X1 U750 ( .A1(n757), .A2(KEYINPUT47), .ZN(n667) );
  XNOR2_X1 U751 ( .A(n667), .B(KEYINPUT81), .ZN(n668) );
  NAND2_X1 U752 ( .A1(n668), .A2(KEYINPUT90), .ZN(n669) );
  NAND2_X1 U753 ( .A1(n741), .A2(n669), .ZN(n676) );
  XNOR2_X1 U754 ( .A(n672), .B(KEYINPUT112), .ZN(n674) );
  AND2_X1 U755 ( .A1(n675), .A2(n676), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n678), .A2(n677), .ZN(n679) );
  INV_X1 U757 ( .A(KEYINPUT48), .ZN(n682) );
  INV_X1 U758 ( .A(n684), .ZN(n687) );
  NAND2_X1 U759 ( .A1(n687), .A2(n686), .ZN(n690) );
  INV_X1 U760 ( .A(KEYINPUT111), .ZN(n688) );
  XNOR2_X1 U761 ( .A(n688), .B(KEYINPUT43), .ZN(n689) );
  XNOR2_X1 U762 ( .A(n690), .B(n689), .ZN(n692) );
  NAND2_X1 U763 ( .A1(n692), .A2(n691), .ZN(n705) );
  INV_X1 U764 ( .A(KEYINPUT94), .ZN(n693) );
  INV_X1 U765 ( .A(n695), .ZN(n697) );
  NAND2_X1 U766 ( .A1(n697), .A2(KEYINPUT2), .ZN(n698) );
  BUF_X1 U767 ( .A(n700), .Z(n701) );
  NAND2_X1 U768 ( .A1(n783), .A2(KEYINPUT2), .ZN(n702) );
  INV_X1 U769 ( .A(G952), .ZN(n704) );
  AND2_X1 U770 ( .A1(n704), .A2(G953), .ZN(n795) );
  XNOR2_X1 U771 ( .A(n705), .B(G140), .ZN(G42) );
  XOR2_X1 U772 ( .A(G122), .B(n706), .Z(G24) );
  XOR2_X1 U773 ( .A(G125), .B(KEYINPUT37), .Z(n707) );
  XNOR2_X1 U774 ( .A(n708), .B(n707), .ZN(G27) );
  XNOR2_X1 U775 ( .A(n709), .B(G131), .ZN(G33) );
  NAND2_X1 U776 ( .A1(n723), .A2(G210), .ZN(n714) );
  XNOR2_X1 U777 ( .A(KEYINPUT96), .B(KEYINPUT54), .ZN(n710) );
  XNOR2_X1 U778 ( .A(n710), .B(KEYINPUT55), .ZN(n711) );
  XNOR2_X1 U779 ( .A(n415), .B(n711), .ZN(n713) );
  XNOR2_X1 U780 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X2 U781 ( .A1(n715), .A2(n795), .ZN(n716) );
  XNOR2_X1 U782 ( .A(n716), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U783 ( .A1(n723), .A2(G475), .ZN(n720) );
  XNOR2_X1 U784 ( .A(KEYINPUT99), .B(KEYINPUT59), .ZN(n717) );
  XNOR2_X1 U785 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X2 U786 ( .A1(n721), .A2(n795), .ZN(n722) );
  XNOR2_X1 U787 ( .A(n722), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U788 ( .A1(n791), .A2(G469), .ZN(n727) );
  XNOR2_X1 U789 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n724) );
  XNOR2_X1 U790 ( .A(n366), .B(n724), .ZN(n726) );
  XNOR2_X1 U791 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U792 ( .A1(n728), .A2(n795), .ZN(G54) );
  XOR2_X1 U793 ( .A(G101), .B(n729), .Z(G3) );
  INV_X1 U794 ( .A(n731), .ZN(n743) );
  NAND2_X1 U795 ( .A1(n730), .A2(n743), .ZN(n732) );
  XNOR2_X1 U796 ( .A(n732), .B(n424), .ZN(G6) );
  XOR2_X1 U797 ( .A(KEYINPUT26), .B(KEYINPUT115), .Z(n734) );
  NAND2_X1 U798 ( .A1(n745), .A2(n730), .ZN(n733) );
  XNOR2_X1 U799 ( .A(n734), .B(n733), .ZN(n736) );
  XOR2_X1 U800 ( .A(G107), .B(KEYINPUT27), .Z(n735) );
  XNOR2_X1 U801 ( .A(n736), .B(n735), .ZN(G9) );
  XNOR2_X1 U802 ( .A(G110), .B(n737), .ZN(G12) );
  XOR2_X1 U803 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n739) );
  NAND2_X1 U804 ( .A1(n745), .A2(n741), .ZN(n738) );
  XNOR2_X1 U805 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U806 ( .A(G128), .B(n740), .ZN(G30) );
  NAND2_X1 U807 ( .A1(n741), .A2(n743), .ZN(n742) );
  XNOR2_X1 U808 ( .A(n742), .B(G146), .ZN(G48) );
  NAND2_X1 U809 ( .A1(n743), .A2(n746), .ZN(n744) );
  XNOR2_X1 U810 ( .A(n744), .B(n430), .ZN(G15) );
  NAND2_X1 U811 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U812 ( .A(n747), .B(G116), .ZN(G18) );
  XOR2_X1 U813 ( .A(G134), .B(n748), .Z(n749) );
  XNOR2_X1 U814 ( .A(n749), .B(KEYINPUT117), .ZN(G36) );
  BUF_X1 U815 ( .A(n750), .Z(n762) );
  NOR2_X1 U816 ( .A1(n762), .A2(n776), .ZN(n751) );
  NOR2_X1 U817 ( .A1(G953), .A2(n751), .ZN(n785) );
  NOR2_X1 U818 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U819 ( .A1(n755), .A2(n754), .ZN(n759) );
  NOR2_X1 U820 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U821 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U822 ( .A(KEYINPUT119), .B(n760), .Z(n761) );
  NOR2_X1 U823 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U824 ( .A(n763), .B(KEYINPUT120), .ZN(n778) );
  XNOR2_X1 U825 ( .A(n764), .B(KEYINPUT50), .ZN(n772) );
  NOR2_X1 U826 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U827 ( .A(n767), .B(KEYINPUT49), .ZN(n768) );
  XNOR2_X1 U828 ( .A(n768), .B(KEYINPUT118), .ZN(n770) );
  NAND2_X1 U829 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U830 ( .A1(n772), .A2(n771), .ZN(n773) );
  OR2_X1 U831 ( .A1(n773), .A2(n367), .ZN(n774) );
  XNOR2_X1 U832 ( .A(KEYINPUT51), .B(n774), .ZN(n775) );
  NOR2_X1 U833 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U834 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U835 ( .A(n779), .B(KEYINPUT121), .Z(n780) );
  XNOR2_X1 U836 ( .A(KEYINPUT52), .B(n780), .ZN(n781) );
  NAND2_X1 U837 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U838 ( .A(KEYINPUT53), .B(n786), .Z(G75) );
  NAND2_X1 U839 ( .A1(n791), .A2(G478), .ZN(n789) );
  XNOR2_X1 U840 ( .A(n787), .B(KEYINPUT122), .ZN(n788) );
  XNOR2_X1 U841 ( .A(n789), .B(n788), .ZN(n790) );
  NOR2_X1 U842 ( .A1(n795), .A2(n790), .ZN(G63) );
  NAND2_X1 U843 ( .A1(n791), .A2(G217), .ZN(n793) );
  XNOR2_X1 U844 ( .A(n793), .B(n792), .ZN(n794) );
  NOR2_X1 U845 ( .A1(n795), .A2(n794), .ZN(G66) );
  INV_X1 U846 ( .A(n796), .ZN(n797) );
  NAND2_X1 U847 ( .A1(n797), .A2(n812), .ZN(n802) );
  NAND2_X1 U848 ( .A1(G953), .A2(G224), .ZN(n798) );
  XNOR2_X1 U849 ( .A(KEYINPUT61), .B(n798), .ZN(n799) );
  NAND2_X1 U850 ( .A1(n799), .A2(G898), .ZN(n800) );
  XOR2_X1 U851 ( .A(KEYINPUT123), .B(n800), .Z(n801) );
  NAND2_X1 U852 ( .A1(n802), .A2(n801), .ZN(n807) );
  XNOR2_X1 U853 ( .A(n803), .B(G110), .ZN(n805) );
  NOR2_X1 U854 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U855 ( .A(n807), .B(n806), .ZN(G69) );
  XOR2_X1 U856 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n808) );
  XNOR2_X1 U857 ( .A(n809), .B(n808), .ZN(n810) );
  XOR2_X1 U858 ( .A(n409), .B(n810), .Z(n814) );
  XNOR2_X1 U859 ( .A(n701), .B(n814), .ZN(n813) );
  NAND2_X1 U860 ( .A1(n813), .A2(n812), .ZN(n819) );
  XNOR2_X1 U861 ( .A(G227), .B(n814), .ZN(n815) );
  NAND2_X1 U862 ( .A1(n815), .A2(G900), .ZN(n816) );
  XNOR2_X1 U863 ( .A(KEYINPUT126), .B(n816), .ZN(n817) );
  NAND2_X1 U864 ( .A1(n817), .A2(G953), .ZN(n818) );
  NAND2_X1 U865 ( .A1(n819), .A2(n818), .ZN(G72) );
  XOR2_X1 U866 ( .A(G119), .B(n820), .Z(n821) );
  XNOR2_X1 U867 ( .A(KEYINPUT127), .B(n821), .ZN(G21) );
endmodule

