//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950;
  XNOR2_X1  g000(.A(KEYINPUT72), .B(G197gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G204gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n203), .B(new_n204), .C1(KEYINPUT22), .C2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(KEYINPUT73), .ZN(new_n210));
  XOR2_X1   g009(.A(new_n208), .B(new_n210), .Z(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G141gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT75), .B(G141gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(new_n212), .ZN(new_n215));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n219), .B2(KEYINPUT2), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G141gat), .B(G148gat), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n216), .B(new_n219), .C1(new_n222), .C2(KEYINPUT2), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(KEYINPUT74), .B(KEYINPUT29), .Z(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n211), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(new_n223), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n208), .B(new_n210), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n225), .B1(new_n231), .B2(new_n227), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n229), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n233), .B1(G228gat), .B2(G233gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(G228gat), .A2(G233gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n225), .B1(new_n231), .B2(KEYINPUT29), .ZN(new_n236));
  AOI211_X1 g035(.A(new_n235), .B(new_n229), .C1(new_n230), .C2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G78gat), .B(G106gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT31), .B(G50gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(G22gat), .ZN(new_n242));
  INV_X1    g041(.A(G22gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(KEYINPUT77), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n242), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n238), .B(new_n245), .Z(new_n246));
  XNOR2_X1  g045(.A(G1gat), .B(G29gat), .ZN(new_n247));
  INV_X1    g046(.A(G85gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT0), .B(G57gat), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n249), .B(new_n250), .Z(new_n251));
  XNOR2_X1  g050(.A(G127gat), .B(G134gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(KEYINPUT68), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n230), .A2(KEYINPUT3), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n226), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G225gat), .A2(G233gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT76), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n256), .A2(new_n224), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n256), .B2(new_n224), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n259), .B(new_n262), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT5), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n257), .A2(new_n230), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n256), .A2(new_n224), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n261), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n251), .B(new_n269), .C1(new_n274), .C2(new_n268), .ZN(new_n275));
  INV_X1    g074(.A(new_n251), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n268), .B1(new_n267), .B2(new_n273), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n271), .A2(KEYINPUT4), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n256), .B1(KEYINPUT3), .B2(new_n230), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n278), .A2(new_n264), .B1(new_n279), .B2(new_n226), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT5), .B1(new_n280), .B2(new_n262), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n276), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n275), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n277), .A2(new_n281), .A3(new_n276), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT6), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT27), .B(G183gat), .ZN(new_n289));
  INV_X1    g088(.A(G190gat), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT66), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n291), .A2(KEYINPUT28), .ZN(new_n292));
  NOR2_X1   g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n295));
  OR3_X1    g094(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT26), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(KEYINPUT26), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(new_n294), .B2(KEYINPUT26), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n291), .A2(KEYINPUT28), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n292), .A2(new_n300), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT64), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n307));
  INV_X1    g106(.A(G183gat), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(new_n290), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT65), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n294), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n294), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT65), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n306), .A2(new_n316), .A3(new_n309), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n311), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT25), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n309), .A2(new_n304), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n315), .A2(KEYINPUT25), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n303), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n322), .B1(new_n318), .B2(new_n319), .ZN(new_n327));
  INV_X1    g126(.A(new_n303), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(new_n227), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n326), .B(new_n231), .C1(new_n330), .C2(new_n325), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n324), .B1(new_n329), .B2(KEYINPUT29), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n332), .A2(new_n326), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n333), .B2(new_n231), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n335));
  XNOR2_X1  g134(.A(G8gat), .B(G36gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(G64gat), .B(G92gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n334), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n334), .A2(new_n339), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n331), .B(new_n338), .C1(new_n333), .C2(new_n231), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(KEYINPUT30), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n288), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n246), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT36), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n257), .ZN(new_n347));
  INV_X1    g146(.A(G227gat), .ZN(new_n348));
  INV_X1    g147(.A(G233gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n256), .B1(new_n327), .B2(new_n328), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G71gat), .B(G99gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(G43gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT70), .B(G15gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  XOR2_X1   g155(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(KEYINPUT32), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT71), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n352), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n363), .B2(new_n356), .ZN(new_n364));
  INV_X1    g163(.A(new_n356), .ZN(new_n365));
  AOI211_X1 g164(.A(KEYINPUT71), .B(new_n365), .C1(new_n352), .C2(new_n362), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n359), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT34), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n347), .A2(new_n351), .ZN(new_n369));
  INV_X1    g168(.A(new_n350), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT34), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n373), .B(new_n359), .C1(new_n364), .C2(new_n366), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n368), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n372), .B1(new_n368), .B2(new_n374), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n346), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n368), .A2(new_n374), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n371), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n368), .A2(new_n372), .A3(new_n374), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(KEYINPUT36), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n345), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n332), .A2(new_n326), .A3(new_n231), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n329), .A2(new_n324), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n323), .A2(new_n228), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n386), .B2(new_n324), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n384), .B(KEYINPUT37), .C1(new_n387), .C2(new_n231), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT37), .ZN(new_n391));
  INV_X1    g190(.A(new_n331), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n231), .B1(new_n332), .B2(new_n326), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n326), .B1(new_n330), .B2(new_n325), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n211), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n396), .A2(KEYINPUT78), .A3(KEYINPUT37), .A4(new_n384), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n390), .A2(new_n338), .A3(new_n394), .A4(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT38), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n339), .B1(new_n334), .B2(new_n391), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n392), .A2(new_n393), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n401), .B2(KEYINPUT37), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n398), .A2(new_n399), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n286), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n288), .B2(new_n404), .ZN(new_n406));
  INV_X1    g205(.A(new_n341), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n403), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n280), .A2(new_n262), .ZN(new_n409));
  OR2_X1    g208(.A1(new_n409), .A2(KEYINPUT39), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n409), .B(KEYINPUT39), .C1(new_n261), .C2(new_n272), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n276), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT40), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n343), .A2(new_n275), .A3(new_n340), .A4(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n412), .A2(new_n413), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n246), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n383), .B1(new_n408), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n405), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n419), .B1(new_n287), .B2(KEYINPUT79), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n398), .A2(new_n399), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n402), .A2(new_n400), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n341), .B(new_n420), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n415), .A2(new_n416), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n423), .A2(KEYINPUT80), .A3(new_n246), .A4(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n382), .A2(new_n418), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n238), .B(new_n245), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n375), .A2(new_n376), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT35), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n343), .A2(new_n340), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .A4(new_n406), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n379), .A2(new_n344), .A3(new_n246), .A4(new_n380), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT35), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n436));
  INV_X1    g235(.A(G29gat), .ZN(new_n437));
  INV_X1    g236(.A(G36gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G29gat), .A2(G36gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(G43gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(G50gat), .ZN(new_n445));
  INV_X1    g244(.A(G50gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(G43gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n447), .A3(KEYINPUT15), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n443), .A2(new_n449), .A3(KEYINPUT81), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT81), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n439), .A2(new_n440), .B1(G29gat), .B2(G36gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(new_n448), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n447), .ZN(new_n455));
  AND2_X1   g254(.A1(KEYINPUT83), .A2(G50gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(KEYINPUT83), .A2(G50gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n458), .B2(new_n444), .ZN(new_n459));
  XOR2_X1   g258(.A(KEYINPUT82), .B(KEYINPUT15), .Z(new_n460));
  OAI211_X1 g259(.A(new_n452), .B(new_n448), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n454), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT17), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n454), .A2(KEYINPUT17), .A3(new_n461), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT93), .ZN(new_n466));
  NAND2_X1  g265(.A1(G99gat), .A2(G106gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(G99gat), .A2(G106gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT92), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G99gat), .ZN(new_n472));
  INV_X1    g271(.A(G106gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT92), .B1(new_n474), .B2(new_n467), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n466), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n470), .B1(new_n468), .B2(new_n469), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(KEYINPUT92), .A3(new_n467), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT93), .ZN(new_n479));
  INV_X1    g278(.A(G92gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n248), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n467), .A2(KEYINPUT8), .ZN(new_n482));
  NAND2_X1  g281(.A1(G85gat), .A2(G92gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT7), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n486));
  AND4_X1   g285(.A1(new_n481), .A2(new_n482), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n476), .A2(new_n479), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n477), .A2(new_n478), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n482), .A2(new_n485), .A3(new_n481), .A4(new_n486), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n466), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n464), .A2(new_n465), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(G232gat), .A2(G233gat), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n462), .A2(new_n492), .B1(KEYINPUT41), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n494), .A2(new_n290), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n290), .B1(new_n494), .B2(new_n496), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n206), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n494), .A2(new_n496), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G190gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n494), .A2(new_n290), .A3(new_n496), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(G218gat), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(new_n503), .A3(KEYINPUT91), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n495), .A2(KEYINPUT41), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(KEYINPUT90), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n506), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n499), .A2(new_n503), .A3(KEYINPUT91), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G134gat), .B(G162gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(new_n511), .A3(new_n509), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G64gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G57gat), .ZN(new_n517));
  INV_X1    g316(.A(G57gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G64gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT89), .ZN(new_n521));
  NAND2_X1  g320(.A1(G71gat), .A2(G78gat), .ZN(new_n522));
  OR2_X1    g321(.A1(G71gat), .A2(G78gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT9), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n517), .A2(new_n519), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n521), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AND3_X1   g327(.A1(KEYINPUT88), .A2(G71gat), .A3(G78gat), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT88), .B1(G71gat), .B2(G78gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(G57gat), .B(G64gat), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n531), .B(new_n523), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT21), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(new_n205), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n540));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541));
  INV_X1    g340(.A(G1gat), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n542), .A2(KEYINPUT84), .A3(KEYINPUT16), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT84), .B1(new_n542), .B2(KEYINPUT16), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT85), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  OR3_X1    g346(.A1(new_n541), .A2(KEYINPUT86), .A3(G1gat), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(G8gat), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G8gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT84), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT16), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(G1gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n542), .A2(KEYINPUT84), .A3(KEYINPUT16), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT87), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(new_n541), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n556), .B2(new_n541), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n551), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n541), .A2(G1gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n551), .A2(KEYINPUT86), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n561), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n550), .B(new_n566), .C1(new_n536), .C2(new_n535), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n567), .A2(G183gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(G183gat), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n540), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n569), .A3(new_n540), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n539), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G127gat), .B(G155gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(new_n572), .A3(new_n539), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n577), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n571), .A2(new_n572), .A3(new_n539), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(new_n573), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n515), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n515), .A2(new_n583), .A3(KEYINPUT94), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n464), .A2(new_n550), .A3(new_n566), .A4(new_n465), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n545), .A2(KEYINPUT87), .ZN(new_n590));
  AOI21_X1  g389(.A(G8gat), .B1(new_n590), .B2(new_n558), .ZN(new_n591));
  NOR3_X1   g390(.A1(new_n591), .A2(new_n562), .A3(new_n564), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n545), .A2(new_n546), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT85), .B1(new_n556), .B2(new_n541), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n551), .B1(new_n595), .B2(new_n548), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n462), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n589), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT18), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n550), .A2(new_n566), .A3(new_n454), .A4(new_n461), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n598), .B(KEYINPUT13), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n589), .A2(new_n597), .A3(KEYINPUT18), .A4(new_n598), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n601), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609));
  INV_X1    g408(.A(G197gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT11), .B(G169gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n601), .A2(new_n606), .A3(new_n607), .A4(new_n614), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n488), .A2(new_n535), .A3(new_n491), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n489), .B1(new_n487), .B2(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n490), .A2(KEYINPUT95), .A3(new_n477), .A4(new_n478), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n621), .A2(new_n534), .A3(new_n528), .A4(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT96), .B(KEYINPUT10), .Z(new_n624));
  NAND3_X1  g423(.A1(new_n619), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n535), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n492), .A2(KEYINPUT10), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n619), .A2(new_n623), .ZN(new_n631));
  INV_X1    g430(.A(new_n629), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT97), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n635), .A3(new_n632), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n630), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT98), .B(G176gat), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G204gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n637), .B(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n588), .A2(new_n618), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n435), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n287), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(new_n542), .ZN(G1324gat));
  NOR2_X1   g446(.A1(new_n645), .A2(new_n430), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT16), .B(G8gat), .Z(new_n649));
  AND2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n650), .A2(KEYINPUT42), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(KEYINPUT42), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n651), .B(new_n652), .C1(new_n551), .C2(new_n648), .ZN(G1325gat));
  INV_X1    g452(.A(G15gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n377), .A2(new_n381), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n645), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n645), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n375), .A2(new_n376), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n656), .B1(new_n654), .B2(new_n659), .ZN(G1326gat));
  INV_X1    g459(.A(KEYINPUT99), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n661), .B1(new_n657), .B2(new_n427), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n645), .A2(KEYINPUT99), .A3(new_n246), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT43), .B(G22gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  INV_X1    g465(.A(new_n515), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n435), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n583), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n618), .A2(new_n643), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n437), .A3(new_n288), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n515), .A2(KEYINPUT44), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n435), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n426), .A2(new_n434), .A3(KEYINPUT100), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n435), .B2(new_n667), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n683), .A2(new_n287), .A3(new_n671), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n674), .B1(new_n684), .B2(new_n437), .ZN(G1328gat));
  INV_X1    g484(.A(new_n430), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n672), .A2(new_n438), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n683), .A2(new_n430), .A3(new_n671), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n689), .B(KEYINPUT101), .C1(new_n690), .C2(new_n438), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n687), .B(KEYINPUT46), .ZN(new_n693));
  INV_X1    g492(.A(new_n679), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT100), .B1(new_n426), .B2(new_n434), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n675), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n682), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n671), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n438), .B1(new_n698), .B2(new_n686), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n692), .B1(new_n693), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n691), .A2(new_n700), .ZN(G1329gat));
  INV_X1    g500(.A(new_n655), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n698), .A2(KEYINPUT103), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n671), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n702), .B(new_n704), .C1(new_n680), .C2(new_n682), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n703), .A2(new_n707), .A3(G43gat), .ZN(new_n708));
  INV_X1    g507(.A(new_n658), .ZN(new_n709));
  NOR4_X1   g508(.A1(new_n668), .A2(G43gat), .A3(new_n709), .A4(new_n671), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n708), .A2(KEYINPUT47), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n444), .B1(new_n698), .B2(new_n702), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(new_n710), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(G1330gat));
  INV_X1    g515(.A(new_n458), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n427), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT104), .Z(new_n719));
  NAND2_X1  g518(.A1(new_n672), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n683), .A2(new_n246), .A3(new_n671), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n721), .B2(new_n717), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(KEYINPUT48), .B(new_n720), .C1(new_n721), .C2(new_n717), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1331gat));
  NAND2_X1  g525(.A1(new_n678), .A2(new_n679), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n616), .A2(new_n617), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n588), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n727), .A2(new_n643), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n287), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT105), .B(G57gat), .Z(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1332gat));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n430), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  AND2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n734), .B2(new_n735), .ZN(G1333gat));
  INV_X1    g537(.A(new_n730), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G71gat), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n730), .A2(new_n709), .ZN(new_n741));
  OAI22_X1  g540(.A1(new_n740), .A2(new_n655), .B1(new_n741), .B2(G71gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g542(.A1(new_n730), .A2(new_n246), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT106), .B(G78gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n583), .A2(new_n728), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT51), .B1(new_n668), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n435), .A2(new_n750), .A3(new_n667), .A4(new_n747), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n749), .A2(new_n643), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n288), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n747), .A2(new_n643), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT107), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n696), .B2(new_n697), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(new_n248), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n753), .B1(new_n759), .B2(new_n288), .ZN(G1336gat));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n686), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT108), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n763), .A2(KEYINPUT108), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n752), .A2(new_n480), .A3(new_n686), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n762), .A2(new_n764), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n480), .B1(new_n757), .B2(new_n686), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n749), .A2(new_n480), .A3(new_n643), .A4(new_n751), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n430), .ZN(new_n770));
  OAI211_X1 g569(.A(KEYINPUT108), .B(new_n763), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n767), .A2(new_n771), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n758), .B2(new_n655), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n752), .A2(new_n472), .A3(new_n658), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(G1338gat));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n757), .A2(new_n776), .A3(new_n427), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n427), .B(new_n755), .C1(new_n680), .C2(new_n682), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT110), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n779), .A3(G106gat), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n246), .A2(G106gat), .ZN(new_n781));
  AND4_X1   g580(.A1(new_n643), .A2(new_n749), .A3(new_n751), .A4(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(KEYINPUT53), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n778), .A2(KEYINPUT109), .A3(G106gat), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT109), .B1(new_n778), .B2(G106gat), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n785), .A2(new_n786), .A3(new_n782), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n603), .B2(new_n605), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n597), .A2(new_n602), .A3(KEYINPUT112), .A4(new_n604), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n589), .A2(new_n597), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n791), .B(new_n792), .C1(new_n793), .C2(new_n598), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n613), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n643), .A3(new_n617), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n625), .A2(new_n632), .A3(new_n627), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n625), .A2(new_n627), .A3(KEYINPUT111), .A4(new_n632), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n799), .A2(new_n630), .A3(KEYINPUT54), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n632), .B1(new_n625), .B2(new_n627), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n641), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n637), .A2(new_n642), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n801), .A2(KEYINPUT55), .A3(new_n804), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n796), .B1(new_n618), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n796), .B(KEYINPUT113), .C1(new_n618), .C2(new_n810), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n515), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n795), .A2(new_n617), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n810), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n513), .A2(new_n817), .A3(new_n514), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n815), .A2(KEYINPUT114), .A3(new_n818), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n669), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n643), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n586), .A2(new_n618), .A3(new_n824), .A4(new_n587), .ZN(new_n825));
  AOI211_X1 g624(.A(new_n709), .B(new_n427), .C1(new_n823), .C2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n686), .A2(new_n287), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n728), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n643), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g631(.A1(new_n828), .A2(new_n583), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(G127gat), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n833), .B(new_n835), .Z(G1342gat));
  NAND2_X1  g635(.A1(new_n828), .A2(new_n667), .ZN(new_n837));
  OR3_X1    g636(.A1(new_n837), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(G134gat), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT56), .B1(new_n837), .B2(G134gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(G1343gat));
  AND3_X1   g640(.A1(new_n815), .A2(KEYINPUT114), .A3(new_n818), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT114), .B1(new_n815), .B2(new_n818), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n842), .A2(new_n843), .A3(new_n583), .ZN(new_n844));
  INV_X1    g643(.A(new_n825), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n427), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(KEYINPUT116), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n246), .B1(new_n823), .B2(new_n825), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(KEYINPUT57), .ZN(new_n851));
  NOR2_X1   g650(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n805), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n805), .A2(new_n852), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n728), .A2(new_n853), .A3(new_n808), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n796), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT118), .B1(new_n515), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n515), .A2(KEYINPUT118), .A3(new_n856), .ZN(new_n858));
  AOI211_X1 g657(.A(new_n857), .B(new_n858), .C1(new_n667), .C2(new_n817), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n825), .B1(new_n859), .B2(new_n583), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(KEYINPUT57), .A3(new_n427), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n848), .A2(new_n851), .A3(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n655), .A2(new_n827), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n728), .A3(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n862), .A2(KEYINPUT121), .A3(new_n728), .A4(new_n863), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n214), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n846), .A2(new_n702), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n827), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(G141gat), .A3(new_n618), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  XOR2_X1   g671(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n873));
  NAND3_X1  g672(.A1(new_n868), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n864), .A2(new_n875), .A3(new_n214), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n864), .B2(new_n214), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n877), .A3(new_n871), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n874), .B1(new_n878), .B2(new_n879), .ZN(G1344gat));
  INV_X1    g679(.A(new_n870), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n212), .A3(new_n643), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n825), .B(KEYINPUT122), .Z(new_n884));
  NAND2_X1  g683(.A1(new_n515), .A2(new_n856), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n583), .B1(new_n885), .B2(new_n818), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n847), .B(new_n427), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n846), .A2(KEYINPUT57), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n887), .A2(new_n643), .A3(new_n863), .A4(new_n888), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n889), .A2(KEYINPUT123), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n212), .B1(new_n889), .B2(KEYINPUT123), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n883), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n862), .A2(new_n863), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT59), .B(new_n212), .C1(new_n893), .C2(new_n643), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n882), .B1(new_n892), .B2(new_n894), .ZN(G1345gat));
  AOI21_X1  g694(.A(G155gat), .B1(new_n881), .B2(new_n583), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n669), .A2(new_n217), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n893), .B2(new_n897), .ZN(G1346gat));
  NAND3_X1  g697(.A1(new_n893), .A2(G162gat), .A3(new_n667), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n218), .B1(new_n870), .B2(new_n515), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT124), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n899), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1347gat));
  NOR2_X1   g704(.A1(new_n430), .A2(new_n288), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n826), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(G169gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n908), .A3(new_n728), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n906), .B(KEYINPUT125), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n826), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G169gat), .B1(new_n911), .B2(new_n618), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n912), .ZN(G1348gat));
  AOI21_X1  g712(.A(G176gat), .B1(new_n907), .B2(new_n643), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n911), .A2(new_n824), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(G176gat), .B2(new_n915), .ZN(G1349gat));
  INV_X1    g715(.A(new_n911), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n308), .B1(new_n917), .B2(new_n583), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n583), .A2(new_n289), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n907), .B2(new_n919), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT60), .Z(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n911), .B2(new_n515), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT61), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n290), .A3(new_n667), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1351gat));
  NAND4_X1  g724(.A1(new_n887), .A2(new_n655), .A3(new_n888), .A4(new_n910), .ZN(new_n926));
  OAI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n618), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n869), .A2(new_n906), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n610), .A3(new_n728), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n931), .B(new_n932), .ZN(G1352gat));
  NOR3_X1   g732(.A1(new_n928), .A2(G204gat), .A3(new_n824), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT62), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n887), .A2(new_n643), .A3(new_n888), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n655), .A2(new_n910), .ZN(new_n937));
  OAI21_X1  g736(.A(G204gat), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n938), .ZN(G1353gat));
  OAI21_X1  g738(.A(G211gat), .B1(new_n926), .B2(new_n669), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g741(.A(KEYINPUT63), .B(G211gat), .C1(new_n926), .C2(new_n669), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(KEYINPUT127), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n205), .A3(new_n583), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n940), .A2(new_n946), .A3(new_n941), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(G1354gat));
  OAI21_X1  g747(.A(G218gat), .B1(new_n926), .B2(new_n515), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n929), .A2(new_n206), .A3(new_n667), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1355gat));
endmodule


