//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  OAI211_X1 g006(.A(G128), .B(new_n189), .C1(new_n190), .C2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n194), .B(new_n195), .C1(KEYINPUT1), .C2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n193), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G137), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT11), .A3(G134), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(G137), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n201), .A2(new_n203), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(G134), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n205), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT65), .B1(new_n208), .B2(G131), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n210));
  AOI211_X1 g024(.A(new_n210), .B(new_n204), .C1(new_n207), .C2(new_n205), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n198), .B(new_n206), .C1(new_n209), .C2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n213));
  INV_X1    g027(.A(G113), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT67), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT2), .A3(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n214), .ZN(new_n219));
  INV_X1    g033(.A(G119), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G116), .ZN(new_n221));
  INV_X1    g035(.A(G116), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G119), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n218), .A2(new_n219), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n221), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(new_n221), .B2(new_n223), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n215), .A2(new_n217), .B1(new_n213), .B2(new_n214), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n224), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G143), .B(G146), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(KEYINPUT0), .B2(G128), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n233), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT0), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT64), .B1(new_n238), .B2(new_n196), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n239), .B(new_n232), .C1(new_n190), .C2(new_n192), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G131), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n206), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n212), .A2(new_n231), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT69), .B(G953), .ZN(new_n248));
  INV_X1    g062(.A(G237), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(G210), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n212), .B2(new_n246), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n241), .B1(new_n244), .B2(new_n206), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n193), .A2(new_n197), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n206), .B1(new_n209), .B2(new_n211), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI211_X1 g075(.A(KEYINPUT66), .B(new_n206), .C1(new_n209), .C2(new_n211), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n256), .B1(new_n263), .B2(new_n255), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n247), .B(new_n254), .C1(new_n264), .C2(new_n231), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT31), .B1(new_n265), .B2(KEYINPUT71), .ZN(new_n266));
  INV_X1    g080(.A(new_n247), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n200), .A2(G137), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n202), .A2(G134), .ZN(new_n269));
  OAI21_X1  g083(.A(G131), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n210), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n208), .A2(KEYINPUT65), .A3(G131), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n271), .A2(new_n272), .B1(new_n204), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n198), .B1(new_n274), .B2(KEYINPUT66), .ZN(new_n275));
  INV_X1    g089(.A(new_n262), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n255), .B(new_n246), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n256), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n267), .B1(new_n279), .B2(new_n230), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT31), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .A4(new_n254), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n266), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n246), .B1(new_n275), .B2(new_n276), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n230), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT73), .B1(new_n263), .B2(new_n231), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n288), .A3(new_n247), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n247), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n254), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n187), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT32), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n231), .B1(new_n246), .B2(new_n212), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT28), .B1(new_n267), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n293), .A3(new_n254), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT29), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n254), .B2(new_n280), .ZN(new_n303));
  INV_X1    g117(.A(new_n293), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n254), .A2(new_n305), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n304), .B(new_n306), .C1(new_n289), .C2(new_n290), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n298), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G472), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n304), .B1(new_n289), .B2(new_n290), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n266), .B(new_n283), .C1(new_n310), .C2(new_n254), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT32), .A3(new_n187), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n297), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n297), .A2(new_n309), .A3(KEYINPUT74), .A4(new_n312), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT81), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT22), .B(G137), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT79), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n248), .A2(G221), .A3(G234), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n320), .B(new_n321), .Z(new_n322));
  XNOR2_X1  g136(.A(G119), .B(G128), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT75), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT24), .B(G110), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(KEYINPUT76), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT23), .B1(new_n196), .B2(G119), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n220), .B2(G128), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n327), .B1(G110), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G125), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT78), .ZN(new_n340));
  XNOR2_X1  g154(.A(G125), .B(G140), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(G146), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT16), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(new_n335), .A3(G125), .ZN(new_n346));
  OAI211_X1 g160(.A(G146), .B(new_n346), .C1(new_n339), .C2(new_n345), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n334), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n333), .A2(G110), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n346), .B1(new_n339), .B2(new_n345), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n191), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n347), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n351), .B(new_n354), .C1(new_n324), .C2(new_n326), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n322), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n350), .A2(KEYINPUT80), .A3(new_n355), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n356), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT80), .A3(new_n322), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G217), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(G234), .B2(new_n298), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n318), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(KEYINPUT81), .B(new_n367), .C1(new_n360), .C2(new_n363), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n358), .A2(new_n359), .ZN(new_n372));
  AOI21_X1  g186(.A(G902), .B1(new_n372), .B2(new_n362), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n366), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI211_X1 g189(.A(KEYINPUT25), .B(G902), .C1(new_n372), .C2(new_n362), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n371), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT82), .B1(new_n317), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n377), .A2(new_n371), .ZN(new_n381));
  AOI211_X1 g195(.A(new_n380), .B(new_n381), .C1(new_n315), .C2(new_n316), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G104), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  INV_X1    g201(.A(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(KEYINPUT3), .A3(G104), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G101), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n384), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n388), .A2(G107), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n385), .A2(KEYINPUT3), .A3(G104), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT3), .B1(new_n385), .B2(G104), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G101), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n384), .A3(G101), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n230), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G122), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n385), .A2(G104), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n392), .B1(new_n394), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n391), .B2(new_n392), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT5), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n226), .A2(new_n227), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n222), .A2(G119), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n214), .B1(new_n408), .B2(new_n406), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n224), .B(new_n405), .C1(new_n407), .C2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n401), .A2(new_n402), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT86), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT86), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n401), .A2(new_n411), .A3(new_n414), .A4(new_n402), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(KEYINPUT6), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n402), .B1(new_n401), .B2(new_n411), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT85), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT6), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n419), .A3(KEYINPUT6), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n416), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n337), .B1(new_n237), .B2(new_n240), .ZN(new_n424));
  AOI21_X1  g238(.A(G125), .B1(new_n193), .B2(new_n197), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT87), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n425), .A2(KEYINPUT87), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G224), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(G953), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT88), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n428), .B(new_n431), .Z(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n423), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G210), .B1(G237), .B2(G902), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n413), .A2(new_n415), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT7), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n426), .A2(new_n427), .A3(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n392), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n394), .A2(new_n403), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G101), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n224), .B(new_n443), .C1(new_n407), .C2(new_n410), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n221), .A2(new_n223), .A3(KEYINPUT5), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n409), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n224), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n405), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n402), .B(KEYINPUT8), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n439), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n438), .B1(new_n426), .B2(new_n427), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n436), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n434), .A2(new_n298), .A3(new_n435), .A4(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n435), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n417), .B(new_n420), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n432), .B1(new_n457), .B2(new_n416), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n298), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G214), .B1(G237), .B2(G902), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT89), .ZN(new_n464));
  INV_X1    g278(.A(G469), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n399), .A2(new_n242), .A3(new_n400), .ZN(new_n466));
  INV_X1    g280(.A(new_n245), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n440), .A2(new_n197), .A3(new_n193), .A4(new_n442), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT10), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n198), .A2(KEYINPUT10), .A3(new_n405), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n466), .A2(new_n467), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT83), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n468), .B(KEYINPUT10), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n475), .A2(KEYINPUT83), .A3(new_n467), .A4(new_n466), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n248), .A2(G227), .ZN(new_n478));
  XNOR2_X1  g292(.A(G110), .B(G140), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n443), .A2(new_n258), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n467), .B1(new_n481), .B2(new_n468), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT12), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n477), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n399), .A2(new_n242), .A3(new_n400), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n471), .A2(new_n470), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT84), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT84), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n466), .A2(new_n488), .A3(new_n470), .A4(new_n471), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n245), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n480), .B1(new_n477), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n465), .B(new_n298), .C1(new_n484), .C2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n465), .A2(new_n298), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n477), .A2(new_n490), .A3(new_n480), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n477), .A2(new_n483), .ZN(new_n496));
  OAI211_X1 g310(.A(G469), .B(new_n495), .C1(new_n496), .C2(new_n480), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n492), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G221), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT9), .B(G234), .Z(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(new_n298), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n464), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT93), .B(G952), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(G953), .ZN(new_n507));
  NAND2_X1  g321(.A1(G234), .A2(G237), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n248), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(G902), .A3(new_n508), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT21), .B(G898), .Z(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n510), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(G475), .A2(G902), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(KEYINPUT69), .A2(G953), .ZN(new_n519));
  NOR2_X1   g333(.A1(KEYINPUT69), .A2(G953), .ZN(new_n520));
  OAI211_X1 g334(.A(G214), .B(new_n249), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n188), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n248), .A2(G143), .A3(G214), .A4(new_n249), .ZN(new_n523));
  NAND2_X1  g337(.A1(KEYINPUT18), .A2(G131), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n341), .A2(new_n191), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n525), .B1(new_n344), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT18), .ZN(new_n528));
  AOI211_X1 g342(.A(new_n528), .B(new_n204), .C1(new_n522), .C2(new_n523), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT90), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n204), .B1(new_n522), .B2(new_n523), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT18), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n339), .A2(KEYINPUT78), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n341), .A2(new_n342), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n191), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n526), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT90), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n532), .A2(new_n537), .A3(new_n538), .A4(new_n525), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n522), .A2(new_n523), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(G131), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT19), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n341), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n340), .A2(new_n343), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n545), .B2(new_n543), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n348), .B1(new_n546), .B2(new_n191), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(G113), .B(G122), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(new_n388), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n354), .B1(KEYINPUT17), .B2(new_n531), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n542), .B2(KEYINPUT17), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n540), .A2(new_n555), .A3(new_n551), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n518), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT20), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT91), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n540), .A2(new_n555), .A3(new_n551), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n551), .B1(new_n540), .B2(new_n548), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n517), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT91), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT20), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n559), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G475), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n551), .B1(new_n540), .B2(new_n555), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n569), .B2(new_n298), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(G116), .B(G122), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(new_n385), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n196), .A2(G143), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n200), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n188), .A2(G128), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n574), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n578), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n222), .A2(G122), .ZN(new_n582));
  AND2_X1   g396(.A1(KEYINPUT14), .A2(G107), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n573), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n578), .B(G134), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n572), .A2(new_n583), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n581), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n500), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n590), .A2(new_n365), .A3(G953), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n581), .B(new_n591), .C1(new_n585), .C2(new_n588), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT92), .ZN(new_n596));
  INV_X1    g410(.A(G478), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(KEYINPUT15), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  OAI22_X1  g413(.A1(new_n595), .A2(KEYINPUT92), .B1(KEYINPUT15), .B2(new_n597), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n599), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n566), .A2(new_n571), .A3(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n505), .A2(new_n516), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n383), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT94), .B(G101), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G3));
  NOR2_X1   g420(.A1(new_n381), .A2(new_n516), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n298), .B1(new_n284), .B2(new_n294), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G472), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n295), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(new_n503), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n595), .A2(G478), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n593), .A2(new_n594), .ZN(new_n613));
  NAND2_X1  g427(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n597), .A2(G902), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n612), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n566), .B2(new_n571), .ZN(new_n620));
  INV_X1    g434(.A(new_n462), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n458), .A2(new_n459), .A3(new_n456), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n622), .B2(KEYINPUT95), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT95), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n455), .A2(new_n460), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n607), .A2(new_n611), .A3(new_n620), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G104), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  AND2_X1   g445(.A1(new_n566), .A2(new_n571), .ZN(new_n632));
  INV_X1    g446(.A(new_n516), .ZN(new_n633));
  INV_X1    g447(.A(new_n601), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n632), .A2(KEYINPUT98), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n566), .A2(new_n634), .A3(new_n571), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n636), .B1(new_n637), .B2(new_n516), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n381), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n627), .A3(new_n611), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n322), .A2(KEYINPUT36), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n356), .A2(KEYINPUT99), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n356), .A2(KEYINPUT99), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n646), .ZN(new_n648));
  INV_X1    g462(.A(new_n643), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n648), .A2(new_n649), .A3(new_n644), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n367), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(new_n375), .B2(new_n376), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n653), .A2(new_n602), .A3(new_n516), .ZN(new_n654));
  INV_X1    g468(.A(new_n610), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n464), .A2(new_n654), .A3(new_n504), .A4(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  INV_X1    g472(.A(new_n317), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n626), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n653), .A2(new_n503), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n509), .B1(new_n512), .B2(G900), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n637), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  XNOR2_X1  g481(.A(new_n662), .B(KEYINPUT39), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n504), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n254), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n280), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n267), .A2(new_n299), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n298), .B1(new_n675), .B2(new_n254), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n297), .A2(new_n312), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n566), .A2(new_n571), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n653), .A2(new_n679), .A3(new_n634), .A4(new_n462), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n461), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n671), .A2(new_n678), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  NAND2_X1  g499(.A1(new_n620), .A2(new_n662), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n686), .A2(new_n503), .A3(new_n653), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n660), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  AOI21_X1  g503(.A(new_n381), .B1(new_n315), .B2(new_n316), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n298), .B1(new_n484), .B2(new_n491), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(KEYINPUT102), .A3(new_n492), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n691), .A2(new_n694), .A3(G469), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n633), .A3(new_n502), .ZN(new_n697));
  INV_X1    g511(.A(new_n619), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n679), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n697), .A2(new_n699), .A3(new_n626), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n690), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND4_X1  g517(.A1(new_n696), .A2(new_n502), .A3(new_n625), .A4(new_n623), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n659), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n639), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n654), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  AND2_X1   g523(.A1(new_n300), .A2(new_n293), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n266), .B(new_n283), .C1(new_n254), .C2(new_n710), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n608), .A2(G472), .B1(new_n187), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n378), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n679), .A2(new_n634), .A3(new_n623), .A4(new_n625), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n713), .A2(new_n697), .A3(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n715), .B(G122), .Z(G24));
  NAND2_X1  g530(.A1(new_n492), .A2(KEYINPUT102), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n477), .A2(new_n480), .A3(new_n483), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n466), .A2(new_n470), .A3(new_n471), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n467), .B1(new_n719), .B2(KEYINPUT84), .ZN(new_n720));
  AOI22_X1  g534(.A1(new_n720), .A2(new_n489), .B1(new_n474), .B2(new_n476), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n718), .B1(new_n721), .B2(new_n480), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n465), .B1(new_n722), .B2(new_n298), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n695), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n502), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n626), .ZN(new_n727));
  INV_X1    g541(.A(new_n686), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n711), .A2(new_n187), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n609), .A2(new_n652), .A3(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n727), .A2(KEYINPUT103), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT103), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n712), .A2(new_n620), .A3(new_n652), .A4(new_n662), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n732), .B1(new_n733), .B2(new_n704), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  NAND2_X1  g550(.A1(new_n313), .A2(new_n378), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT107), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n313), .A2(new_n739), .A3(new_n378), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n455), .A2(new_n460), .A3(new_n462), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n480), .B1(new_n477), .B2(new_n483), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n495), .B1(new_n743), .B2(KEYINPUT104), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT104), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n721), .A2(new_n745), .A3(new_n480), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(G469), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n492), .A2(new_n494), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n744), .A2(KEYINPUT105), .A3(G469), .A4(new_n746), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT106), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n749), .A2(new_n750), .A3(KEYINPUT106), .A4(new_n751), .ZN(new_n755));
  AOI211_X1 g569(.A(new_n501), .B(new_n742), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n741), .A2(new_n728), .A3(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n690), .A2(new_n756), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n686), .A2(KEYINPUT42), .ZN(new_n759));
  AOI22_X1  g573(.A1(KEYINPUT42), .A2(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G131), .ZN(G33));
  NAND3_X1  g575(.A1(new_n690), .A2(new_n756), .A3(new_n664), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n497), .B1(new_n764), .B2(new_n465), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n744), .A2(new_n746), .ZN(new_n766));
  AOI22_X1  g580(.A1(KEYINPUT108), .A2(new_n765), .B1(new_n766), .B2(KEYINPUT45), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n765), .A2(KEYINPUT108), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n493), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(KEYINPUT46), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n492), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n769), .B2(KEYINPUT46), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n501), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n668), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n632), .A2(new_n698), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n776), .B1(KEYINPUT109), .B2(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n779));
  NAND3_X1  g593(.A1(new_n632), .A2(new_n698), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n655), .A2(new_n653), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(KEYINPUT44), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n742), .B(KEYINPUT110), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT44), .B1(new_n781), .B2(new_n782), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n775), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n202), .ZN(G39));
  NAND2_X1  g602(.A1(new_n769), .A2(KEYINPUT46), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n492), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n502), .B1(new_n790), .B2(new_n770), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT47), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT47), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n774), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n317), .A2(new_n378), .A3(new_n686), .A4(new_n742), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT111), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  XOR2_X1   g614(.A(new_n696), .B(KEYINPUT49), .Z(new_n801));
  NAND4_X1  g615(.A1(new_n682), .A2(new_n378), .A3(new_n502), .A4(new_n462), .ZN(new_n802));
  OR4_X1    g616(.A1(new_n678), .A2(new_n801), .A3(new_n776), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n804));
  INV_X1    g618(.A(new_n733), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n455), .A2(new_n460), .A3(new_n462), .A4(new_n662), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n632), .A2(new_n807), .A3(KEYINPUT114), .A4(new_n601), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n602), .B2(new_n806), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n808), .A2(new_n661), .A3(new_n810), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n805), .A2(new_n756), .B1(new_n811), .B2(new_n317), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n715), .B1(new_n690), .B2(new_n700), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n317), .B(new_n727), .C1(new_n639), .C2(new_n654), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n762), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n637), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n699), .A2(KEYINPUT112), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n699), .A2(KEYINPUT112), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n607), .A2(new_n464), .A3(new_n611), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n656), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n383), .B2(new_n603), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n815), .A2(new_n823), .A3(new_n760), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n317), .B(new_n627), .C1(new_n665), .C2(new_n687), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n651), .B(new_n662), .C1(new_n375), .C2(new_n376), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(KEYINPUT115), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(KEYINPUT115), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n827), .A2(new_n714), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n501), .B1(new_n754), .B2(new_n755), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n678), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n825), .A2(new_n735), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n825), .A2(new_n735), .A3(new_n831), .A4(KEYINPUT52), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n804), .B1(new_n824), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n757), .A2(KEYINPUT42), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n758), .A2(new_n759), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n812), .A2(new_n813), .A3(new_n762), .A4(new_n814), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n834), .A2(new_n835), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(KEYINPUT53), .A3(new_n843), .A4(new_n823), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n837), .A2(KEYINPUT116), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n824), .A2(new_n836), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT53), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n848), .A3(KEYINPUT54), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n837), .A2(KEYINPUT117), .A3(new_n844), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n851), .B(new_n804), .C1(new_n824), .C2(new_n836), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT54), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n849), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g669(.A(KEYINPUT118), .B(KEYINPUT54), .C1(new_n850), .C2(new_n852), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n381), .A2(new_n678), .A3(new_n509), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n726), .A2(new_n742), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n620), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n781), .A2(new_n378), .A3(new_n510), .A4(new_n712), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n860), .B(new_n507), .C1(new_n704), .C2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n509), .B1(new_n778), .B2(new_n780), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n863), .A2(new_n858), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n741), .ZN(new_n869));
  OR3_X1    g683(.A1(new_n868), .A2(KEYINPUT48), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT48), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n862), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n682), .A2(new_n502), .A3(new_n621), .A4(new_n696), .ZN(new_n873));
  OR3_X1    g687(.A1(new_n861), .A2(KEYINPUT50), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT50), .B1(new_n861), .B2(new_n873), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n859), .A2(new_n632), .A3(new_n619), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n730), .B1(new_n866), .B2(new_n867), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n792), .A2(new_n794), .B1(new_n501), .B2(new_n696), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n863), .A2(new_n378), .A3(new_n712), .A4(new_n784), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(KEYINPUT119), .A3(KEYINPUT51), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT51), .B1(new_n881), .B2(KEYINPUT119), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n872), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n855), .A2(new_n856), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(G952), .A2(G953), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT121), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n803), .B1(new_n886), .B2(new_n888), .ZN(G75));
  NAND4_X1  g703(.A1(new_n850), .A2(G210), .A3(G902), .A4(new_n852), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n423), .A2(new_n433), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n458), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n890), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n890), .B2(new_n891), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n248), .A2(G952), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G51));
  XNOR2_X1  g712(.A(new_n493), .B(KEYINPUT57), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n850), .A2(KEYINPUT54), .A3(new_n852), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(new_n853), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n722), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n850), .A2(new_n852), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n767), .A2(new_n768), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT122), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(G902), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n897), .B1(new_n902), .B2(new_n906), .ZN(G54));
  AND2_X1   g721(.A1(KEYINPUT58), .A2(G475), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n903), .A2(G902), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n553), .A2(new_n556), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n909), .A2(new_n911), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n913), .A3(new_n897), .ZN(G60));
  INV_X1    g728(.A(new_n617), .ZN(new_n915));
  NAND2_X1  g729(.A1(G478), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT59), .Z(new_n917));
  NOR2_X1   g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n900), .B2(new_n853), .ZN(new_n919));
  INV_X1    g733(.A(new_n897), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n917), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n855), .B2(new_n856), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n923), .B2(new_n915), .ZN(G63));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n925));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT60), .Z(new_n927));
  NAND3_X1  g741(.A1(new_n850), .A2(new_n852), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n364), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n647), .A2(new_n650), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n920), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n925), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n928), .A2(new_n931), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n934), .A2(KEYINPUT61), .A3(new_n920), .A4(new_n929), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n933), .A2(new_n935), .ZN(G66));
  OAI21_X1  g750(.A(G953), .B1(new_n515), .B2(new_n429), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n823), .A2(new_n813), .A3(new_n814), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(new_n511), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT123), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n457), .B(new_n416), .C1(G898), .C2(new_n248), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G69));
  XOR2_X1   g756(.A(new_n546), .B(KEYINPUT124), .Z(new_n943));
  XNOR2_X1  g757(.A(new_n264), .B(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(G227), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n248), .B1(new_n946), .B2(G900), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n787), .B1(new_n796), .B2(new_n798), .ZN(new_n948));
  INV_X1    g762(.A(new_n714), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n774), .A2(new_n668), .A3(new_n949), .A4(new_n741), .ZN(new_n950));
  AND4_X1   g764(.A1(new_n735), .A2(new_n950), .A3(new_n762), .A4(new_n825), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n948), .A2(new_n760), .A3(new_n951), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n952), .A2(new_n511), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n944), .B1(new_n945), .B2(new_n511), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n947), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n684), .A2(new_n825), .A3(new_n735), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT62), .Z(new_n957));
  NOR3_X1   g771(.A1(new_n820), .A2(new_n669), .A3(new_n742), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n383), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n948), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n948), .A2(new_n957), .A3(KEYINPUT125), .A4(new_n959), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n248), .A3(new_n944), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n955), .A2(new_n965), .ZN(G72));
  NAND2_X1  g780(.A1(G472), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT63), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n280), .A2(new_n254), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n969), .B2(new_n265), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n845), .A2(new_n848), .A3(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n971), .A2(KEYINPUT127), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n962), .A2(new_n938), .A3(new_n963), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n968), .B(KEYINPUT126), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n673), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n974), .B1(new_n952), .B2(new_n938), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n280), .A2(new_n672), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n920), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n971), .A2(KEYINPUT127), .ZN(new_n980));
  NOR4_X1   g794(.A1(new_n972), .A2(new_n976), .A3(new_n979), .A4(new_n980), .ZN(G57));
endmodule


