//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  XOR2_X1   g000(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT24), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n210));
  INV_X1    g009(.A(G169gat), .ZN(new_n211));
  INV_X1    g010(.A(G176gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n209), .A2(new_n210), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n202), .B1(new_n207), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n208), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(KEYINPUT23), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(new_n214), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n203), .B(KEYINPUT24), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n209), .A2(KEYINPUT25), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n222), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n221), .B1(new_n220), .B2(new_n214), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n216), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n218), .A2(new_n232), .A3(new_n219), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n233), .B(new_n214), .C1(new_n232), .C2(new_n208), .ZN(new_n234));
  AOI21_X1  g033(.A(G190gat), .B1(new_n223), .B2(KEYINPUT27), .ZN(new_n235));
  OR2_X1    g034(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(G183gat), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT28), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT27), .B(G183gat), .Z(new_n240));
  INV_X1    g039(.A(KEYINPUT28), .ZN(new_n241));
  NOR3_X1   g040(.A1(new_n240), .A2(new_n241), .A3(G190gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n203), .B(new_n234), .C1(new_n239), .C2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n231), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G226gat), .A2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT29), .B1(new_n231), .B2(new_n243), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n250), .A2(KEYINPUT71), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(KEYINPUT71), .ZN(new_n252));
  XNOR2_X1  g051(.A(G197gat), .B(G204gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G211gat), .B(G218gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n251), .A2(new_n255), .A3(new_n252), .A4(new_n253), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n249), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n247), .B(new_n259), .C1(new_n246), .C2(new_n248), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT37), .ZN(new_n264));
  XNOR2_X1  g063(.A(G8gat), .B(G36gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n265), .B(new_n266), .Z(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT37), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n261), .A2(new_n262), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n264), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT83), .B(KEYINPUT38), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n264), .A2(new_n268), .A3(new_n272), .A4(new_n270), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT2), .ZN(new_n277));
  INV_X1    g076(.A(G155gat), .ZN(new_n278));
  INV_X1    g077(.A(G162gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281));
  INV_X1    g080(.A(G141gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G148gat), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n280), .A2(new_n281), .B1(new_n283), .B2(KEYINPUT73), .ZN(new_n284));
  XNOR2_X1  g083(.A(G141gat), .B(G148gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G148gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(G141gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n277), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G155gat), .B(G162gat), .Z(new_n291));
  AOI22_X1  g090(.A1(new_n284), .A2(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G113gat), .ZN(new_n293));
  INV_X1    g092(.A(G120gat), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT1), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n293), .B2(new_n294), .ZN(new_n296));
  XNOR2_X1  g095(.A(G127gat), .B(G134gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n297), .B(new_n295), .C1(new_n293), .C2(new_n294), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n299), .A2(KEYINPUT69), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT69), .B1(new_n299), .B2(new_n300), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n292), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n284), .A2(new_n287), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n292), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n299), .A2(new_n300), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n292), .A2(new_n311), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n309), .A2(new_n312), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n308), .A2(new_n313), .A3(new_n304), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(KEYINPUT5), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n305), .A2(new_n315), .A3(new_n317), .A4(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n316), .B1(new_n303), .B2(new_n304), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n324), .A2(KEYINPUT76), .A3(new_n315), .A4(new_n320), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n292), .B(new_n313), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT5), .B1(new_n327), .B2(new_n318), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT75), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n292), .A2(new_n300), .A3(new_n299), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n319), .B1(new_n330), .B2(new_n304), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n315), .B(new_n331), .C1(new_n304), .C2(new_n303), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n333), .B(KEYINPUT5), .C1(new_n327), .C2(new_n318), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT0), .ZN(new_n338));
  XNOR2_X1  g137(.A(G57gat), .B(G85gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT6), .ZN(new_n342));
  INV_X1    g141(.A(new_n340), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n335), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n336), .A2(KEYINPUT6), .A3(new_n340), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n261), .A2(new_n262), .A3(new_n267), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n276), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n318), .B1(new_n324), .B2(new_n315), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n327), .A2(new_n318), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT39), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT39), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n340), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n350), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT40), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT81), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n360), .B1(new_n354), .B2(new_n356), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(KEYINPUT82), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n359), .A2(new_n362), .B1(new_n340), .B2(new_n336), .ZN(new_n363));
  OAI22_X1  g162(.A1(KEYINPUT82), .A2(new_n361), .B1(new_n357), .B2(new_n358), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n263), .A2(new_n268), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT30), .A4(new_n267), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT30), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n347), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n365), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  AND4_X1   g170(.A1(new_n365), .A2(new_n370), .A3(new_n366), .A4(new_n367), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n363), .B(new_n364), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G78gat), .B(G106gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT31), .B(G50gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n314), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT77), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n314), .A2(new_n381), .A3(new_n378), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n260), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT29), .B1(new_n257), .B2(new_n258), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n308), .B1(new_n384), .B2(KEYINPUT3), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n383), .A2(G228gat), .A3(G233gat), .A4(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(KEYINPUT78), .B(G22gat), .Z(new_n387));
  NAND2_X1  g186(.A1(new_n379), .A2(new_n260), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n385), .ZN(new_n389));
  INV_X1    g188(.A(G228gat), .ZN(new_n390));
  INV_X1    g189(.A(G233gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n386), .A2(new_n387), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n387), .B1(new_n386), .B2(new_n392), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n377), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n386), .A2(new_n392), .A3(new_n396), .A4(new_n387), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n386), .A2(new_n392), .ZN(new_n398));
  INV_X1    g197(.A(G22gat), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n397), .B(new_n376), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n393), .A2(new_n396), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n395), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n349), .A2(new_n373), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n345), .A2(new_n346), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT72), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n368), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n366), .A2(new_n367), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT72), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n404), .A2(new_n406), .A3(new_n370), .A4(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n402), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT36), .ZN(new_n411));
  XNOR2_X1  g210(.A(G15gat), .B(G43gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(G71gat), .B(G99gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n301), .A2(new_n302), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n244), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G227gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(new_n391), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n415), .A2(new_n231), .A3(new_n243), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n414), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(KEYINPUT32), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n421), .B(KEYINPUT32), .C1(new_n422), .C2(new_n414), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n419), .ZN(new_n428));
  INV_X1    g227(.A(new_n417), .ZN(new_n429));
  INV_X1    g228(.A(new_n420), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT34), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT34), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n433), .B(new_n428), .C1(new_n429), .C2(new_n430), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n427), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n427), .A2(new_n435), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n411), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n435), .A2(KEYINPUT70), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT70), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n432), .A2(new_n441), .A3(new_n434), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n427), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n435), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(new_n426), .A3(new_n425), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(KEYINPUT36), .A3(new_n445), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n409), .A2(new_n410), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n371), .A2(new_n372), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n402), .A2(new_n445), .A3(new_n436), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT35), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n404), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n402), .A2(new_n443), .A3(new_n445), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT35), .B1(new_n409), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n403), .A2(new_n447), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G15gat), .B(G22gat), .ZN(new_n455));
  INV_X1    g254(.A(G1gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT16), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(G8gat), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n458), .B(new_n459), .C1(G1gat), .C2(new_n455), .ZN(new_n460));
  INV_X1    g259(.A(G15gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G22gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n399), .A2(G15gat), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n457), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(G1gat), .B1(new_n462), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g264(.A(G8gat), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(G50gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G43gat), .ZN(new_n469));
  INV_X1    g268(.A(G43gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G50gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT15), .ZN(new_n472));
  INV_X1    g271(.A(G29gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT14), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT14), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(G29gat), .ZN(new_n476));
  INV_X1    g275(.A(G36gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n472), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n477), .B1(new_n473), .B2(KEYINPUT14), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n475), .A2(G29gat), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT85), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n469), .A2(new_n471), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n470), .A2(KEYINPUT85), .A3(G50gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT84), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT84), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT15), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n483), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n480), .B1(new_n492), .B2(new_n472), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT17), .B1(new_n493), .B2(KEYINPUT86), .ZN(new_n494));
  INV_X1    g293(.A(new_n472), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n469), .A2(new_n471), .A3(new_n484), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT84), .B(KEYINPUT15), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n486), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n495), .B1(new_n498), .B2(new_n483), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT17), .ZN(new_n501));
  NOR4_X1   g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .A4(new_n480), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n467), .B1(new_n494), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G229gat), .A2(G233gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n460), .A2(new_n466), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n493), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT18), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n504), .B(KEYINPUT13), .Z(new_n510));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n483), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n512), .A2(new_n496), .B1(new_n478), .B2(new_n479), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n511), .B1(new_n513), .B2(new_n495), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n467), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n493), .A2(new_n505), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT87), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n467), .A2(new_n514), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n506), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(KEYINPUT87), .A3(new_n510), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n503), .A2(KEYINPUT18), .A3(new_n504), .A4(new_n506), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(G197gat), .ZN(new_n527));
  XOR2_X1   g326(.A(KEYINPUT11), .B(G169gat), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(KEYINPUT12), .Z(new_n530));
  NAND2_X1  g329(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(KEYINPUT86), .B(new_n511), .C1(new_n513), .C2(new_n495), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n501), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n493), .A2(KEYINPUT86), .A3(KEYINPUT17), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n505), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n504), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n535), .A2(new_n536), .A3(new_n515), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n537), .A2(KEYINPUT18), .B1(new_n519), .B2(new_n522), .ZN(new_n538));
  INV_X1    g337(.A(new_n530), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n539), .A3(new_n509), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n531), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n454), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(KEYINPUT41), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(KEYINPUT90), .Z(new_n546));
  XNOR2_X1  g345(.A(G190gat), .B(G218gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT95), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n546), .B(new_n548), .Z(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551));
  AND2_X1   g350(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n552));
  NOR2_X1   g351(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT7), .ZN(new_n557));
  NAND2_X1  g356(.A1(G85gat), .A2(G92gat), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(KEYINPUT91), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(KEYINPUT91), .B2(new_n558), .ZN(new_n560));
  OAI211_X1 g359(.A(KEYINPUT93), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G99gat), .B(G106gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT94), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n565), .A2(KEYINPUT8), .ZN(new_n566));
  NOR2_X1   g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(KEYINPUT8), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n569), .B(KEYINPUT94), .C1(G85gat), .C2(G92gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n562), .A2(new_n563), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n563), .B1(new_n562), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n574), .A2(new_n493), .B1(KEYINPUT41), .B2(new_n544), .ZN(new_n575));
  OAI22_X1  g374(.A1(new_n494), .A2(new_n502), .B1(new_n572), .B2(new_n573), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n547), .A2(KEYINPUT95), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n580), .A2(new_n581), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n550), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(new_n549), .A3(new_n582), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G57gat), .B(G64gat), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n589), .A2(new_n590), .B1(KEYINPUT88), .B2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G71gat), .B(G78gat), .Z(new_n593));
  AND2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G127gat), .B(G155gat), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n467), .B1(new_n596), .B2(new_n597), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT89), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n602), .B(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n588), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n611), .B(new_n612), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n596), .B1(new_n572), .B2(new_n573), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n562), .A2(new_n571), .ZN(new_n617));
  INV_X1    g416(.A(new_n563), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n592), .B(new_n593), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n562), .A2(new_n563), .A3(new_n571), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n616), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n616), .A2(new_n622), .A3(KEYINPUT96), .A4(new_n623), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n574), .A2(KEYINPUT10), .A3(new_n620), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n615), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n616), .A2(new_n622), .ZN(new_n631));
  INV_X1    g430(.A(new_n615), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n614), .B1(new_n635), .B2(KEYINPUT97), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n637), .A3(new_n613), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n610), .A2(new_n639), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n640), .A2(KEYINPUT98), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(KEYINPUT98), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n543), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n404), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(new_n456), .ZN(G1324gat));
  INV_X1    g445(.A(new_n448), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n543), .A2(new_n647), .A3(new_n643), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n648), .A2(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(KEYINPUT99), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT16), .B(G8gat), .Z(new_n652));
  AOI21_X1  g451(.A(KEYINPUT42), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n649), .A2(G8gat), .A3(new_n650), .ZN(new_n654));
  INV_X1    g453(.A(new_n644), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n655), .A2(KEYINPUT42), .A3(new_n647), .A4(new_n652), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n658), .B1(new_n653), .B2(new_n657), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(G1325gat));
  NAND2_X1  g460(.A1(new_n439), .A2(new_n446), .ZN(new_n662));
  OAI21_X1  g461(.A(G15gat), .B1(new_n644), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n437), .A2(new_n438), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n461), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(new_n644), .B2(new_n665), .ZN(G1326gat));
  NOR2_X1   g465(.A1(new_n644), .A2(new_n402), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT43), .B(G22gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  INV_X1    g468(.A(new_n588), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n639), .A2(new_n609), .ZN(new_n671));
  NOR4_X1   g470(.A1(new_n454), .A2(new_n542), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n404), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(new_n473), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT45), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n454), .B2(new_n670), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n409), .A2(new_n410), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n354), .A2(new_n356), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n350), .B(KEYINPUT40), .C1(new_n679), .C2(new_n360), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n364), .A2(new_n680), .A3(new_n341), .ZN(new_n681));
  INV_X1    g480(.A(new_n371), .ZN(new_n682));
  INV_X1    g481(.A(new_n372), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n402), .B1(new_n276), .B2(new_n348), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n678), .B(new_n662), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n451), .A2(new_n453), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(KEYINPUT44), .A3(new_n588), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n677), .A2(new_n689), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n531), .A2(new_n540), .A3(KEYINPUT101), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT101), .B1(new_n531), .B2(new_n540), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n671), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G29gat), .B1(new_n695), .B2(new_n404), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n675), .A2(new_n696), .ZN(G1328gat));
  NAND3_X1  g496(.A1(new_n672), .A2(new_n477), .A3(new_n647), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n699), .B2(KEYINPUT46), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(KEYINPUT46), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n700), .B(new_n701), .Z(new_n702));
  NOR2_X1   g501(.A1(new_n695), .A2(new_n448), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n703), .A2(KEYINPUT103), .ZN(new_n704));
  OAI21_X1  g503(.A(G36gat), .B1(new_n703), .B2(KEYINPUT103), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(G1329gat));
  NOR3_X1   g505(.A1(new_n695), .A2(new_n470), .A3(new_n662), .ZN(new_n707));
  AOI21_X1  g506(.A(G43gat), .B1(new_n672), .B2(new_n664), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g509(.A1(new_n677), .A2(new_n689), .A3(new_n410), .A4(new_n694), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G50gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n672), .A2(new_n468), .A3(new_n410), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n714), .A2(KEYINPUT105), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(KEYINPUT105), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(KEYINPUT48), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  OAI22_X1  g520(.A1(new_n715), .A2(new_n716), .B1(KEYINPUT48), .B2(new_n719), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1331gat));
  INV_X1    g522(.A(new_n639), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n688), .A2(new_n610), .A3(new_n724), .A4(new_n693), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n404), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(G57gat), .Z(G1332gat));
  XOR2_X1   g526(.A(new_n725), .B(KEYINPUT106), .Z(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n647), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT49), .B(G64gat), .Z(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(G1333gat));
  INV_X1    g531(.A(new_n662), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n728), .A2(G71gat), .A3(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n725), .A2(new_n438), .A3(new_n437), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n736));
  INV_X1    g535(.A(G71gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n735), .B2(KEYINPUT107), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n734), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g539(.A1(new_n728), .A2(new_n410), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G78gat), .ZN(G1335gat));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n688), .A2(new_n588), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n539), .B1(new_n538), .B2(new_n509), .ZN(new_n746));
  AND4_X1   g545(.A1(new_n539), .A2(new_n509), .A3(new_n524), .A4(new_n523), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n531), .A2(new_n540), .A3(KEYINPUT101), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n609), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n743), .B1(new_n744), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n688), .A2(KEYINPUT51), .A3(new_n588), .A4(new_n752), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(new_n639), .ZN(new_n759));
  INV_X1    g558(.A(G85gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n760), .A3(new_n673), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n753), .A2(new_n639), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n677), .A2(new_n689), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT108), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n677), .A2(new_n689), .A3(new_n765), .A4(new_n762), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n764), .A2(new_n673), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n761), .B1(new_n760), .B2(new_n767), .ZN(G1336gat));
  NOR2_X1   g567(.A1(new_n448), .A2(G92gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n759), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(G92gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n763), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n647), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n764), .A2(new_n647), .A3(new_n766), .ZN(new_n776));
  AOI22_X1  g575(.A1(new_n759), .A2(new_n769), .B1(G92gat), .B2(new_n776), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n772), .A2(new_n775), .B1(new_n777), .B2(new_n771), .ZN(G1337gat));
  INV_X1    g577(.A(G99gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n759), .A2(new_n779), .A3(new_n664), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n764), .A2(new_n733), .A3(new_n766), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n779), .B2(new_n781), .ZN(G1338gat));
  OAI21_X1  g581(.A(G106gat), .B1(new_n763), .B2(new_n402), .ZN(new_n783));
  XNOR2_X1  g582(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n639), .A2(G106gat), .A3(new_n402), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n783), .B(new_n784), .C1(new_n758), .C2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n764), .A2(new_n410), .A3(new_n766), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G106gat), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n785), .B(KEYINPUT109), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n754), .B2(new_n756), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n788), .B1(new_n795), .B2(KEYINPUT53), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n793), .B1(new_n789), .B2(G106gat), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n797), .A2(KEYINPUT110), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n787), .B1(new_n796), .B2(new_n799), .ZN(G1339gat));
  NOR2_X1   g599(.A1(new_n634), .A2(new_n614), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n624), .A2(new_n625), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n802), .A2(new_n632), .A3(new_n627), .A4(new_n628), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n630), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n805), .B(new_n615), .C1(new_n626), .C2(new_n629), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n614), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n801), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n804), .A2(KEYINPUT55), .A3(new_n614), .A4(new_n806), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n750), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n504), .B1(new_n503), .B2(new_n506), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n521), .A2(new_n510), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n529), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n540), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n636), .A2(new_n638), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n588), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n630), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n806), .A2(new_n614), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n808), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n801), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n810), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n588), .A2(new_n815), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n609), .B1(new_n817), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n640), .A2(new_n750), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n448), .A2(new_n673), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n452), .ZN(new_n832));
  AOI21_X1  g631(.A(G113gat), .B1(new_n832), .B2(new_n750), .ZN(new_n833));
  INV_X1    g632(.A(new_n449), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n542), .A2(new_n293), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(G1340gat));
  NAND3_X1  g636(.A1(new_n832), .A2(new_n294), .A3(new_n724), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n724), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n839), .A2(KEYINPUT112), .A3(G120gat), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT112), .B1(new_n839), .B2(G120gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  XOR2_X1   g641(.A(new_n842), .B(KEYINPUT113), .Z(G1341gat));
  INV_X1    g642(.A(new_n832), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(G127gat), .A3(new_n609), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n835), .A2(new_n751), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(G127gat), .B2(new_n846), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT114), .Z(G1342gat));
  NOR3_X1   g647(.A1(new_n844), .A2(G134gat), .A3(new_n670), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT56), .ZN(new_n850));
  INV_X1    g649(.A(new_n831), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n449), .A3(new_n588), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(G134gat), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(KEYINPUT115), .Z(new_n854));
  NAND2_X1  g653(.A1(new_n850), .A2(new_n854), .ZN(G1343gat));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n402), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n820), .A2(new_n541), .A3(new_n821), .A4(new_n810), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n816), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n670), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n824), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n861), .A2(KEYINPUT117), .A3(new_n670), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n751), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n859), .B1(new_n866), .B2(new_n826), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n816), .B1(new_n822), .B2(new_n693), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n670), .ZN(new_n869));
  INV_X1    g668(.A(new_n824), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n826), .B1(new_n871), .B2(new_n609), .ZN(new_n872));
  OAI211_X1 g671(.A(KEYINPUT116), .B(new_n858), .C1(new_n872), .C2(new_n402), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n402), .B1(new_n825), .B2(new_n827), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(KEYINPUT57), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n867), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n733), .A2(new_n829), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n750), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G141gat), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n875), .A2(new_n282), .A3(new_n541), .A4(new_n878), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT118), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n857), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n857), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n877), .A2(new_n541), .A3(new_n878), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(G141gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n856), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(G141gat), .ZN(new_n889));
  INV_X1    g688(.A(new_n885), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n882), .B1(new_n879), .B2(G141gat), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n891), .B(KEYINPUT119), .C1(new_n857), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n888), .A2(new_n893), .ZN(G1344gat));
  AND2_X1   g693(.A1(new_n875), .A2(new_n878), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n288), .A3(new_n724), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n877), .A2(new_n878), .ZN(new_n897));
  AOI211_X1 g696(.A(KEYINPUT59), .B(new_n288), .C1(new_n897), .C2(new_n724), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n862), .A2(new_n870), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n609), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n641), .A2(new_n542), .A3(new_n642), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n410), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n858), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n875), .A2(KEYINPUT57), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n639), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n878), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n899), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n896), .B1(new_n898), .B2(new_n911), .ZN(G1345gat));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n278), .A3(new_n751), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n897), .A2(new_n751), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n278), .ZN(G1346gat));
  NOR2_X1   g714(.A1(new_n670), .A2(new_n279), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n733), .A2(new_n402), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n851), .A2(new_n588), .A3(new_n917), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n897), .A2(new_n916), .B1(new_n279), .B2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n448), .A2(new_n673), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n828), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n452), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(G169gat), .B1(new_n924), .B2(new_n750), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n920), .B(KEYINPUT121), .Z(new_n926));
  NOR3_X1   g725(.A1(new_n926), .A2(new_n872), .A3(new_n834), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n542), .A2(new_n211), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(G1348gat));
  INV_X1    g728(.A(new_n927), .ZN(new_n930));
  OAI21_X1  g729(.A(G176gat), .B1(new_n930), .B2(new_n639), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n724), .A2(new_n212), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n923), .B2(new_n932), .ZN(G1349gat));
  NOR3_X1   g732(.A1(new_n923), .A2(new_n240), .A3(new_n609), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n223), .B1(new_n927), .B2(new_n751), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1350gat));
  AOI21_X1  g737(.A(new_n224), .B1(new_n927), .B2(new_n588), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT61), .Z(new_n940));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n224), .A3(new_n588), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1351gat));
  AND2_X1   g741(.A1(new_n921), .A2(new_n917), .ZN(new_n943));
  AOI21_X1  g742(.A(G197gat), .B1(new_n943), .B2(new_n750), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n907), .A2(new_n908), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n926), .A2(new_n733), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n541), .A2(G197gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(G1352gat));
  XNOR2_X1  g749(.A(KEYINPUT123), .B(G204gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n951), .B1(new_n909), .B2(new_n946), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n921), .A2(new_n724), .A3(new_n917), .A4(new_n951), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT62), .ZN(new_n955));
  OR3_X1    g754(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n952), .B2(new_n955), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1353gat));
  OAI21_X1  g757(.A(G211gat), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(new_n947), .B2(new_n609), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(KEYINPUT125), .A3(KEYINPUT63), .ZN(new_n962));
  NAND2_X1  g761(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n960), .B(new_n963), .C1(new_n947), .C2(new_n609), .ZN(new_n964));
  INV_X1    g763(.A(G211gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n943), .A2(new_n965), .A3(new_n751), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n962), .A2(new_n964), .A3(new_n966), .ZN(G1354gat));
  AOI21_X1  g766(.A(G218gat), .B1(new_n943), .B2(new_n588), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n968), .B(KEYINPUT126), .Z(new_n969));
  NAND2_X1  g768(.A1(new_n588), .A2(G218gat), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n970), .B1(new_n948), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n947), .A2(KEYINPUT127), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(G1355gat));
endmodule


