

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(n655), .A2(n614), .ZN(n864) );
  AND2_X1 U554 ( .A1(G2104), .A2(G2105), .ZN(n955) );
  XNOR2_X1 U555 ( .A(KEYINPUT70), .B(n607), .ZN(n860) );
  INV_X1 U556 ( .A(n557), .ZN(G160) );
  AND2_X1 U557 ( .A1(n769), .A2(n768), .ZN(n520) );
  NOR2_X2 U558 ( .A1(n573), .A2(n572), .ZN(n744) );
  INV_X1 U559 ( .A(n771), .ZN(n781) );
  AND2_X1 U560 ( .A1(n788), .A2(G137), .ZN(n635) );
  XNOR2_X1 U561 ( .A(G2104), .B(KEYINPUT66), .ZN(n626) );
  AND2_X1 U562 ( .A1(n677), .A2(G40), .ZN(n555) );
  OR2_X1 U563 ( .A1(n567), .A2(KEYINPUT32), .ZN(n564) );
  INV_X1 U564 ( .A(KEYINPUT33), .ZN(n592) );
  AND2_X1 U565 ( .A1(n711), .A2(n682), .ZN(n683) );
  OR2_X1 U566 ( .A1(n764), .A2(n719), .ZN(n721) );
  NAND2_X1 U567 ( .A1(n579), .A2(n571), .ZN(n574) );
  AND2_X1 U568 ( .A1(n739), .A2(KEYINPUT29), .ZN(n571) );
  XNOR2_X1 U569 ( .A(n535), .B(n534), .ZN(n750) );
  INV_X1 U570 ( .A(KEYINPUT94), .ZN(n534) );
  NAND2_X1 U571 ( .A1(n741), .A2(n742), .ZN(n535) );
  AND2_X1 U572 ( .A1(n550), .A2(KEYINPUT64), .ZN(n549) );
  NAND2_X1 U573 ( .A1(n548), .A2(n555), .ZN(n547) );
  NAND2_X1 U574 ( .A1(n557), .A2(KEYINPUT64), .ZN(n556) );
  OR2_X1 U575 ( .A1(n761), .A2(KEYINPUT32), .ZN(n563) );
  AND2_X1 U576 ( .A1(n568), .A2(G8), .ZN(n567) );
  OR2_X1 U577 ( .A1(G286), .A2(n569), .ZN(n568) );
  OR2_X1 U578 ( .A1(n772), .A2(n593), .ZN(n589) );
  NAND2_X1 U579 ( .A1(n772), .A2(n591), .ZN(n590) );
  OR2_X1 U580 ( .A1(n1052), .A2(n593), .ZN(n591) );
  AND2_X1 U581 ( .A1(n522), .A2(n592), .ZN(n586) );
  NAND2_X1 U582 ( .A1(n595), .A2(n594), .ZN(n956) );
  NAND2_X1 U583 ( .A1(n526), .A2(n597), .ZN(n594) );
  NAND2_X1 U584 ( .A1(n596), .A2(KEYINPUT67), .ZN(n595) );
  NAND2_X1 U585 ( .A1(n537), .A2(n1039), .ZN(n776) );
  XNOR2_X1 U586 ( .A(n539), .B(n538), .ZN(n537) );
  INV_X1 U587 ( .A(KEYINPUT102), .ZN(n538) );
  INV_X1 U588 ( .A(KEYINPUT97), .ZN(n687) );
  OR2_X1 U589 ( .A1(n740), .A2(n1064), .ZN(n722) );
  BUF_X1 U590 ( .A(n711), .Z(n740) );
  NOR2_X1 U591 ( .A1(G168), .A2(n748), .ZN(n749) );
  AND2_X1 U592 ( .A1(n556), .A2(n554), .ZN(n553) );
  NAND2_X1 U593 ( .A1(G160), .A2(n525), .ZN(n551) );
  NAND2_X1 U594 ( .A1(n549), .A2(n547), .ZN(n554) );
  AND2_X1 U595 ( .A1(n565), .A2(n561), .ZN(n560) );
  NAND2_X1 U596 ( .A1(n564), .A2(n562), .ZN(n561) );
  NAND2_X1 U597 ( .A1(n567), .A2(n563), .ZN(n562) );
  NAND2_X1 U598 ( .A1(n762), .A2(n528), .ZN(n558) );
  INV_X1 U599 ( .A(KEYINPUT32), .ZN(n559) );
  AND2_X1 U600 ( .A1(n764), .A2(G8), .ZN(n771) );
  INV_X1 U601 ( .A(KEYINPUT67), .ZN(n602) );
  OR2_X1 U602 ( .A1(n626), .A2(n625), .ZN(n596) );
  INV_X1 U603 ( .A(n626), .ZN(n597) );
  NAND2_X1 U604 ( .A1(n540), .A2(n587), .ZN(n539) );
  AND2_X1 U605 ( .A1(n585), .A2(n530), .ZN(n540) );
  INV_X1 U606 ( .A(G125), .ZN(n599) );
  INV_X1 U607 ( .A(G651), .ZN(n614) );
  AND2_X1 U608 ( .A1(n622), .A2(n621), .ZN(n604) );
  BUF_X1 U609 ( .A(n956), .Z(n536) );
  NOR2_X2 U610 ( .A1(G2104), .A2(G2105), .ZN(n624) );
  AND2_X1 U611 ( .A1(n546), .A2(n581), .ZN(n545) );
  NOR2_X1 U612 ( .A1(n582), .A2(n529), .ZN(n581) );
  NAND2_X1 U613 ( .A1(n544), .A2(n523), .ZN(n543) );
  NOR2_X1 U614 ( .A1(G651), .A2(G543), .ZN(n865) );
  NOR2_X1 U615 ( .A1(G651), .A2(n655), .ZN(n859) );
  INV_X1 U616 ( .A(KEYINPUT6), .ZN(n611) );
  XOR2_X1 U617 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  OR2_X1 U618 ( .A1(n819), .A2(n829), .ZN(n521) );
  AND2_X1 U619 ( .A1(n772), .A2(KEYINPUT65), .ZN(n522) );
  AND2_X1 U620 ( .A1(n521), .A2(KEYINPUT105), .ZN(n523) );
  OR2_X1 U621 ( .A1(n784), .A2(n783), .ZN(n524) );
  AND2_X1 U622 ( .A1(n678), .A2(n552), .ZN(n525) );
  AND2_X1 U623 ( .A1(G2105), .A2(n602), .ZN(n526) );
  XOR2_X1 U624 ( .A(n743), .B(KEYINPUT95), .Z(n527) );
  AND2_X1 U625 ( .A1(n567), .A2(n559), .ZN(n528) );
  NOR2_X1 U626 ( .A1(n820), .A2(n829), .ZN(n529) );
  OR2_X1 U627 ( .A1(n781), .A2(n774), .ZN(n530) );
  AND2_X1 U628 ( .A1(n583), .A2(n592), .ZN(n531) );
  NAND2_X1 U629 ( .A1(n1052), .A2(n593), .ZN(n532) );
  AND2_X1 U630 ( .A1(G160), .A2(G40), .ZN(n533) );
  INV_X1 U631 ( .A(KEYINPUT65), .ZN(n593) );
  AND2_X1 U632 ( .A1(n576), .A2(n527), .ZN(n575) );
  INV_X1 U633 ( .A(n570), .ZN(n762) );
  NAND2_X1 U634 ( .A1(n570), .A2(n566), .ZN(n565) );
  XNOR2_X2 U635 ( .A(n756), .B(KEYINPUT101), .ZN(n570) );
  NOR2_X1 U636 ( .A1(n542), .A2(KEYINPUT105), .ZN(n541) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n573) );
  NOR2_X1 U638 ( .A1(n684), .A2(n683), .ZN(n686) );
  XNOR2_X2 U639 ( .A(n776), .B(KEYINPUT104), .ZN(n580) );
  NOR2_X1 U640 ( .A1(n781), .A2(G1966), .ZN(n766) );
  NAND2_X1 U641 ( .A1(n637), .A2(n636), .ZN(n557) );
  NOR2_X1 U642 ( .A1(n736), .A2(n731), .ZN(n737) );
  NAND2_X1 U643 ( .A1(n580), .A2(n524), .ZN(n544) );
  NAND2_X1 U644 ( .A1(n580), .A2(n541), .ZN(n546) );
  INV_X1 U645 ( .A(n524), .ZN(n542) );
  NAND2_X1 U646 ( .A1(n545), .A2(n543), .ZN(n833) );
  INV_X1 U647 ( .A(n604), .ZN(n548) );
  NAND2_X1 U648 ( .A1(n631), .A2(n555), .ZN(n550) );
  NAND2_X1 U649 ( .A1(n604), .A2(n632), .ZN(n678) );
  NAND2_X1 U650 ( .A1(n678), .A2(n677), .ZN(n818) );
  NAND2_X4 U651 ( .A1(n553), .A2(n551), .ZN(n764) );
  AND2_X1 U652 ( .A1(n555), .A2(n679), .ZN(n552) );
  NAND2_X1 U653 ( .A1(n560), .A2(n558), .ZN(n769) );
  AND2_X1 U654 ( .A1(n761), .A2(KEYINPUT32), .ZN(n566) );
  INV_X1 U655 ( .A(n761), .ZN(n569) );
  NAND2_X1 U656 ( .A1(n520), .A2(n586), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n734), .A2(n735), .ZN(n579) );
  NOR2_X1 U658 ( .A1(n579), .A2(KEYINPUT29), .ZN(n572) );
  NAND2_X1 U659 ( .A1(n578), .A2(n577), .ZN(n576) );
  INV_X1 U660 ( .A(KEYINPUT29), .ZN(n577) );
  INV_X1 U661 ( .A(n739), .ZN(n578) );
  NOR2_X1 U662 ( .A1(n521), .A2(KEYINPUT105), .ZN(n582) );
  NAND2_X1 U663 ( .A1(n584), .A2(n531), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n588), .A2(n532), .ZN(n583) );
  NAND2_X1 U665 ( .A1(n520), .A2(n588), .ZN(n584) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n588) );
  INV_X1 U667 ( .A(n956), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n600), .A2(n598), .ZN(n636) );
  NAND2_X1 U669 ( .A1(n603), .A2(n599), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n601), .A2(n603), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n766), .A2(n745), .ZN(n746) );
  NOR2_X1 U672 ( .A1(n635), .A2(n605), .ZN(n603) );
  AND2_X1 U673 ( .A1(G113), .A2(n955), .ZN(n605) );
  NOR2_X1 U674 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n685) );
  NOR2_X1 U675 ( .A1(n773), .A2(n770), .ZN(n1052) );
  INV_X1 U676 ( .A(KEYINPUT75), .ZN(n693) );
  INV_X1 U677 ( .A(KEYINPUT17), .ZN(n623) );
  XNOR2_X1 U678 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U679 ( .A(n696), .B(n695), .ZN(n701) );
  XNOR2_X1 U680 ( .A(n612), .B(n611), .ZN(n619) );
  INV_X1 U681 ( .A(n716), .ZN(n1057) );
  NOR2_X1 U682 ( .A1(n644), .A2(n643), .ZN(G171) );
  NOR2_X1 U683 ( .A1(G543), .A2(n614), .ZN(n606) );
  XOR2_X1 U684 ( .A(KEYINPUT1), .B(n606), .Z(n607) );
  NAND2_X1 U685 ( .A1(G63), .A2(n860), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n608), .B(KEYINPUT76), .ZN(n610) );
  XOR2_X1 U687 ( .A(G543), .B(KEYINPUT0), .Z(n655) );
  NAND2_X1 U688 ( .A1(G51), .A2(n859), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n865), .A2(G89), .ZN(n613) );
  XNOR2_X1 U691 ( .A(n613), .B(KEYINPUT4), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G76), .A2(n864), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n617), .B(KEYINPUT5), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n620), .B(KEYINPUT7), .ZN(G168) );
  INV_X1 U697 ( .A(G2105), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n956), .A2(G126), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n955), .A2(G114), .ZN(n621) );
  XNOR2_X2 U700 ( .A(n624), .B(n623), .ZN(n788) );
  NAND2_X1 U701 ( .A1(n788), .A2(G138), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n628) );
  INV_X1 U703 ( .A(KEYINPUT68), .ZN(n627) );
  XNOR2_X2 U704 ( .A(n628), .B(n627), .ZN(n785) );
  NAND2_X1 U705 ( .A1(n785), .A2(G102), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n631) );
  INV_X1 U707 ( .A(n631), .ZN(n632) );
  INV_X1 U708 ( .A(n678), .ZN(G164) );
  NAND2_X1 U709 ( .A1(n785), .A2(G101), .ZN(n634) );
  INV_X1 U710 ( .A(KEYINPUT23), .ZN(n633) );
  XNOR2_X1 U711 ( .A(n634), .B(n633), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n859), .A2(G52), .ZN(n639) );
  NAND2_X1 U713 ( .A1(G64), .A2(n860), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n644) );
  NAND2_X1 U715 ( .A1(G77), .A2(n864), .ZN(n641) );
  NAND2_X1 U716 ( .A1(G90), .A2(n865), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U718 ( .A(KEYINPUT9), .B(n642), .Z(n643) );
  AND2_X1 U719 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U720 ( .A(G57), .ZN(G237) );
  INV_X1 U721 ( .A(G69), .ZN(G235) );
  INV_X1 U722 ( .A(G108), .ZN(G238) );
  INV_X1 U723 ( .A(G120), .ZN(G236) );
  INV_X1 U724 ( .A(G132), .ZN(G219) );
  INV_X1 U725 ( .A(G82), .ZN(G220) );
  NAND2_X1 U726 ( .A1(n865), .A2(G86), .ZN(n646) );
  NAND2_X1 U727 ( .A1(G61), .A2(n860), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U729 ( .A(KEYINPUT82), .B(n647), .ZN(n651) );
  NAND2_X1 U730 ( .A1(G73), .A2(n864), .ZN(n648) );
  XNOR2_X1 U731 ( .A(n648), .B(KEYINPUT83), .ZN(n649) );
  XNOR2_X1 U732 ( .A(n649), .B(KEYINPUT2), .ZN(n650) );
  NOR2_X1 U733 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U734 ( .A1(n859), .A2(G48), .ZN(n652) );
  NAND2_X1 U735 ( .A1(n653), .A2(n652), .ZN(G305) );
  NAND2_X1 U736 ( .A1(G74), .A2(G651), .ZN(n654) );
  XNOR2_X1 U737 ( .A(n654), .B(KEYINPUT80), .ZN(n658) );
  NAND2_X1 U738 ( .A1(G87), .A2(n655), .ZN(n656) );
  XOR2_X1 U739 ( .A(KEYINPUT81), .B(n656), .Z(n657) );
  NAND2_X1 U740 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U741 ( .A1(n860), .A2(n659), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n859), .A2(G49), .ZN(n660) );
  NAND2_X1 U743 ( .A1(n661), .A2(n660), .ZN(G288) );
  NAND2_X1 U744 ( .A1(G75), .A2(n864), .ZN(n663) );
  NAND2_X1 U745 ( .A1(G88), .A2(n865), .ZN(n662) );
  NAND2_X1 U746 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U747 ( .A(KEYINPUT84), .B(n664), .Z(n668) );
  NAND2_X1 U748 ( .A1(n860), .A2(G62), .ZN(n666) );
  NAND2_X1 U749 ( .A1(n859), .A2(G50), .ZN(n665) );
  AND2_X1 U750 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U751 ( .A1(n668), .A2(n667), .ZN(G303) );
  INV_X1 U752 ( .A(G303), .ZN(G166) );
  NAND2_X1 U753 ( .A1(n859), .A2(G47), .ZN(n670) );
  NAND2_X1 U754 ( .A1(G60), .A2(n860), .ZN(n669) );
  NAND2_X1 U755 ( .A1(n670), .A2(n669), .ZN(n673) );
  NAND2_X1 U756 ( .A1(G72), .A2(n864), .ZN(n671) );
  XNOR2_X1 U757 ( .A(KEYINPUT69), .B(n671), .ZN(n672) );
  NOR2_X1 U758 ( .A1(n673), .A2(n672), .ZN(n675) );
  NAND2_X1 U759 ( .A1(n865), .A2(G85), .ZN(n674) );
  NAND2_X1 U760 ( .A1(n675), .A2(n674), .ZN(G290) );
  INV_X1 U761 ( .A(G1384), .ZN(n677) );
  INV_X1 U762 ( .A(KEYINPUT64), .ZN(n679) );
  INV_X1 U763 ( .A(G1341), .ZN(n680) );
  AND2_X1 U764 ( .A1(n680), .A2(KEYINPUT26), .ZN(n681) );
  AND2_X1 U765 ( .A1(n764), .A2(n681), .ZN(n684) );
  INV_X1 U766 ( .A(n764), .ZN(n711) );
  NAND2_X1 U767 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n682) );
  NOR2_X1 U768 ( .A1(n686), .A2(n685), .ZN(n688) );
  XNOR2_X1 U769 ( .A(n688), .B(n687), .ZN(n717) );
  NAND2_X1 U770 ( .A1(n865), .A2(G81), .ZN(n689) );
  XOR2_X1 U771 ( .A(KEYINPUT12), .B(n689), .Z(n692) );
  NAND2_X1 U772 ( .A1(n864), .A2(G68), .ZN(n690) );
  XOR2_X1 U773 ( .A(n690), .B(KEYINPUT74), .Z(n691) );
  NOR2_X1 U774 ( .A1(n692), .A2(n691), .ZN(n696) );
  INV_X1 U775 ( .A(KEYINPUT13), .ZN(n694) );
  NAND2_X1 U776 ( .A1(G56), .A2(n860), .ZN(n697) );
  XNOR2_X1 U777 ( .A(n697), .B(KEYINPUT14), .ZN(n699) );
  NAND2_X1 U778 ( .A1(G43), .A2(n859), .ZN(n698) );
  AND2_X1 U779 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U780 ( .A1(n701), .A2(n700), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n859), .A2(G54), .ZN(n703) );
  NAND2_X1 U782 ( .A1(G66), .A2(n860), .ZN(n702) );
  NAND2_X1 U783 ( .A1(n703), .A2(n702), .ZN(n707) );
  NAND2_X1 U784 ( .A1(G79), .A2(n864), .ZN(n705) );
  NAND2_X1 U785 ( .A1(G92), .A2(n865), .ZN(n704) );
  NAND2_X1 U786 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U787 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U788 ( .A(n708), .B(KEYINPUT15), .ZN(n1042) );
  NOR2_X1 U789 ( .A1(n716), .A2(n1042), .ZN(n709) );
  NAND2_X1 U790 ( .A1(n717), .A2(n709), .ZN(n710) );
  XNOR2_X1 U791 ( .A(n710), .B(KEYINPUT98), .ZN(n715) );
  NAND2_X1 U792 ( .A1(n764), .A2(G1348), .ZN(n713) );
  NAND2_X1 U793 ( .A1(n740), .A2(G2067), .ZN(n712) );
  NAND2_X1 U794 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U795 ( .A1(n715), .A2(n714), .ZN(n735) );
  NAND2_X1 U796 ( .A1(n717), .A2(n1057), .ZN(n718) );
  NAND2_X1 U797 ( .A1(n718), .A2(n1042), .ZN(n733) );
  INV_X1 U798 ( .A(G2072), .ZN(n719) );
  XOR2_X1 U799 ( .A(KEYINPUT27), .B(KEYINPUT96), .Z(n720) );
  XNOR2_X1 U800 ( .A(n721), .B(n720), .ZN(n723) );
  INV_X1 U801 ( .A(G1956), .ZN(n1064) );
  NAND2_X1 U802 ( .A1(n723), .A2(n722), .ZN(n736) );
  NAND2_X1 U803 ( .A1(G65), .A2(n860), .ZN(n726) );
  NAND2_X1 U804 ( .A1(G78), .A2(n864), .ZN(n724) );
  XOR2_X1 U805 ( .A(KEYINPUT71), .B(n724), .Z(n725) );
  NAND2_X1 U806 ( .A1(n726), .A2(n725), .ZN(n730) );
  NAND2_X1 U807 ( .A1(G53), .A2(n859), .ZN(n728) );
  NAND2_X1 U808 ( .A1(G91), .A2(n865), .ZN(n727) );
  NAND2_X1 U809 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U810 ( .A1(n730), .A2(n729), .ZN(n1046) );
  INV_X1 U811 ( .A(n1046), .ZN(n731) );
  NAND2_X1 U812 ( .A1(n736), .A2(n731), .ZN(n732) );
  XNOR2_X1 U813 ( .A(n732), .B(KEYINPUT28), .ZN(n738) );
  AND2_X1 U814 ( .A1(n733), .A2(n738), .ZN(n734) );
  NAND2_X1 U815 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U816 ( .A1(n764), .A2(G1961), .ZN(n742) );
  XOR2_X1 U817 ( .A(KEYINPUT25), .B(G2078), .Z(n998) );
  NAND2_X1 U818 ( .A1(n740), .A2(n998), .ZN(n741) );
  NAND2_X1 U819 ( .A1(n750), .A2(G171), .ZN(n743) );
  XNOR2_X1 U820 ( .A(n744), .B(KEYINPUT99), .ZN(n755) );
  NOR2_X1 U821 ( .A1(n764), .A2(G2084), .ZN(n745) );
  NAND2_X1 U822 ( .A1(n746), .A2(G8), .ZN(n747) );
  XNOR2_X1 U823 ( .A(n747), .B(KEYINPUT30), .ZN(n748) );
  XNOR2_X1 U824 ( .A(n749), .B(KEYINPUT100), .ZN(n752) );
  NOR2_X1 U825 ( .A1(n750), .A2(G171), .ZN(n751) );
  NOR2_X1 U826 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U827 ( .A(KEYINPUT31), .B(n753), .Z(n754) );
  NAND2_X1 U828 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U829 ( .A1(n764), .A2(G2090), .ZN(n757) );
  NOR2_X1 U830 ( .A1(n757), .A2(G166), .ZN(n760) );
  INV_X1 U831 ( .A(G1971), .ZN(n758) );
  NAND2_X1 U832 ( .A1(n771), .A2(n758), .ZN(n759) );
  NAND2_X1 U833 ( .A1(n760), .A2(n759), .ZN(n761) );
  INV_X1 U834 ( .A(G2084), .ZN(n1019) );
  NAND2_X1 U835 ( .A1(n1019), .A2(G8), .ZN(n763) );
  NOR2_X1 U836 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U837 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U838 ( .A1(n762), .A2(n767), .ZN(n768) );
  NOR2_X1 U839 ( .A1(G288), .A2(G1976), .ZN(n773) );
  NOR2_X1 U840 ( .A1(G303), .A2(G1971), .ZN(n770) );
  NAND2_X1 U841 ( .A1(G288), .A2(G1976), .ZN(n1047) );
  AND2_X1 U842 ( .A1(n771), .A2(n1047), .ZN(n772) );
  NAND2_X1 U843 ( .A1(n773), .A2(KEYINPUT33), .ZN(n774) );
  XNOR2_X1 U844 ( .A(G1981), .B(KEYINPUT103), .ZN(n775) );
  XNOR2_X1 U845 ( .A(G305), .B(n775), .ZN(n1039) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U847 ( .A1(G8), .A2(n777), .ZN(n778) );
  NAND2_X1 U848 ( .A1(n781), .A2(n778), .ZN(n779) );
  NOR2_X1 U849 ( .A1(n520), .A2(n779), .ZN(n784) );
  NOR2_X1 U850 ( .A1(G305), .A2(G1981), .ZN(n780) );
  XNOR2_X1 U851 ( .A(n780), .B(KEYINPUT24), .ZN(n782) );
  NOR2_X1 U852 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U853 ( .A(G2067), .B(KEYINPUT37), .ZN(n827) );
  BUF_X1 U854 ( .A(n785), .Z(n786) );
  NAND2_X1 U855 ( .A1(n786), .A2(G104), .ZN(n787) );
  XOR2_X1 U856 ( .A(KEYINPUT89), .B(n787), .Z(n790) );
  NAND2_X1 U857 ( .A1(n788), .A2(G140), .ZN(n789) );
  NAND2_X1 U858 ( .A1(n790), .A2(n789), .ZN(n792) );
  XNOR2_X1 U859 ( .A(KEYINPUT90), .B(KEYINPUT34), .ZN(n791) );
  XNOR2_X1 U860 ( .A(n792), .B(n791), .ZN(n797) );
  NAND2_X1 U861 ( .A1(G116), .A2(n955), .ZN(n794) );
  NAND2_X1 U862 ( .A1(G128), .A2(n536), .ZN(n793) );
  NAND2_X1 U863 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U864 ( .A(KEYINPUT35), .B(n795), .Z(n796) );
  NOR2_X1 U865 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U866 ( .A(KEYINPUT36), .B(n798), .ZN(n965) );
  NOR2_X1 U867 ( .A1(n827), .A2(n965), .ZN(n1033) );
  NAND2_X1 U868 ( .A1(G107), .A2(n955), .ZN(n800) );
  NAND2_X1 U869 ( .A1(G119), .A2(n536), .ZN(n799) );
  NAND2_X1 U870 ( .A1(n800), .A2(n799), .ZN(n804) );
  NAND2_X1 U871 ( .A1(G131), .A2(n788), .ZN(n802) );
  NAND2_X1 U872 ( .A1(n786), .A2(G95), .ZN(n801) );
  NAND2_X1 U873 ( .A1(n802), .A2(n801), .ZN(n803) );
  OR2_X1 U874 ( .A1(n804), .A2(n803), .ZN(n950) );
  NAND2_X1 U875 ( .A1(G1991), .A2(n950), .ZN(n805) );
  XNOR2_X1 U876 ( .A(n805), .B(KEYINPUT91), .ZN(n816) );
  NAND2_X1 U877 ( .A1(n786), .A2(G105), .ZN(n807) );
  XOR2_X1 U878 ( .A(KEYINPUT93), .B(KEYINPUT38), .Z(n806) );
  XNOR2_X1 U879 ( .A(n807), .B(n806), .ZN(n814) );
  NAND2_X1 U880 ( .A1(G141), .A2(n788), .ZN(n809) );
  NAND2_X1 U881 ( .A1(G129), .A2(n536), .ZN(n808) );
  NAND2_X1 U882 ( .A1(n809), .A2(n808), .ZN(n812) );
  NAND2_X1 U883 ( .A1(n955), .A2(G117), .ZN(n810) );
  XOR2_X1 U884 ( .A(KEYINPUT92), .B(n810), .Z(n811) );
  NOR2_X1 U885 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U886 ( .A1(n814), .A2(n813), .ZN(n945) );
  AND2_X1 U887 ( .A1(G1996), .A2(n945), .ZN(n815) );
  NOR2_X1 U888 ( .A1(n816), .A2(n815), .ZN(n1023) );
  INV_X1 U889 ( .A(n1023), .ZN(n817) );
  NOR2_X1 U890 ( .A1(n1033), .A2(n817), .ZN(n819) );
  NAND2_X1 U891 ( .A1(n818), .A2(n533), .ZN(n829) );
  XNOR2_X1 U892 ( .A(G290), .B(G1986), .ZN(n1054) );
  INV_X1 U893 ( .A(n1054), .ZN(n820) );
  INV_X1 U894 ( .A(n1033), .ZN(n826) );
  NOR2_X1 U895 ( .A1(G1996), .A2(n945), .ZN(n1013) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U897 ( .A1(G1991), .A2(n950), .ZN(n1016) );
  NOR2_X1 U898 ( .A1(n821), .A2(n1016), .ZN(n822) );
  NOR2_X1 U899 ( .A1(n817), .A2(n822), .ZN(n823) );
  NOR2_X1 U900 ( .A1(n1013), .A2(n823), .ZN(n824) );
  XNOR2_X1 U901 ( .A(n824), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U902 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U903 ( .A1(n827), .A2(n965), .ZN(n1030) );
  NAND2_X1 U904 ( .A1(n828), .A2(n1030), .ZN(n831) );
  INV_X1 U905 ( .A(n829), .ZN(n830) );
  NAND2_X1 U906 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U907 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U908 ( .A(n834), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U909 ( .A1(G7), .A2(G661), .ZN(n835) );
  XNOR2_X1 U910 ( .A(n835), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U911 ( .A(G223), .B(KEYINPUT73), .ZN(n898) );
  NAND2_X1 U912 ( .A1(n898), .A2(G567), .ZN(n836) );
  XOR2_X1 U913 ( .A(KEYINPUT11), .B(n836), .Z(G234) );
  NAND2_X1 U914 ( .A1(n1057), .A2(G860), .ZN(G153) );
  INV_X1 U915 ( .A(G171), .ZN(G301) );
  NAND2_X1 U916 ( .A1(G868), .A2(G301), .ZN(n838) );
  INV_X1 U917 ( .A(G868), .ZN(n871) );
  NAND2_X1 U918 ( .A1(n1042), .A2(n871), .ZN(n837) );
  NAND2_X1 U919 ( .A1(n838), .A2(n837), .ZN(G284) );
  XOR2_X1 U920 ( .A(n1046), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U921 ( .A1(G299), .A2(G868), .ZN(n840) );
  NOR2_X1 U922 ( .A1(G286), .A2(n871), .ZN(n839) );
  NOR2_X1 U923 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U924 ( .A(KEYINPUT77), .B(n841), .Z(G297) );
  INV_X1 U925 ( .A(G860), .ZN(n842) );
  NAND2_X1 U926 ( .A1(G559), .A2(n842), .ZN(n843) );
  XNOR2_X1 U927 ( .A(KEYINPUT78), .B(n843), .ZN(n844) );
  INV_X1 U928 ( .A(n1042), .ZN(n970) );
  NAND2_X1 U929 ( .A1(n844), .A2(n970), .ZN(n845) );
  XNOR2_X1 U930 ( .A(KEYINPUT16), .B(n845), .ZN(G148) );
  NAND2_X1 U931 ( .A1(n970), .A2(G868), .ZN(n846) );
  NOR2_X1 U932 ( .A1(G559), .A2(n846), .ZN(n848) );
  AND2_X1 U933 ( .A1(n871), .A2(n1057), .ZN(n847) );
  NOR2_X1 U934 ( .A1(n848), .A2(n847), .ZN(G282) );
  NAND2_X1 U935 ( .A1(G135), .A2(n788), .ZN(n850) );
  NAND2_X1 U936 ( .A1(G111), .A2(n955), .ZN(n849) );
  NAND2_X1 U937 ( .A1(n850), .A2(n849), .ZN(n855) );
  NAND2_X1 U938 ( .A1(G123), .A2(n536), .ZN(n851) );
  XNOR2_X1 U939 ( .A(n851), .B(KEYINPUT18), .ZN(n853) );
  NAND2_X1 U940 ( .A1(n786), .A2(G99), .ZN(n852) );
  NAND2_X1 U941 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U942 ( .A1(n855), .A2(n854), .ZN(n1015) );
  XNOR2_X1 U943 ( .A(n1015), .B(G2096), .ZN(n857) );
  INV_X1 U944 ( .A(G2100), .ZN(n856) );
  NAND2_X1 U945 ( .A1(n857), .A2(n856), .ZN(G156) );
  NAND2_X1 U946 ( .A1(G559), .A2(n970), .ZN(n858) );
  XOR2_X1 U947 ( .A(n1057), .B(n858), .Z(n880) );
  NOR2_X1 U948 ( .A1(n880), .A2(G860), .ZN(n870) );
  NAND2_X1 U949 ( .A1(n859), .A2(G55), .ZN(n862) );
  NAND2_X1 U950 ( .A1(G67), .A2(n860), .ZN(n861) );
  NAND2_X1 U951 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U952 ( .A(KEYINPUT79), .B(n863), .ZN(n869) );
  NAND2_X1 U953 ( .A1(G80), .A2(n864), .ZN(n867) );
  NAND2_X1 U954 ( .A1(G93), .A2(n865), .ZN(n866) );
  AND2_X1 U955 ( .A1(n867), .A2(n866), .ZN(n868) );
  NAND2_X1 U956 ( .A1(n869), .A2(n868), .ZN(n873) );
  XOR2_X1 U957 ( .A(n870), .B(n873), .Z(G145) );
  NAND2_X1 U958 ( .A1(n871), .A2(n873), .ZN(n872) );
  XNOR2_X1 U959 ( .A(n872), .B(KEYINPUT86), .ZN(n883) );
  XOR2_X1 U960 ( .A(n873), .B(G299), .Z(n879) );
  XNOR2_X1 U961 ( .A(KEYINPUT19), .B(G305), .ZN(n874) );
  XNOR2_X1 U962 ( .A(n874), .B(G288), .ZN(n875) );
  XNOR2_X1 U963 ( .A(KEYINPUT85), .B(n875), .ZN(n877) );
  XNOR2_X1 U964 ( .A(G290), .B(G166), .ZN(n876) );
  XNOR2_X1 U965 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U966 ( .A(n879), .B(n878), .ZN(n969) );
  XNOR2_X1 U967 ( .A(n969), .B(n880), .ZN(n881) );
  NAND2_X1 U968 ( .A1(G868), .A2(n881), .ZN(n882) );
  NAND2_X1 U969 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U970 ( .A(KEYINPUT87), .B(n884), .Z(G295) );
  NAND2_X1 U971 ( .A1(G2078), .A2(G2084), .ZN(n885) );
  XOR2_X1 U972 ( .A(KEYINPUT20), .B(n885), .Z(n886) );
  NAND2_X1 U973 ( .A1(G2090), .A2(n886), .ZN(n887) );
  XNOR2_X1 U974 ( .A(KEYINPUT21), .B(n887), .ZN(n888) );
  NAND2_X1 U975 ( .A1(n888), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U976 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U977 ( .A1(G220), .A2(G219), .ZN(n889) );
  XOR2_X1 U978 ( .A(KEYINPUT22), .B(n889), .Z(n890) );
  NOR2_X1 U979 ( .A1(G218), .A2(n890), .ZN(n891) );
  NAND2_X1 U980 ( .A1(G96), .A2(n891), .ZN(n902) );
  NAND2_X1 U981 ( .A1(n902), .A2(G2106), .ZN(n896) );
  NOR2_X1 U982 ( .A1(G236), .A2(G238), .ZN(n893) );
  NOR2_X1 U983 ( .A1(G235), .A2(G237), .ZN(n892) );
  NAND2_X1 U984 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U985 ( .A(KEYINPUT88), .B(n894), .ZN(n903) );
  NAND2_X1 U986 ( .A1(n903), .A2(G567), .ZN(n895) );
  NAND2_X1 U987 ( .A1(n896), .A2(n895), .ZN(n904) );
  NAND2_X1 U988 ( .A1(G483), .A2(G661), .ZN(n897) );
  NOR2_X1 U989 ( .A1(n904), .A2(n897), .ZN(n901) );
  NAND2_X1 U990 ( .A1(n901), .A2(G36), .ZN(G176) );
  NAND2_X1 U991 ( .A1(G2106), .A2(n898), .ZN(G217) );
  AND2_X1 U992 ( .A1(G15), .A2(G2), .ZN(n899) );
  NAND2_X1 U993 ( .A1(G661), .A2(n899), .ZN(G259) );
  NAND2_X1 U994 ( .A1(G3), .A2(G1), .ZN(n900) );
  NAND2_X1 U995 ( .A1(n901), .A2(n900), .ZN(G188) );
  INV_X1 U997 ( .A(G96), .ZN(G221) );
  NOR2_X1 U998 ( .A1(n903), .A2(n902), .ZN(G325) );
  INV_X1 U999 ( .A(G325), .ZN(G261) );
  INV_X1 U1000 ( .A(n904), .ZN(G319) );
  XOR2_X1 U1001 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G2678), .B(KEYINPUT43), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U1004 ( .A(KEYINPUT42), .B(G2090), .Z(n908) );
  XNOR2_X1 U1005 ( .A(G2067), .B(G2072), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1007 ( .A(n910), .B(n909), .Z(n912) );
  XNOR2_X1 U1008 ( .A(G2096), .B(G2100), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n914) );
  XOR2_X1 U1010 ( .A(G2078), .B(G2084), .Z(n913) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(G227) );
  XOR2_X1 U1012 ( .A(G1981), .B(G1966), .Z(n916) );
  XNOR2_X1 U1013 ( .A(G1996), .B(G1991), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n926) );
  XOR2_X1 U1015 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n918) );
  XNOR2_X1 U1016 ( .A(G1961), .B(KEYINPUT110), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n918), .B(n917), .ZN(n922) );
  XOR2_X1 U1018 ( .A(G1976), .B(G1971), .Z(n920) );
  XNOR2_X1 U1019 ( .A(G1986), .B(G1956), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1021 ( .A(n922), .B(n921), .Z(n924) );
  XNOR2_X1 U1022 ( .A(G2474), .B(KEYINPUT41), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(n924), .B(n923), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n926), .B(n925), .ZN(G229) );
  NAND2_X1 U1025 ( .A1(G136), .A2(n788), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(G112), .A2(n955), .ZN(n927) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n934) );
  NAND2_X1 U1028 ( .A1(G124), .A2(n536), .ZN(n929) );
  XOR2_X1 U1029 ( .A(KEYINPUT113), .B(n929), .Z(n930) );
  XNOR2_X1 U1030 ( .A(n930), .B(KEYINPUT44), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n786), .A2(G100), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(G162) );
  NAND2_X1 U1034 ( .A1(G142), .A2(n788), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n786), .A2(G106), .ZN(n935) );
  NAND2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(n937), .B(KEYINPUT45), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(G130), .A2(n536), .ZN(n938) );
  NAND2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(n955), .A2(G118), .ZN(n940) );
  XOR2_X1 U1041 ( .A(KEYINPUT114), .B(n940), .Z(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n954) );
  XOR2_X1 U1043 ( .A(KEYINPUT46), .B(KEYINPUT116), .Z(n944) );
  XNOR2_X1 U1044 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(n944), .B(n943), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(n1015), .B(n945), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(G160), .B(G164), .ZN(n946) );
  XNOR2_X1 U1048 ( .A(n947), .B(n946), .ZN(n948) );
  XNOR2_X1 U1049 ( .A(n949), .B(n948), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(n950), .B(G162), .ZN(n951) );
  XNOR2_X1 U1051 ( .A(n952), .B(n951), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(n954), .B(n953), .ZN(n967) );
  NAND2_X1 U1053 ( .A1(G115), .A2(n955), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(G127), .A2(n536), .ZN(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(n959), .B(KEYINPUT47), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(n786), .A2(G103), .ZN(n960) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(G139), .A2(n788), .ZN(n962) );
  XNOR2_X1 U1060 ( .A(KEYINPUT115), .B(n962), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n1024) );
  XNOR2_X1 U1062 ( .A(n965), .B(n1024), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(n967), .B(n966), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(G37), .A2(n968), .ZN(G395) );
  XOR2_X1 U1065 ( .A(n969), .B(G286), .Z(n972) );
  XNOR2_X1 U1066 ( .A(n970), .B(G171), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(n972), .B(n971), .ZN(n973) );
  XOR2_X1 U1068 ( .A(n1057), .B(n973), .Z(n974) );
  NOR2_X1 U1069 ( .A1(G37), .A2(n974), .ZN(G397) );
  XNOR2_X1 U1070 ( .A(G2443), .B(G2427), .ZN(n984) );
  XOR2_X1 U1071 ( .A(G2430), .B(KEYINPUT107), .Z(n976) );
  XNOR2_X1 U1072 ( .A(G2454), .B(G2435), .ZN(n975) );
  XNOR2_X1 U1073 ( .A(n976), .B(n975), .ZN(n980) );
  XOR2_X1 U1074 ( .A(G2438), .B(KEYINPUT106), .Z(n978) );
  XNOR2_X1 U1075 ( .A(G1341), .B(G1348), .ZN(n977) );
  XNOR2_X1 U1076 ( .A(n978), .B(n977), .ZN(n979) );
  XOR2_X1 U1077 ( .A(n980), .B(n979), .Z(n982) );
  XNOR2_X1 U1078 ( .A(G2451), .B(G2446), .ZN(n981) );
  XNOR2_X1 U1079 ( .A(n982), .B(n981), .ZN(n983) );
  XNOR2_X1 U1080 ( .A(n984), .B(n983), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n985), .A2(G14), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(G319), .A2(n991), .ZN(n988) );
  NOR2_X1 U1083 ( .A1(G227), .A2(G229), .ZN(n986) );
  XNOR2_X1 U1084 ( .A(KEYINPUT49), .B(n986), .ZN(n987) );
  NOR2_X1 U1085 ( .A1(n988), .A2(n987), .ZN(n990) );
  NOR2_X1 U1086 ( .A1(G395), .A2(G397), .ZN(n989) );
  NAND2_X1 U1087 ( .A1(n990), .A2(n989), .ZN(G225) );
  INV_X1 U1088 ( .A(G225), .ZN(G308) );
  INV_X1 U1089 ( .A(n991), .ZN(G401) );
  XNOR2_X1 U1090 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n1099) );
  XOR2_X1 U1091 ( .A(G32), .B(G1996), .Z(n1002) );
  XOR2_X1 U1092 ( .A(G1991), .B(G25), .Z(n992) );
  NAND2_X1 U1093 ( .A1(G28), .A2(n992), .ZN(n993) );
  XNOR2_X1 U1094 ( .A(n993), .B(KEYINPUT119), .ZN(n997) );
  XNOR2_X1 U1095 ( .A(G2067), .B(G26), .ZN(n995) );
  XNOR2_X1 U1096 ( .A(G2072), .B(G33), .ZN(n994) );
  NOR2_X1 U1097 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1098 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XNOR2_X1 U1099 ( .A(G27), .B(n998), .ZN(n999) );
  NOR2_X1 U1100 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1101 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1102 ( .A(KEYINPUT53), .B(n1003), .ZN(n1007) );
  XOR2_X1 U1103 ( .A(G34), .B(KEYINPUT120), .Z(n1005) );
  XNOR2_X1 U1104 ( .A(G2084), .B(KEYINPUT54), .ZN(n1004) );
  XNOR2_X1 U1105 ( .A(n1005), .B(n1004), .ZN(n1006) );
  NAND2_X1 U1106 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XNOR2_X1 U1107 ( .A(G35), .B(G2090), .ZN(n1008) );
  NOR2_X1 U1108 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1109 ( .A(KEYINPUT55), .B(n1010), .Z(n1011) );
  NOR2_X1 U1110 ( .A1(G29), .A2(n1011), .ZN(n1097) );
  XOR2_X1 U1111 ( .A(G2090), .B(G162), .Z(n1012) );
  NOR2_X1 U1112 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1113 ( .A(KEYINPUT51), .B(n1014), .Z(n1018) );
  NOR2_X1 U1114 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1115 ( .A1(n1018), .A2(n1017), .ZN(n1021) );
  XNOR2_X1 U1116 ( .A(G160), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1117 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1118 ( .A1(n1023), .A2(n1022), .ZN(n1029) );
  XOR2_X1 U1119 ( .A(G2072), .B(n1024), .Z(n1026) );
  XOR2_X1 U1120 ( .A(G164), .B(G2078), .Z(n1025) );
  NOR2_X1 U1121 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1122 ( .A(KEYINPUT50), .B(n1027), .Z(n1028) );
  NOR2_X1 U1123 ( .A1(n1029), .A2(n1028), .ZN(n1031) );
  NAND2_X1 U1124 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1125 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1126 ( .A(KEYINPUT52), .B(n1034), .ZN(n1036) );
  INV_X1 U1127 ( .A(KEYINPUT55), .ZN(n1035) );
  NAND2_X1 U1128 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1129 ( .A1(n1037), .A2(G29), .ZN(n1038) );
  XOR2_X1 U1130 ( .A(KEYINPUT118), .B(n1038), .Z(n1094) );
  XNOR2_X1 U1131 ( .A(G16), .B(KEYINPUT56), .ZN(n1063) );
  XNOR2_X1 U1132 ( .A(G1966), .B(G168), .ZN(n1040) );
  NAND2_X1 U1133 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1134 ( .A(n1041), .B(KEYINPUT57), .ZN(n1061) );
  XOR2_X1 U1135 ( .A(n1042), .B(G1348), .Z(n1044) );
  XNOR2_X1 U1136 ( .A(G171), .B(G1961), .ZN(n1043) );
  NAND2_X1 U1137 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XNOR2_X1 U1138 ( .A(KEYINPUT121), .B(n1045), .ZN(n1056) );
  XNOR2_X1 U1139 ( .A(n1046), .B(G1956), .ZN(n1048) );
  NAND2_X1 U1140 ( .A1(n1048), .A2(n1047), .ZN(n1050) );
  AND2_X1 U1141 ( .A1(G303), .A2(G1971), .ZN(n1049) );
  NOR2_X1 U1142 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  NAND2_X1 U1143 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
  NOR2_X1 U1144 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
  NAND2_X1 U1145 ( .A1(n1056), .A2(n1055), .ZN(n1059) );
  XOR2_X1 U1146 ( .A(n1057), .B(G1341), .Z(n1058) );
  NOR2_X1 U1147 ( .A1(n1059), .A2(n1058), .ZN(n1060) );
  NAND2_X1 U1148 ( .A1(n1061), .A2(n1060), .ZN(n1062) );
  NAND2_X1 U1149 ( .A1(n1063), .A2(n1062), .ZN(n1092) );
  INV_X1 U1150 ( .A(G16), .ZN(n1090) );
  XNOR2_X1 U1151 ( .A(n1064), .B(G20), .ZN(n1072) );
  XOR2_X1 U1152 ( .A(G1981), .B(G6), .Z(n1067) );
  XOR2_X1 U1153 ( .A(G19), .B(KEYINPUT122), .Z(n1065) );
  XNOR2_X1 U1154 ( .A(G1341), .B(n1065), .ZN(n1066) );
  NAND2_X1 U1155 ( .A1(n1067), .A2(n1066), .ZN(n1070) );
  XOR2_X1 U1156 ( .A(KEYINPUT59), .B(G1348), .Z(n1068) );
  XNOR2_X1 U1157 ( .A(G4), .B(n1068), .ZN(n1069) );
  NOR2_X1 U1158 ( .A1(n1070), .A2(n1069), .ZN(n1071) );
  NAND2_X1 U1159 ( .A1(n1072), .A2(n1071), .ZN(n1073) );
  XNOR2_X1 U1160 ( .A(n1073), .B(KEYINPUT123), .ZN(n1074) );
  XOR2_X1 U1161 ( .A(KEYINPUT60), .B(n1074), .Z(n1076) );
  XNOR2_X1 U1162 ( .A(G1961), .B(G5), .ZN(n1075) );
  NOR2_X1 U1163 ( .A1(n1076), .A2(n1075), .ZN(n1086) );
  XNOR2_X1 U1164 ( .A(G1971), .B(G22), .ZN(n1078) );
  XNOR2_X1 U1165 ( .A(G1976), .B(G23), .ZN(n1077) );
  NOR2_X1 U1166 ( .A1(n1078), .A2(n1077), .ZN(n1079) );
  XOR2_X1 U1167 ( .A(KEYINPUT124), .B(n1079), .Z(n1081) );
  XNOR2_X1 U1168 ( .A(G1986), .B(G24), .ZN(n1080) );
  NOR2_X1 U1169 ( .A1(n1081), .A2(n1080), .ZN(n1082) );
  XOR2_X1 U1170 ( .A(KEYINPUT58), .B(n1082), .Z(n1084) );
  XNOR2_X1 U1171 ( .A(G1966), .B(G21), .ZN(n1083) );
  NOR2_X1 U1172 ( .A1(n1084), .A2(n1083), .ZN(n1085) );
  NAND2_X1 U1173 ( .A1(n1086), .A2(n1085), .ZN(n1087) );
  XNOR2_X1 U1174 ( .A(n1087), .B(KEYINPUT61), .ZN(n1088) );
  XNOR2_X1 U1175 ( .A(KEYINPUT125), .B(n1088), .ZN(n1089) );
  NAND2_X1 U1176 ( .A1(n1090), .A2(n1089), .ZN(n1091) );
  NAND2_X1 U1177 ( .A1(n1092), .A2(n1091), .ZN(n1093) );
  NOR2_X1 U1178 ( .A1(n1094), .A2(n1093), .ZN(n1095) );
  NAND2_X1 U1179 ( .A1(n1095), .A2(G11), .ZN(n1096) );
  NOR2_X1 U1180 ( .A1(n1097), .A2(n1096), .ZN(n1098) );
  XNOR2_X1 U1181 ( .A(n1099), .B(n1098), .ZN(n1100) );
  XNOR2_X1 U1182 ( .A(KEYINPUT62), .B(n1100), .ZN(G150) );
  INV_X1 U1183 ( .A(G150), .ZN(G311) );
endmodule

