//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT66), .A2(G134), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT66), .A2(G134), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n193), .B1(new_n196), .B2(G137), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n192), .B1(new_n194), .B2(new_n195), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n197), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n203), .B1(new_n197), .B2(new_n202), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n212), .A3(G143), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n209), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n219));
  OAI21_X1  g033(.A(G128), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n213), .A2(G128), .A3(new_n222), .A4(new_n215), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G107), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT78), .B1(new_n225), .B2(G104), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT78), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G107), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(G104), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G101), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(G107), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n225), .A2(KEYINPUT3), .A3(G104), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT3), .B1(new_n225), .B2(G104), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n233), .B(new_n234), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n224), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT79), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n232), .A2(new_n240), .A3(new_n237), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n219), .A2(KEYINPUT68), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT1), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n243), .B1(new_n213), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n210), .A2(new_n212), .ZN(new_n249));
  INV_X1    g063(.A(G143), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n218), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n223), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n240), .B1(new_n232), .B2(new_n237), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n242), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT80), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n239), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n213), .A2(new_n247), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G128), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT64), .B(G146), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n217), .B1(new_n259), .B2(G143), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n214), .B1(new_n259), .B2(G143), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n247), .A2(new_n243), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n258), .A2(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n232), .A2(new_n237), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT79), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n265), .A3(new_n241), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(KEYINPUT80), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n208), .B1(new_n256), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT12), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n264), .B1(new_n223), .B2(new_n221), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n266), .B2(KEYINPUT80), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n254), .A2(new_n255), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n207), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT12), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT10), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n239), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(KEYINPUT10), .B(new_n252), .C1(new_n242), .C2(new_n253), .ZN(new_n278));
  AND2_X1   g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n213), .A2(new_n215), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(KEYINPUT0), .A2(G128), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n280), .B1(new_n251), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(G101), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(G101), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT4), .A3(new_n237), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n285), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n277), .A2(new_n278), .A3(new_n207), .A4(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G953), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G227), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n294), .B(KEYINPUT77), .ZN(new_n295));
  XNOR2_X1  g109(.A(G110), .B(G140), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n269), .A2(new_n275), .A3(new_n292), .A4(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n278), .A2(new_n277), .A3(new_n291), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n300), .A2(new_n208), .ZN(new_n301));
  INV_X1    g115(.A(new_n292), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n297), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI211_X1 g117(.A(G469), .B(G902), .C1(new_n299), .C2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G469), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n292), .B1(new_n273), .B2(new_n274), .ZN(new_n306));
  AOI211_X1 g120(.A(KEYINPUT12), .B(new_n207), .C1(new_n271), .C2(new_n272), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n297), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n301), .A2(new_n302), .A3(new_n297), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n305), .B1(new_n311), .B2(new_n190), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT81), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n304), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n269), .A2(new_n275), .A3(new_n292), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n309), .B1(new_n315), .B2(new_n297), .ZN(new_n316));
  OAI21_X1  g130(.A(G469), .B1(new_n316), .B2(G902), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT81), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n191), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G110), .B(G122), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G113), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n323));
  INV_X1    g137(.A(G119), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n324), .A2(G116), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n322), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(G116), .B(G119), .Z(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(new_n323), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT2), .B(G113), .Z(new_n329));
  XNOR2_X1  g143(.A(G116), .B(G119), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(new_n265), .B2(new_n241), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n329), .B(new_n330), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n290), .A2(new_n334), .A3(new_n288), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n321), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n327), .A2(new_n323), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n337), .A2(new_n326), .B1(new_n330), .B2(new_n329), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n242), .B2(new_n253), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n290), .A2(new_n334), .A3(new_n288), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(new_n320), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(KEYINPUT6), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n284), .A2(G125), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n344), .B(new_n223), .C1(new_n248), .C2(new_n251), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n293), .A2(G224), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n347), .B(KEYINPUT85), .Z(new_n348));
  XOR2_X1   g162(.A(new_n346), .B(new_n348), .Z(new_n349));
  INV_X1    g163(.A(KEYINPUT6), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(new_n321), .C1(new_n333), .C2(new_n335), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n342), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n320), .B(KEYINPUT8), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n330), .A2(KEYINPUT5), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n326), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n331), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n265), .B2(new_n241), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n338), .A2(new_n238), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n347), .A2(KEYINPUT7), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n346), .B(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(KEYINPUT86), .B(new_n353), .C1(new_n357), .C2(new_n358), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n361), .A2(new_n363), .A3(new_n341), .A4(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n352), .A2(new_n190), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(G210), .B1(G237), .B2(G902), .ZN(new_n367));
  XOR2_X1   g181(.A(new_n367), .B(KEYINPUT87), .Z(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n352), .A2(new_n190), .A3(new_n365), .A4(new_n368), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(G214), .B1(G237), .B2(G902), .ZN(new_n374));
  XOR2_X1   g188(.A(new_n374), .B(KEYINPUT82), .Z(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT83), .ZN(new_n376));
  NAND2_X1  g190(.A1(G234), .A2(G237), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(G952), .A3(new_n293), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(KEYINPUT92), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(G902), .A3(G953), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT21), .B(G898), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n373), .A2(new_n376), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G140), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G125), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n344), .A2(G140), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT75), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .A4(KEYINPUT16), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT16), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT16), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n387), .A3(G125), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT75), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n209), .B(new_n391), .C1(new_n392), .C2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n388), .A2(new_n389), .ZN(new_n398));
  OAI211_X1 g212(.A(KEYINPUT75), .B(new_n394), .C1(new_n398), .C2(new_n393), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n209), .B1(new_n399), .B2(new_n391), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(G237), .A2(G953), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n402), .A2(G143), .A3(G214), .ZN(new_n403));
  AOI21_X1  g217(.A(G143), .B1(new_n402), .B2(G214), .ZN(new_n404));
  OAI21_X1  g218(.A(G131), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G237), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n293), .A3(G214), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n250), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n402), .A2(G143), .A3(G214), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n203), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n405), .A2(new_n410), .A3(KEYINPUT88), .A4(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT88), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n405), .A2(new_n410), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(KEYINPUT17), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n408), .A2(new_n409), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT17), .A3(G131), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n401), .A2(new_n412), .A3(new_n415), .A4(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n388), .A2(new_n389), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n259), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n209), .B2(new_n419), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n416), .A2(KEYINPUT18), .A3(G131), .ZN(new_n422));
  NAND2_X1  g236(.A1(KEYINPUT18), .A2(G131), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n408), .A2(new_n409), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G113), .B(G122), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(G104), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(KEYINPUT89), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n190), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n418), .B2(new_n425), .ZN(new_n433));
  OAI21_X1  g247(.A(G475), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n425), .A2(new_n428), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n419), .B(KEYINPUT19), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n400), .B1(new_n259), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n414), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n426), .B2(new_n429), .ZN(new_n440));
  NOR2_X1   g254(.A1(G475), .A2(G902), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n435), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n428), .B1(new_n418), .B2(new_n425), .ZN(new_n443));
  INV_X1    g257(.A(new_n441), .ZN(new_n444));
  NOR4_X1   g258(.A1(new_n443), .A2(new_n439), .A3(KEYINPUT20), .A4(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n434), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n189), .A2(G217), .A3(new_n293), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G122), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G116), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n225), .B1(new_n451), .B2(KEYINPUT14), .ZN(new_n452));
  XNOR2_X1  g266(.A(G116), .B(G122), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n250), .A2(G128), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n243), .A2(G143), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n195), .B2(new_n194), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n196), .A2(new_n455), .A3(new_n456), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT91), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT91), .B1(new_n458), .B2(new_n459), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n454), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n453), .B(new_n225), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT13), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n455), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n456), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n455), .A2(new_n465), .ZN(new_n468));
  OAI21_X1  g282(.A(G134), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n459), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n196), .A2(KEYINPUT90), .A3(new_n455), .A4(new_n456), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n464), .A2(new_n469), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n449), .B1(new_n463), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n463), .A2(new_n449), .A3(new_n473), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G478), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT15), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n476), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n190), .B1(new_n482), .B2(new_n474), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n479), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n447), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n386), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n319), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G472), .ZN(new_n490));
  OR2_X1    g304(.A1(KEYINPUT66), .A2(G134), .ZN(new_n491));
  NAND2_X1  g305(.A1(KEYINPUT66), .A2(G134), .ZN(new_n492));
  AOI21_X1  g306(.A(G137), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n192), .A2(G134), .ZN(new_n494));
  OAI21_X1  g308(.A(G131), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n204), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT69), .B1(new_n263), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT69), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n252), .A2(new_n498), .A3(new_n204), .A4(new_n495), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n285), .B1(new_n205), .B2(new_n206), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n497), .A2(KEYINPUT30), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n197), .A2(new_n202), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G131), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n284), .B1(new_n503), .B2(new_n204), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT67), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n258), .A2(new_n260), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n496), .A2(new_n505), .B1(new_n506), .B2(new_n223), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n204), .A2(KEYINPUT67), .A3(new_n495), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n501), .B(new_n334), .C1(new_n509), .C2(KEYINPUT30), .ZN(new_n510));
  INV_X1    g324(.A(new_n334), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n497), .A2(new_n511), .A3(new_n499), .A4(new_n500), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n402), .A2(G210), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT27), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT26), .B(G101), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n512), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n496), .A2(new_n505), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n252), .A3(new_n508), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n511), .B1(new_n521), .B2(new_n500), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT28), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT71), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n252), .A2(new_n204), .A3(new_n495), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n524), .B1(new_n526), .B2(new_n504), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n500), .A2(KEYINPUT71), .A3(new_n525), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n511), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n523), .A2(new_n531), .A3(new_n517), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n518), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n500), .A2(new_n525), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n334), .B1(new_n535), .B2(new_n524), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT28), .B1(new_n536), .B2(new_n528), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n334), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n512), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n540), .B2(KEYINPUT28), .ZN(new_n541));
  INV_X1    g355(.A(new_n517), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n533), .ZN(new_n543));
  AOI21_X1  g357(.A(G902), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n490), .B1(new_n534), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(G472), .A2(G902), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n508), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT67), .B1(new_n204), .B2(new_n495), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n549), .A2(new_n550), .A3(new_n263), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n334), .B1(new_n551), .B2(new_n504), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n530), .B1(new_n552), .B2(new_n512), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n542), .B1(new_n553), .B2(new_n537), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT72), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n523), .A2(new_n531), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT72), .A3(new_n542), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n513), .A2(KEYINPUT70), .A3(KEYINPUT31), .A4(new_n517), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n510), .A2(KEYINPUT70), .A3(new_n512), .A4(new_n517), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT31), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AOI211_X1 g378(.A(KEYINPUT32), .B(new_n548), .C1(new_n559), .C2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT32), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT72), .B1(new_n557), .B2(new_n542), .ZN(new_n567));
  AOI211_X1 g381(.A(new_n555), .B(new_n517), .C1(new_n523), .C2(new_n531), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n561), .A2(new_n562), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n561), .A2(new_n562), .ZN(new_n570));
  OAI22_X1  g384(.A1(new_n567), .A2(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n566), .B1(new_n571), .B2(new_n547), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n546), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  XOR2_X1   g387(.A(KEYINPUT24), .B(G110), .Z(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT74), .ZN(new_n575));
  XNOR2_X1  g389(.A(G119), .B(G128), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT23), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n324), .B2(G128), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n243), .A2(KEYINPUT23), .A3(G119), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n578), .B(new_n579), .C1(G119), .C2(new_n243), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n575), .A2(new_n576), .B1(G110), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n397), .B2(new_n400), .ZN(new_n582));
  OAI22_X1  g396(.A1(new_n575), .A2(new_n576), .B1(G110), .B2(new_n580), .ZN(new_n583));
  INV_X1    g397(.A(new_n400), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n420), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT22), .B(G137), .ZN(new_n587));
  INV_X1    g401(.A(G234), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n187), .A2(new_n588), .A3(G953), .ZN(new_n589));
  XOR2_X1   g403(.A(new_n587), .B(new_n589), .Z(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n582), .A2(new_n585), .A3(new_n590), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n190), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT25), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(G217), .B1(new_n588), .B2(G902), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT73), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n592), .A2(new_n593), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n598), .A2(G902), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n573), .A2(KEYINPUT76), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT76), .B1(new_n573), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n489), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  AOI21_X1  g421(.A(new_n490), .B1(new_n571), .B2(new_n190), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n556), .A2(new_n558), .B1(new_n560), .B2(new_n563), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n548), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n319), .A2(new_n603), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n477), .B2(G478), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n483), .A2(KEYINPUT94), .A3(new_n478), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT93), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n448), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n475), .B2(new_n476), .ZN(new_n621));
  INV_X1    g435(.A(new_n620), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n482), .A2(new_n474), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n478), .A2(G902), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n617), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n447), .ZN(new_n628));
  INV_X1    g442(.A(new_n375), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n370), .A2(new_n371), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n628), .A2(new_n631), .A3(new_n385), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n613), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT95), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NOR2_X1   g450(.A1(new_n630), .A2(new_n384), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT96), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n445), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n440), .A2(new_n441), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT20), .ZN(new_n641));
  INV_X1    g455(.A(new_n445), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n642), .A3(KEYINPUT96), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n485), .A2(new_n434), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n637), .A2(new_n639), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n613), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT35), .B(G107), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  OR2_X1    g462(.A1(new_n608), .A2(new_n610), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n591), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n586), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n601), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n599), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n489), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  INV_X1    g472(.A(new_n379), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n659), .B1(new_n660), .B2(new_n381), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n644), .A2(new_n643), .A3(new_n639), .A4(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n630), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n573), .A2(new_n319), .A3(new_n653), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  INV_X1    g480(.A(KEYINPUT98), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT97), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT32), .B1(new_n609), .B2(new_n548), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n571), .A2(new_n566), .A3(new_n547), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n513), .A2(new_n517), .ZN(new_n672));
  INV_X1    g486(.A(new_n540), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n672), .B1(new_n517), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n490), .B1(new_n674), .B2(new_n190), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n668), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  AOI211_X1 g491(.A(KEYINPUT97), .B(new_n675), .C1(new_n669), .C2(new_n670), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n667), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n676), .B1(new_n565), .B2(new_n572), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT97), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n671), .A2(new_n668), .A3(new_n676), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(KEYINPUT98), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n661), .B(KEYINPUT39), .Z(new_n685));
  NAND2_X1  g499(.A1(new_n319), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n372), .B(KEYINPUT38), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n375), .B1(new_n481), .B2(new_n484), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n446), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n690), .A2(new_n654), .A3(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n684), .A2(new_n687), .A3(new_n688), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  NAND2_X1  g509(.A1(new_n617), .A2(new_n626), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n696), .A2(new_n446), .A3(new_n662), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT99), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n631), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n696), .A2(new_n446), .A3(new_n662), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT99), .B1(new_n700), .B2(new_n630), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n573), .A2(new_n319), .A3(new_n653), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  NAND2_X1  g518(.A1(new_n299), .A2(new_n303), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n190), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  INV_X1    g521(.A(new_n191), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n705), .A2(new_n305), .A3(new_n190), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n632), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n573), .A2(new_n603), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT100), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n603), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n671), .B2(new_n546), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(KEYINPUT100), .A3(new_n711), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NOR2_X1   g534(.A1(new_n645), .A2(new_n710), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n573), .A3(new_n603), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT101), .B(G116), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G18));
  NOR2_X1   g538(.A1(new_n710), .A2(new_n630), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n487), .A2(new_n384), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n573), .A2(new_n653), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  NAND3_X1  g542(.A1(new_n373), .A2(new_n692), .A3(new_n385), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n710), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n541), .A2(new_n517), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n548), .B1(new_n564), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n571), .A2(new_n190), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n732), .B1(new_n733), .B2(G472), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n730), .A2(new_n734), .A3(KEYINPUT102), .A4(new_n603), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT102), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n569), .A2(new_n570), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n541), .A2(new_n517), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n547), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(G902), .B1(new_n559), .B2(new_n564), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n603), .B(new_n739), .C1(new_n740), .C2(new_n490), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n305), .B1(new_n705), .B2(new_n190), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n304), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n370), .A2(new_n446), .A3(new_n371), .A4(new_n691), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n384), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n745), .A3(new_n708), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n736), .B1(new_n741), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n735), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  NOR4_X1   g563(.A1(new_n608), .A2(new_n654), .A3(new_n732), .A4(new_n700), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n725), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G125), .ZN(G27));
  NOR2_X1   g566(.A1(new_n373), .A2(new_n375), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT103), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(new_n308), .B2(new_n310), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT103), .B1(new_n315), .B2(new_n297), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n756), .A2(new_n305), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n305), .A2(new_n190), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n709), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n708), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT104), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n754), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n308), .A2(new_n755), .ZN(new_n765));
  OAI211_X1 g579(.A(G469), .B(new_n765), .C1(new_n316), .C2(new_n755), .ZN(new_n766));
  AOI21_X1  g580(.A(G902), .B1(new_n299), .B2(new_n303), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n759), .B1(new_n767), .B2(new_n305), .ZN(new_n768));
  AOI211_X1 g582(.A(new_n763), .B(new_n191), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n716), .A2(new_n697), .A3(new_n764), .A4(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  AOI21_X1  g588(.A(new_n191), .B1(new_n766), .B2(new_n768), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n753), .B1(new_n775), .B2(KEYINPUT104), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n769), .ZN(new_n777));
  INV_X1    g591(.A(new_n663), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n716), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  OAI211_X1 g594(.A(KEYINPUT45), .B(new_n765), .C1(new_n316), .C2(new_n755), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n781), .B(G469), .C1(KEYINPUT45), .C2(new_n316), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n760), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n709), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n783), .A2(new_n784), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n708), .B(new_n685), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT106), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n790), .B(KEYINPUT43), .C1(new_n627), .C2(new_n446), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT43), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n627), .A2(new_n446), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n792), .B1(new_n793), .B2(KEYINPUT106), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n649), .A2(new_n653), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n754), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n789), .B(new_n797), .C1(new_n796), .C2(new_n795), .ZN(new_n798));
  XNOR2_X1  g612(.A(KEYINPUT107), .B(G137), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(G39));
  OAI21_X1  g614(.A(new_n708), .B1(new_n786), .B2(new_n787), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT47), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n573), .A2(new_n603), .A3(new_n700), .A4(new_n754), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  NOR2_X1   g622(.A1(G952), .A2(G953), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n754), .A2(new_n710), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n603), .A3(new_n659), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n684), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n447), .A3(new_n627), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n794), .A2(new_n659), .A3(new_n791), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT111), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n794), .A2(new_n816), .A3(new_n659), .A4(new_n791), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n741), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n710), .A2(new_n629), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT112), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n818), .A2(new_n689), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n818), .A2(new_n820), .A3(KEYINPUT50), .A4(new_n689), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n710), .B(new_n754), .C1(new_n815), .C2(new_n817), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n653), .A3(new_n734), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n813), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n743), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n708), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n753), .B(new_n818), .C1(new_n805), .C2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(KEYINPUT51), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n826), .A2(new_n716), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT48), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n812), .A2(new_n628), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n293), .A2(G952), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n818), .B2(new_n725), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n829), .A2(KEYINPUT113), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n828), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n832), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n840), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n665), .A2(new_n703), .A3(new_n751), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n653), .A2(new_n661), .A3(new_n744), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n775), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n681), .B2(new_n682), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n848), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n313), .B(G469), .C1(new_n316), .C2(G902), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n318), .A2(new_n854), .A3(new_n709), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n855), .A2(new_n708), .A3(new_n664), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n654), .B1(new_n671), .B2(new_n546), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n856), .A2(new_n857), .B1(new_n725), .B2(new_n750), .ZN(new_n858));
  INV_X1    g672(.A(new_n851), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(new_n677), .B2(new_n678), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n858), .A2(new_n860), .A3(KEYINPUT52), .A4(new_n703), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n489), .ZN(new_n863));
  INV_X1    g677(.A(new_n605), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n716), .A2(KEYINPUT76), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT108), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n628), .A2(new_n867), .B1(new_n447), .B2(new_n485), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT108), .B1(new_n627), .B2(new_n447), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n386), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n319), .A3(new_n603), .A4(new_n611), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n656), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n727), .A2(new_n722), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n718), .A2(new_n874), .A3(new_n748), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n862), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT109), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n777), .B2(new_n750), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n877), .A2(new_n764), .A3(new_n750), .A4(new_n770), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n643), .A2(new_n639), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n486), .A2(new_n434), .A3(new_n662), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n754), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n857), .A2(new_n319), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n779), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n773), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n847), .B1(new_n876), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n612), .A2(new_n870), .B1(new_n489), .B2(new_n655), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n606), .A3(KEYINPUT53), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n748), .A2(new_n722), .A3(new_n727), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n718), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n891), .B1(new_n893), .B2(KEYINPUT110), .ZN(new_n894));
  INV_X1    g708(.A(new_n772), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n771), .B(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n779), .B(new_n884), .C1(new_n878), .C2(new_n879), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT110), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n892), .A2(new_n899), .A3(new_n718), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n894), .A2(new_n898), .A3(new_n862), .A4(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n888), .A2(new_n889), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n892), .A2(new_n606), .A3(new_n890), .A4(new_n718), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n853), .B2(new_n861), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(KEYINPUT53), .A3(new_n898), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n888), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n902), .B1(new_n906), .B2(KEYINPUT54), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n809), .B1(new_n846), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT114), .ZN(new_n909));
  INV_X1    g723(.A(new_n684), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n830), .A2(KEYINPUT49), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n830), .A2(KEYINPUT49), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n603), .A2(new_n708), .A3(new_n376), .A4(new_n793), .ZN(new_n913));
  NOR4_X1   g727(.A1(new_n911), .A2(new_n912), .A3(new_n690), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  OR3_X1    g730(.A1(new_n908), .A2(new_n909), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n909), .B1(new_n908), .B2(new_n916), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(G75));
  NOR2_X1   g733(.A1(new_n293), .A2(G952), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n190), .B1(new_n888), .B2(new_n901), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT56), .B1(new_n922), .B2(new_n368), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n342), .A2(new_n351), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n349), .ZN(new_n925));
  XNOR2_X1  g739(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n921), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n923), .B2(new_n927), .ZN(G51));
  XOR2_X1   g743(.A(new_n782), .B(KEYINPUT117), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n922), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n705), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n759), .B(KEYINPUT57), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n889), .B1(new_n888), .B2(new_n901), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n902), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT116), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n934), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT53), .B1(new_n904), .B2(new_n898), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n893), .A2(KEYINPUT110), .ZN(new_n941));
  INV_X1    g755(.A(new_n891), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n941), .A2(new_n900), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n886), .A2(new_n862), .A3(new_n773), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT54), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n888), .A2(new_n901), .A3(new_n889), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n939), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(KEYINPUT116), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n932), .B1(new_n938), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT118), .B1(new_n950), .B2(new_n920), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n705), .B1(new_n948), .B2(KEYINPUT116), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n936), .A2(new_n937), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n931), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT118), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n955), .A3(new_n921), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n951), .A2(new_n956), .ZN(G54));
  NAND3_X1  g771(.A1(new_n922), .A2(KEYINPUT58), .A3(G475), .ZN(new_n958));
  INV_X1    g772(.A(new_n440), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n958), .A2(KEYINPUT119), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n921), .B1(new_n958), .B2(new_n959), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT119), .B1(new_n958), .B2(new_n959), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G60));
  INV_X1    g777(.A(new_n624), .ZN(new_n964));
  NAND2_X1  g778(.A1(G478), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT59), .Z(new_n966));
  AOI211_X1 g780(.A(new_n964), .B(new_n966), .C1(new_n946), .C2(new_n947), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n907), .A2(new_n966), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n920), .B(new_n967), .C1(new_n968), .C2(new_n964), .ZN(G63));
  NAND2_X1  g783(.A1(new_n888), .A2(new_n901), .ZN(new_n970));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT60), .Z(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT120), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n970), .A2(KEYINPUT120), .A3(new_n972), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n920), .B1(new_n977), .B2(new_n651), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n600), .B(KEYINPUT121), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n975), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n978), .A2(KEYINPUT61), .A3(new_n980), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(G66));
  INV_X1    g799(.A(G224), .ZN(new_n986));
  OAI21_X1  g800(.A(G953), .B1(new_n382), .B2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n903), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n987), .B1(new_n988), .B2(G953), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n924), .B1(G898), .B2(new_n293), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT122), .Z(new_n991));
  XNOR2_X1  g805(.A(new_n989), .B(new_n991), .ZN(G69));
  OAI21_X1  g806(.A(new_n501), .B1(new_n509), .B2(KEYINPUT30), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT123), .Z(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(new_n437), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n864), .A2(new_n865), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n754), .B1(new_n868), .B2(new_n869), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n996), .A2(new_n319), .A3(new_n685), .A4(new_n997), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n798), .A2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT62), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n849), .B(KEYINPUT124), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n1001), .A2(new_n694), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n999), .B(new_n807), .C1(new_n1000), .C2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n995), .B1(new_n1004), .B2(G953), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n293), .A2(G900), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n798), .A2(new_n1001), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT126), .ZN(new_n1008));
  AOI211_X1 g822(.A(new_n715), .B(new_n744), .C1(new_n671), .C2(new_n546), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n789), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n807), .A2(new_n773), .A3(new_n779), .A4(new_n1010), .ZN(new_n1011));
  OR2_X1    g825(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1006), .B1(new_n1012), .B2(new_n293), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1005), .B1(new_n1013), .B2(new_n995), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n293), .B1(G227), .B2(G900), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1015), .B(KEYINPUT125), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1014), .B(new_n1016), .ZN(G72));
  XNOR2_X1  g831(.A(new_n513), .B(KEYINPUT127), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n1004), .A2(new_n988), .ZN(new_n1019));
  NAND2_X1  g833(.A1(G472), .A2(G902), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT63), .Z(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n517), .B(new_n1018), .C1(new_n1019), .C2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1021), .B1(new_n1012), .B2(new_n903), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1018), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1024), .A2(new_n542), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1022), .B1(new_n518), .B2(new_n672), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n920), .B1(new_n906), .B2(new_n1027), .ZN(new_n1028));
  AND3_X1   g842(.A1(new_n1023), .A2(new_n1026), .A3(new_n1028), .ZN(G57));
endmodule


