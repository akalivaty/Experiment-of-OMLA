//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G77), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT65), .Z(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n203), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT67), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n214), .B(new_n215), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n213), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT68), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n213), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT66), .B(KEYINPUT0), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n202), .A2(new_n203), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(new_n211), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n230), .B(new_n236), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n226), .A2(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT70), .ZN(new_n244));
  XOR2_X1   g0044(.A(G250), .B(G257), .Z(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n211), .A2(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n234), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(KEYINPUT11), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(KEYINPUT11), .ZN(new_n265));
  INV_X1    g0065(.A(new_n262), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n210), .A2(G20), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(G68), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G13), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G20), .A3(new_n203), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT12), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n264), .A2(new_n265), .A3(new_n271), .A4(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT71), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  INV_X1    g0081(.A(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(KEYINPUT71), .A3(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(G226), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(G232), .A3(G1698), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G97), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n234), .B1(G33), .B2(G41), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT13), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  OAI211_X1 g0099(.A(G1), .B(G13), .C1(new_n282), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n295), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n298), .B1(new_n301), .B2(new_n217), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n293), .A2(new_n294), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n294), .B1(new_n293), .B2(new_n303), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n305), .B2(new_n306), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n276), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT14), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT14), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(G169), .C1(new_n306), .C2(new_n305), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n307), .A2(G179), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n312), .B1(new_n318), .B2(new_n276), .ZN(new_n319));
  INV_X1    g0119(.A(G226), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n298), .B1(new_n301), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n286), .A2(G222), .A3(new_n287), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n286), .A2(G1698), .ZN(new_n323));
  INV_X1    g0123(.A(G223), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n322), .B1(new_n258), .B2(new_n286), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n321), .B1(new_n325), .B2(new_n292), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G179), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n313), .B2(new_n326), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n205), .A2(G20), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT8), .B(G58), .ZN(new_n330));
  INV_X1    g0130(.A(G150), .ZN(new_n331));
  INV_X1    g0131(.A(new_n256), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n330), .A2(new_n259), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n262), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n270), .A2(G50), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n268), .A2(new_n335), .B1(G50), .B2(new_n267), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n328), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  XOR2_X1   g0140(.A(new_n338), .B(KEYINPUT9), .Z(new_n341));
  NOR2_X1   g0141(.A1(new_n326), .A2(new_n310), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n326), .A2(G190), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT10), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT10), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n343), .A2(new_n347), .A3(new_n344), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n340), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n283), .A2(new_n284), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G226), .A2(G1698), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n324), .B2(G1698), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n350), .A2(new_n352), .B1(G33), .B2(G87), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(new_n300), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT75), .ZN(new_n355));
  INV_X1    g0155(.A(G232), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n298), .B1(new_n301), .B2(new_n356), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n355), .A2(G179), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n354), .A2(new_n357), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(G169), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n330), .B1(new_n210), .B2(G20), .ZN(new_n362));
  INV_X1    g0162(.A(new_n267), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n269), .A2(new_n362), .B1(new_n363), .B2(new_n330), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n350), .A2(new_n365), .A3(G20), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n350), .B2(G20), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G68), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G58), .A2(G68), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n231), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G20), .ZN(new_n373));
  INV_X1    g0173(.A(G159), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n373), .A2(KEYINPUT73), .B1(new_n374), .B2(new_n332), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n373), .A2(KEYINPUT73), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n370), .A2(KEYINPUT16), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n262), .ZN(new_n379));
  XOR2_X1   g0179(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(G20), .B1(new_n280), .B2(new_n285), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n367), .B1(new_n382), .B2(KEYINPUT7), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G68), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n381), .B1(new_n384), .B2(new_n377), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n364), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n361), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT18), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n357), .A2(G190), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n355), .A2(new_n389), .B1(G200), .B2(new_n359), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n390), .B(new_n364), .C1(new_n385), .C2(new_n379), .ZN(new_n391));
  XOR2_X1   g0191(.A(new_n391), .B(KEYINPUT17), .Z(new_n392));
  NOR2_X1   g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n394), .A2(new_n259), .B1(new_n211), .B2(new_n258), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n330), .A2(new_n332), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n262), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n397), .B(KEYINPUT72), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n267), .A2(G77), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n269), .A2(G77), .A3(new_n270), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G244), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n298), .B1(new_n301), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n286), .A2(G232), .A3(new_n287), .ZN(new_n404));
  INV_X1    g0204(.A(G107), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n404), .B1(new_n405), .B2(new_n286), .C1(new_n323), .C2(new_n217), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n403), .B1(new_n406), .B2(new_n292), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n407), .A2(new_n308), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(G200), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n401), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n401), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n407), .A2(new_n313), .ZN(new_n412));
  INV_X1    g0212(.A(G179), .ZN(new_n413));
  AOI211_X1 g0213(.A(new_n413), .B(new_n403), .C1(new_n406), .C2(new_n292), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n411), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  AND4_X1   g0216(.A1(new_n319), .A2(new_n349), .A3(new_n393), .A4(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT79), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G283), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(G244), .B(new_n287), .C1(new_n278), .C2(new_n279), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT4), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n422), .A2(new_n402), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n280), .A2(new_n285), .A3(new_n287), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n286), .A2(KEYINPUT76), .A3(G250), .A4(G1698), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n280), .A2(new_n285), .A3(G250), .A4(G1698), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT76), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n426), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT77), .B1(new_n431), .B2(new_n300), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT77), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n428), .B(KEYINPUT76), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n433), .B(new_n292), .C1(new_n434), .C2(new_n426), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n210), .A2(G45), .ZN(new_n436));
  NAND2_X1  g0236(.A1(KEYINPUT5), .A2(G41), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(KEYINPUT5), .A2(G41), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(G257), .A3(new_n300), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT78), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n210), .A2(G45), .ZN(new_n443));
  INV_X1    g0243(.A(new_n439), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(new_n437), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G274), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n441), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n442), .B1(new_n441), .B2(new_n446), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AND4_X1   g0249(.A1(new_n413), .A2(new_n432), .A3(new_n435), .A4(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n267), .A2(G97), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n210), .A2(G33), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n267), .A2(new_n452), .A3(new_n234), .A4(new_n261), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n451), .B1(new_n454), .B2(G97), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT6), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n456), .A2(new_n457), .A3(G107), .ZN(new_n458));
  XNOR2_X1  g0258(.A(G97), .B(G107), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n458), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  OAI22_X1  g0260(.A1(new_n460), .A2(new_n211), .B1(new_n258), .B2(new_n332), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n383), .B2(G107), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n455), .B1(new_n462), .B2(new_n266), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n441), .A2(new_n446), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT78), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n441), .A2(new_n442), .A3(new_n446), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n428), .A2(new_n429), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n428), .A2(new_n429), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n425), .B(new_n423), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n467), .B1(new_n470), .B2(new_n292), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n463), .B1(new_n471), .B2(G169), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n418), .B1(new_n450), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n449), .B1(new_n431), .B2(new_n300), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n459), .A2(new_n456), .ZN(new_n475));
  INV_X1    g0275(.A(new_n458), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n477), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n278), .A2(new_n279), .A3(new_n277), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT71), .B1(new_n283), .B2(new_n284), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n211), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n366), .B1(new_n481), .B2(new_n365), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n478), .B1(new_n482), .B2(new_n405), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n262), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n313), .A2(new_n474), .B1(new_n484), .B2(new_n455), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n432), .A2(new_n435), .A3(new_n413), .A4(new_n449), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(KEYINPUT79), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n432), .A2(new_n435), .A3(new_n449), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G200), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n463), .B1(new_n471), .B2(G190), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n473), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n211), .A2(G107), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT25), .B1(new_n273), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT83), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n273), .A2(new_n494), .A3(KEYINPUT25), .ZN(new_n498));
  OR2_X1    g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(KEYINPUT83), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n499), .A2(new_n500), .B1(G107), .B2(new_n454), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n350), .A2(new_n211), .A3(G87), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT22), .ZN(new_n503));
  INV_X1    g0303(.A(G87), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n504), .A2(KEYINPUT22), .A3(G20), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n280), .A2(new_n285), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n494), .A2(KEYINPUT23), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n494), .A2(KEYINPUT23), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G116), .ZN(new_n510));
  OR3_X1    g0310(.A1(new_n510), .A2(KEYINPUT82), .A3(G20), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT82), .B1(new_n510), .B2(G20), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n508), .A2(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n507), .A2(KEYINPUT24), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n262), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT24), .B1(new_n507), .B2(new_n513), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n501), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(G257), .A2(G1698), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n278), .B2(new_n279), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT84), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(KEYINPUT84), .B(new_n519), .C1(new_n278), .C2(new_n279), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(G250), .B(new_n287), .C1(new_n278), .C2(new_n279), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G294), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT85), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n292), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n524), .B2(new_n527), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT86), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n524), .A2(new_n527), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT85), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT86), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n534), .A2(new_n535), .A3(new_n292), .A4(new_n529), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n445), .A2(new_n292), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G264), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n538), .A2(new_n446), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n532), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G169), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n446), .B(new_n538), .C1(new_n530), .C2(new_n531), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G179), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n518), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n443), .A2(G250), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT80), .B1(new_n292), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT80), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n300), .A2(new_n548), .A3(G250), .A4(new_n443), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n547), .A2(new_n549), .B1(G274), .B2(new_n436), .ZN(new_n550));
  OAI211_X1 g0350(.A(G238), .B(new_n287), .C1(new_n278), .C2(new_n279), .ZN(new_n551));
  OAI211_X1 g0351(.A(G244), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(new_n510), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n292), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(new_n308), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n211), .B1(new_n290), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n504), .A2(new_n457), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(G107), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n211), .B(G68), .C1(new_n278), .C2(new_n279), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n557), .B1(new_n290), .B2(G20), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n262), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n394), .A2(new_n363), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT81), .B1(new_n453), .B2(new_n504), .ZN(new_n566));
  OR3_X1    g0366(.A1(new_n453), .A2(KEYINPUT81), .A3(new_n504), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n564), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n310), .B1(new_n550), .B2(new_n554), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n556), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n555), .A2(G169), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n550), .A2(G179), .A3(new_n554), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n564), .A2(new_n565), .ZN(new_n573));
  INV_X1    g0373(.A(new_n394), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n454), .A2(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n571), .A2(new_n572), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n537), .A2(G270), .B1(G274), .B2(new_n445), .ZN(new_n578));
  INV_X1    g0378(.A(G303), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n280), .B2(new_n285), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G264), .A2(G1698), .ZN(new_n581));
  INV_X1    g0381(.A(G257), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n582), .B2(G1698), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n350), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n292), .B1(new_n580), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n310), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(G190), .B2(new_n587), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n282), .A2(G97), .ZN(new_n590));
  AOI21_X1  g0390(.A(G20), .B1(new_n590), .B2(new_n419), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n211), .A2(new_n218), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n262), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT20), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(KEYINPUT20), .B(new_n262), .C1(new_n591), .C2(new_n592), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n267), .A2(new_n218), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n454), .B2(new_n218), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n589), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n280), .A2(new_n285), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G303), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n300), .B1(new_n602), .B2(new_n584), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n440), .A2(new_n300), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n446), .B1(new_n604), .B2(new_n219), .ZN(new_n605));
  OAI211_X1 g0405(.A(KEYINPUT21), .B(G169), .C1(new_n603), .C2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n578), .A2(new_n586), .A3(G179), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n597), .A2(new_n599), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n587), .A3(G169), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n608), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n577), .A2(new_n600), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n532), .A2(new_n536), .A3(new_n308), .A4(new_n539), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n542), .A2(new_n310), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n517), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n545), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n417), .A2(new_n493), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g0418(.A(new_n618), .B(KEYINPUT87), .Z(G372));
  AND3_X1   g0419(.A1(new_n485), .A2(KEYINPUT79), .A3(new_n486), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT79), .B1(new_n485), .B2(new_n486), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n540), .A2(G169), .B1(new_n543), .B2(G179), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n623), .A2(new_n518), .B1(new_n616), .B2(new_n612), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n622), .A2(new_n491), .A3(new_n624), .A4(new_n577), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n577), .B1(new_n620), .B2(new_n621), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT26), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n577), .A2(new_n485), .A3(new_n628), .A4(new_n486), .ZN(new_n629));
  INV_X1    g0429(.A(new_n576), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n625), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n417), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT88), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT88), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT18), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n387), .B(new_n636), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n392), .A2(new_n312), .ZN(new_n638));
  INV_X1    g0438(.A(new_n415), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n318), .B2(new_n276), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n346), .A2(new_n348), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n340), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n634), .A2(new_n635), .A3(new_n643), .ZN(G369));
  NAND2_X1  g0444(.A1(new_n600), .A2(new_n612), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n273), .A2(new_n211), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n649), .B(KEYINPUT89), .Z(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n609), .ZN(new_n654));
  MUX2_X1   g0454(.A(new_n612), .B(new_n645), .S(new_n654), .Z(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g0456(.A(KEYINPUT90), .B(G330), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT91), .ZN(new_n660));
  INV_X1    g0460(.A(new_n545), .ZN(new_n661));
  INV_X1    g0461(.A(new_n616), .ZN(new_n662));
  INV_X1    g0462(.A(new_n653), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n661), .B(new_n662), .C1(new_n518), .C2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n545), .A2(new_n653), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n653), .A2(new_n612), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n545), .B2(new_n663), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(G399));
  INV_X1    g0473(.A(new_n227), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT92), .B1(new_n676), .B2(new_n232), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n559), .A2(G107), .A3(G116), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(G1), .A3(new_n678), .ZN(new_n679));
  MUX2_X1   g0479(.A(KEYINPUT92), .B(new_n677), .S(new_n679), .Z(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT93), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n614), .A2(new_n615), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n612), .B1(new_n683), .B2(new_n518), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n577), .B1(new_n684), .B2(new_n545), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n492), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n450), .A2(new_n472), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n628), .B1(new_n687), .B2(new_n577), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n686), .A2(new_n576), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(KEYINPUT26), .B2(new_n626), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(KEYINPUT29), .A3(new_n663), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n632), .A2(new_n663), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n530), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n534), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n607), .A2(new_n555), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n471), .A2(new_n697), .A3(new_n538), .A4(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n587), .A2(new_n413), .A3(new_n555), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n488), .A2(new_n542), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n700), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n653), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  XOR2_X1   g0507(.A(KEYINPUT94), .B(KEYINPUT31), .Z(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(KEYINPUT31), .B2(new_n707), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n493), .A2(new_n617), .A3(new_n663), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n658), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n695), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n682), .B1(new_n716), .B2(G1), .ZN(G364));
  NOR2_X1   g0517(.A1(new_n272), .A2(G20), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G45), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT95), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(KEYINPUT95), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n675), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n656), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n211), .A2(G190), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n310), .A2(G179), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n405), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n211), .A2(new_n308), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n413), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n202), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n413), .A2(new_n310), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n735), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI211_X1 g0541(.A(new_n734), .B(new_n738), .C1(G50), .C2(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(KEYINPUT96), .B(G159), .Z(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n731), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT32), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n735), .A2(new_n732), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n748), .A2(KEYINPUT97), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(KEYINPUT97), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n742), .B(new_n747), .C1(new_n504), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n739), .A2(new_n731), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n731), .A2(new_n736), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G68), .A2(new_n754), .B1(new_n756), .B2(G77), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n744), .A2(G190), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G97), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n757), .A2(new_n286), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT33), .B(G317), .ZN(new_n762));
  INV_X1    g0562(.A(new_n745), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n754), .A2(new_n762), .B1(new_n763), .B2(G329), .ZN(new_n764));
  INV_X1    g0564(.A(G294), .ZN(new_n765));
  INV_X1    g0565(.A(new_n759), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n764), .B(new_n601), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n741), .A2(G326), .B1(new_n756), .B2(G311), .ZN(new_n768));
  INV_X1    g0568(.A(new_n737), .ZN(new_n769));
  INV_X1    g0569(.A(new_n733), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G322), .A2(new_n769), .B1(new_n770), .B2(G283), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n768), .B(new_n771), .C1(new_n751), .C2(new_n579), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n752), .A2(new_n761), .B1(new_n767), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n234), .B1(G20), .B2(new_n313), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n674), .A2(new_n218), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n286), .A2(new_n227), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n233), .A2(G45), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n251), .B2(G45), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n674), .A2(new_n350), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n775), .B1(new_n208), .B2(new_n776), .C1(new_n778), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n727), .A2(new_n774), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n773), .A2(new_n774), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n724), .B1(new_n730), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n660), .B1(new_n656), .B2(new_n658), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(new_n785), .B2(new_n724), .ZN(G396));
  OAI21_X1  g0586(.A(KEYINPUT98), .B1(new_n415), .B2(new_n663), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n407), .A2(G179), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n313), .B2(new_n407), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT98), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n789), .A2(new_n790), .A3(new_n411), .A4(new_n653), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n410), .B(new_n415), .C1(new_n401), .C2(new_n663), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT99), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n692), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT100), .Z(new_n797));
  INV_X1    g0597(.A(new_n577), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(new_n473), .B2(new_n487), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n631), .B1(new_n799), .B2(new_n628), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n663), .B(new_n794), .C1(new_n800), .C2(new_n686), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT101), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n632), .A2(KEYINPUT101), .A3(new_n663), .A4(new_n794), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n797), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n714), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n724), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n807), .A2(KEYINPUT102), .A3(new_n714), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(KEYINPUT102), .B1(new_n807), .B2(new_n714), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n774), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n726), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n723), .B1(G77), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n733), .A2(new_n504), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n737), .A2(new_n765), .B1(new_n745), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n817), .B(new_n819), .C1(G116), .C2(new_n756), .ZN(new_n820));
  INV_X1    g0620(.A(new_n751), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G107), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n740), .A2(new_n579), .B1(new_n753), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n286), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n820), .A2(new_n822), .A3(new_n760), .A4(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G143), .A2(new_n769), .B1(new_n754), .B2(G150), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n828), .B2(new_n740), .C1(new_n755), .C2(new_n743), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT34), .Z(new_n830));
  NAND2_X1  g0630(.A1(new_n770), .A2(G68), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n831), .B(new_n350), .C1(new_n832), .C2(new_n745), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G58), .B2(new_n759), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n201), .B2(new_n751), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n826), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n816), .B1(new_n836), .B2(new_n774), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n794), .B2(new_n726), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n813), .A2(new_n838), .ZN(G384));
  INV_X1    g0639(.A(new_n276), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n663), .A2(new_n840), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n841), .B(new_n312), .C1(new_n318), .C2(new_n276), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n276), .B(new_n653), .C1(new_n318), .C2(new_n312), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n377), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n203), .B1(new_n367), .B2(new_n368), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n380), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT105), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(new_n850), .A3(new_n262), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n381), .B1(new_n370), .B2(new_n377), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT105), .B1(new_n852), .B2(new_n266), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n853), .A3(new_n378), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n651), .B1(new_n854), .B2(new_n364), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n388), .B2(new_n392), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  INV_X1    g0657(.A(new_n391), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n854), .A2(new_n364), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n361), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n857), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n386), .A2(new_n650), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n387), .A2(new_n863), .A3(new_n391), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n856), .B(KEYINPUT38), .C1(new_n862), .C2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n860), .A2(new_n650), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n861), .A2(new_n868), .A3(new_n391), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n865), .B1(new_n869), .B2(KEYINPUT37), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n391), .B(KEYINPUT17), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n868), .B1(new_n637), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n867), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT104), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n639), .A2(new_n663), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n805), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n876), .ZN(new_n878));
  AOI211_X1 g0678(.A(KEYINPUT104), .B(new_n878), .C1(new_n803), .C2(new_n804), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n846), .B(new_n874), .C1(new_n877), .C2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n388), .A2(new_n651), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n880), .A2(KEYINPUT106), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT106), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n857), .B1(new_n863), .B2(KEYINPUT107), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(new_n864), .Z(new_n886));
  AOI21_X1  g0686(.A(new_n863), .B1(new_n637), .B2(new_n871), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n867), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n866), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n884), .B1(KEYINPUT39), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n318), .A2(new_n276), .A3(new_n663), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n882), .A2(new_n883), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT109), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n695), .A2(new_n417), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n643), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT108), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n896), .B(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n653), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(KEYINPUT111), .Z(new_n902));
  AOI21_X1  g0702(.A(new_n707), .B1(new_n712), .B2(new_n709), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n841), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n319), .A2(new_n906), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n907), .A2(new_n843), .B1(new_n792), .B2(new_n793), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n905), .A2(new_n874), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n901), .B(KEYINPUT111), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(new_n903), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n794), .B1(new_n842), .B2(new_n844), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n888), .B2(new_n866), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n909), .A2(new_n910), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n905), .A2(new_n417), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n917), .B(new_n918), .Z(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(new_n657), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n900), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n900), .A2(new_n920), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n921), .B(new_n922), .C1(new_n210), .C2(new_n718), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n477), .A2(KEYINPUT35), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G116), .A3(new_n235), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(KEYINPUT35), .B2(new_n477), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n926), .A2(KEYINPUT36), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(KEYINPUT36), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n371), .A2(G77), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n232), .A2(new_n929), .B1(G50), .B2(new_n203), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(G1), .A3(new_n272), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT103), .Z(new_n933));
  NAND2_X1  g0733(.A1(new_n923), .A2(new_n933), .ZN(G367));
  NAND2_X1  g0734(.A1(new_n653), .A2(new_n463), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n493), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n687), .A2(new_n653), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n671), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT112), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT42), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n621), .B(new_n620), .C1(new_n938), .C2(new_n545), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n942), .B(new_n943), .C1(new_n653), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n653), .A2(new_n568), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n798), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n576), .B2(new_n946), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT43), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n949), .B2(new_n948), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n948), .A2(new_n949), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n945), .B2(new_n950), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(new_n668), .A3(new_n938), .ZN(new_n956));
  INV_X1    g0756(.A(new_n938), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n952), .A2(new_n954), .B1(new_n669), .B2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n675), .B(KEYINPUT41), .Z(new_n959));
  NOR2_X1   g0759(.A1(new_n672), .A2(new_n938), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT44), .Z(new_n961));
  NAND2_X1  g0761(.A1(new_n672), .A2(new_n938), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT45), .ZN(new_n963));
  OR3_X1    g0763(.A1(new_n961), .A2(new_n668), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n668), .B1(new_n961), .B2(new_n963), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n667), .A2(new_n670), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n664), .B2(new_n670), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n660), .B(new_n969), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n970), .A2(new_n695), .A3(new_n715), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(KEYINPUT113), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(KEYINPUT113), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n967), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n959), .B1(new_n975), .B2(new_n716), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n956), .B(new_n958), .C1(new_n976), .C2(new_n722), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n948), .A2(new_n727), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n782), .B1(new_n227), .B2(new_n394), .ZN(new_n979));
  INV_X1    g0779(.A(new_n247), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n979), .B1(new_n980), .B2(new_n779), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n724), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n733), .A2(new_n258), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n743), .A2(new_n753), .B1(new_n755), .B2(new_n201), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(G137), .C2(new_n763), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n766), .A2(new_n203), .ZN(new_n986));
  INV_X1    g0786(.A(G143), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n740), .A2(new_n987), .B1(new_n737), .B2(new_n331), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n986), .A2(new_n988), .A3(new_n601), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n985), .B(new_n989), .C1(new_n202), .C2(new_n751), .ZN(new_n990));
  INV_X1    g0790(.A(new_n350), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n740), .B2(new_n818), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n737), .A2(new_n579), .B1(new_n733), .B2(new_n457), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(G107), .C2(new_n759), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n821), .A2(KEYINPUT46), .A3(G116), .ZN(new_n995));
  INV_X1    g0795(.A(G317), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n755), .A2(new_n823), .B1(new_n745), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G294), .B2(new_n754), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n751), .B2(new_n218), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n994), .A2(new_n995), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT47), .B1(new_n990), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n990), .A2(new_n1001), .A3(KEYINPUT47), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n774), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n978), .B(new_n982), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n977), .A2(new_n1005), .ZN(G387));
  INV_X1    g0806(.A(new_n970), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n722), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n674), .A2(new_n405), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n243), .A2(G45), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n330), .B2(G50), .ZN(new_n1012));
  AOI21_X1  g0812(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n678), .A3(new_n1013), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n330), .A2(new_n1011), .A3(G50), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n779), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1009), .B1(new_n678), .B2(new_n776), .C1(new_n1010), .C2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n724), .B1(new_n1017), .B2(new_n782), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n574), .A2(new_n759), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n201), .A2(new_n737), .B1(new_n753), .B2(new_n330), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n991), .B(new_n1020), .C1(G97), .C2(new_n770), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n821), .A2(G77), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n755), .A2(new_n203), .B1(new_n745), .B2(new_n331), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G159), .B2(new_n741), .ZN(new_n1024));
  AND4_X1   g0824(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n737), .A2(new_n996), .B1(new_n755), .B2(new_n579), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1026), .A2(KEYINPUT115), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(KEYINPUT115), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G322), .A2(new_n741), .B1(new_n754), .B2(G311), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n821), .A2(G294), .B1(G283), .B2(new_n759), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(G326), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n991), .B1(new_n745), .B2(new_n1038), .C1(new_n218), .C2(new_n733), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1025), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1018), .B1(new_n814), .B2(new_n1041), .C1(new_n666), .C2(new_n728), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n973), .A2(new_n974), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n675), .B1(new_n1007), .B2(new_n716), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1008), .B(new_n1042), .C1(new_n1044), .C2(new_n1045), .ZN(G393));
  NAND2_X1  g0846(.A1(new_n967), .A2(new_n722), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n782), .B1(new_n457), .B2(new_n227), .C1(new_n780), .C2(new_n254), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n723), .ZN(new_n1049));
  INV_X1    g0849(.A(G322), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n755), .A2(new_n765), .B1(new_n745), .B2(new_n1050), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n734), .B(new_n1051), .C1(G303), .C2(new_n754), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n740), .A2(new_n996), .B1(new_n737), .B2(new_n818), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT52), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n821), .A2(G283), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n286), .B1(G116), .B2(new_n759), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n759), .A2(G77), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n201), .B2(new_n753), .C1(new_n330), .C2(new_n755), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT118), .Z(new_n1060));
  OAI22_X1  g0860(.A1(new_n740), .A2(new_n331), .B1(new_n737), .B2(new_n374), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT51), .Z(new_n1062));
  OR4_X1    g0862(.A1(new_n991), .A2(new_n1060), .A3(new_n817), .A4(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n751), .A2(new_n203), .B1(new_n987), .B2(new_n745), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT117), .Z(new_n1065));
  OAI21_X1  g0865(.A(new_n1057), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1049), .B1(new_n1066), .B2(new_n774), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n938), .B2(new_n728), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1047), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n676), .B1(new_n1044), .B2(new_n967), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1043), .A2(new_n966), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(G390));
  NAND3_X1  g0873(.A1(new_n690), .A2(new_n663), .A3(new_n794), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1074), .A2(new_n876), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n891), .B(new_n889), .C1(new_n1075), .C2(new_n845), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n715), .A2(new_n908), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n805), .A2(new_n876), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(KEYINPUT104), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n805), .A2(new_n875), .A3(new_n876), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n892), .B1(new_n1081), .B2(new_n846), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1076), .B(new_n1077), .C1(new_n1082), .C2(new_n890), .ZN(new_n1083));
  INV_X1    g0883(.A(G330), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n912), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n908), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n846), .B1(new_n877), .B2(new_n879), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n890), .B1(new_n1088), .B2(new_n891), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1076), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1083), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n905), .A2(G330), .A3(new_n417), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n897), .A2(new_n643), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n846), .B1(new_n715), .B2(new_n794), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1081), .B1(new_n1087), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1085), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n845), .B1(new_n1097), .B2(new_n795), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1098), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1094), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1092), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1083), .A2(new_n1091), .A3(new_n1100), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n675), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1083), .A2(new_n1091), .A3(new_n722), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n330), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n723), .B1(new_n1106), .B2(new_n815), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n751), .A2(new_n331), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT53), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n763), .A2(G125), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n286), .B(new_n1110), .C1(new_n201), .C2(new_n733), .ZN(new_n1111));
  INV_X1    g0911(.A(G128), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n740), .A2(new_n1112), .B1(new_n737), .B2(new_n832), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT54), .B(G143), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n753), .A2(new_n828), .B1(new_n755), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n766), .A2(new_n374), .ZN(new_n1116));
  NOR4_X1   g0916(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n737), .A2(new_n218), .B1(new_n755), .B2(new_n457), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n740), .A2(new_n823), .B1(new_n753), .B2(new_n405), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1118), .B(new_n1119), .C1(new_n821), .C2(G87), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n763), .A2(G294), .ZN(new_n1121));
  AND4_X1   g0921(.A1(new_n601), .A2(new_n831), .A3(new_n1121), .A4(new_n1058), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1109), .A2(new_n1117), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1123), .A2(KEYINPUT119), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n814), .B1(new_n1123), .B2(KEYINPUT119), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1107), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n890), .B2(new_n726), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1104), .A2(new_n1105), .A3(new_n1127), .ZN(G378));
  INV_X1    g0928(.A(KEYINPUT121), .ZN(new_n1129));
  XOR2_X1   g0929(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1130));
  NAND2_X1  g0930(.A1(new_n650), .A2(new_n338), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n349), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n349), .A2(new_n1131), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1134), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1130), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n1132), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n917), .B2(G330), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n908), .B1(new_n903), .B2(new_n911), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n866), .A2(new_n873), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n910), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n914), .A2(new_n916), .ZN(new_n1144));
  AND4_X1   g0944(.A1(G330), .A2(new_n1143), .A3(new_n1144), .A4(new_n1139), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1129), .B1(new_n895), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n880), .A2(new_n881), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT106), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n880), .A2(KEYINPUT106), .A3(new_n881), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1150), .A2(new_n1151), .A3(new_n893), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1146), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(KEYINPUT121), .A3(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1146), .A2(new_n1150), .A3(new_n1151), .A4(new_n893), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT122), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n883), .A2(new_n894), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1158), .A2(KEYINPUT122), .A3(new_n1151), .A4(new_n1146), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1147), .A2(new_n1154), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1094), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1103), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT57), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1155), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n1162), .A3(KEYINPUT57), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n675), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n723), .B1(G50), .B2(new_n815), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1139), .A2(new_n726), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G128), .A2(new_n769), .B1(new_n756), .B2(G137), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n832), .B2(new_n753), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n741), .A2(G125), .B1(new_n759), .B2(G150), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT120), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1114), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1172), .B(new_n1174), .C1(new_n821), .C2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT59), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n763), .A2(G124), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n743), .A2(new_n733), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1181), .A2(G33), .A3(G41), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n574), .A2(new_n756), .B1(new_n770), .B2(G58), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1022), .B(new_n1184), .C1(new_n823), .C2(new_n745), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n991), .B(new_n299), .C1(new_n457), .C2(new_n753), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n740), .A2(new_n218), .B1(new_n737), .B2(new_n405), .ZN(new_n1187));
  NOR4_X1   g0987(.A1(new_n1185), .A2(new_n986), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1188), .A2(KEYINPUT58), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(KEYINPUT58), .ZN(new_n1190));
  AOI21_X1  g0990(.A(G50), .B1(new_n282), .B2(new_n299), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n350), .B2(G41), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1183), .A2(new_n1189), .A3(new_n1190), .A4(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1169), .B(new_n1170), .C1(new_n774), .C2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1160), .B2(new_n722), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1168), .A2(new_n1195), .ZN(G375));
  NAND2_X1  g0996(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n722), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n723), .B1(G68), .B2(new_n815), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n754), .A2(new_n1175), .B1(new_n763), .B2(G128), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n331), .B2(new_n755), .C1(new_n751), .C2(new_n374), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G132), .A2(new_n741), .B1(new_n769), .B2(G137), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n991), .B1(new_n770), .B2(G58), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(new_n201), .C2(new_n766), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G294), .A2(new_n741), .B1(new_n754), .B2(G116), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G283), .A2(new_n769), .B1(new_n763), .B2(G303), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(new_n751), .C2(new_n457), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n983), .B1(G107), .B2(new_n756), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(new_n601), .A3(new_n1019), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n1201), .A2(new_n1204), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1199), .B1(new_n1210), .B2(new_n774), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT123), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n846), .B2(new_n726), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1198), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n959), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1096), .A2(new_n1099), .A3(new_n1094), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1101), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n1218), .ZN(G381));
  INV_X1    g1019(.A(G375), .ZN(new_n1220));
  INV_X1    g1020(.A(G378), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n977), .A2(new_n1072), .A3(new_n1005), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(G393), .A2(G396), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1226), .A2(G384), .A3(G381), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n1225), .A3(new_n1227), .ZN(G407));
  OAI211_X1 g1028(.A(G407), .B(G213), .C1(G343), .C2(new_n1222), .ZN(G409));
  AND2_X1   g1029(.A1(new_n1217), .A2(KEYINPUT60), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1217), .A2(KEYINPUT60), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n675), .B(new_n1101), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(G384), .A2(new_n1215), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1215), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n838), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n811), .B2(new_n812), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n652), .A2(G213), .A3(G2897), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1240), .A2(KEYINPUT125), .A3(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT125), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n652), .A2(G213), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1160), .A2(new_n1216), .A3(new_n1162), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1194), .B1(new_n1165), .B2(new_n722), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1221), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G378), .B(new_n1195), .C1(new_n1163), .C2(new_n1167), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1249), .A2(new_n1250), .A3(KEYINPUT124), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT124), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1245), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1244), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G393), .A2(G396), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1072), .B1(new_n977), .B2(new_n1005), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1226), .B(new_n1255), .C1(new_n1225), .C2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1256), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1226), .A2(new_n1255), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1224), .A3(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1257), .A2(new_n1258), .A3(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1249), .A2(new_n1250), .B1(G213), .B2(new_n652), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1238), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1262), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1238), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1245), .B(new_n1267), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1264), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1254), .A2(new_n1266), .A3(new_n1269), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1258), .B1(new_n1271), .B2(new_n1263), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT62), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1268), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1263), .A2(KEYINPUT62), .A3(new_n1267), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1272), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(KEYINPUT126), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1270), .B1(new_n1276), .B2(new_n1278), .ZN(G405));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1238), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1257), .A2(new_n1267), .A3(new_n1261), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1282), .B1(new_n1283), .B2(new_n1223), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1223), .A2(new_n1283), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(G402));
endmodule


