//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G57), .Z(G237));
  XOR2_X1   g015(.A(KEYINPUT68), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT69), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g025(.A1(G221), .A2(G218), .A3(G219), .A4(G220), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(G2106), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n460), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(G100), .A2(G2105), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT70), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n465), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n464), .A2(new_n475), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(G162));
  NAND4_X1  g055(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n475), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT4), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT3), .B(G2104), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n483), .A2(new_n484), .A3(G138), .A4(new_n475), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n461), .A2(new_n463), .A3(G126), .A4(G2105), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n486), .A2(KEYINPUT71), .A3(new_n490), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(G164));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G543), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(new_n499), .A3(G62), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT73), .ZN(new_n501));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n497), .A2(new_n499), .A3(new_n503), .A4(G62), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT74), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT72), .A3(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(G543), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n513), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(G50), .A2(new_n516), .B1(new_n519), .B2(G88), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n505), .A2(new_n521), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n507), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(G166));
  AOI22_X1  g099(.A1(new_n510), .A2(new_n512), .B1(KEYINPUT6), .B2(new_n509), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(G51), .A3(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(G89), .A3(new_n517), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  AND4_X1   g105(.A1(new_n526), .A2(new_n527), .A3(new_n528), .A4(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(new_n509), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n525), .A2(G52), .A3(G543), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n525), .A2(G90), .A3(new_n517), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n536), .B1(new_n534), .B2(new_n535), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n533), .B1(new_n537), .B2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n497), .A2(new_n499), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n525), .A2(G81), .A3(new_n517), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n545), .B(new_n546), .C1(new_n547), .C2(new_n515), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  INV_X1    g130(.A(G91), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n518), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n525), .A2(KEYINPUT76), .A3(new_n517), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n517), .A2(G65), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n509), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n525), .A2(G53), .A3(G543), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(G299));
  NAND4_X1  g142(.A1(new_n526), .A2(new_n527), .A3(new_n528), .A4(new_n530), .ZN(G286));
  AND3_X1   g143(.A1(new_n505), .A2(new_n521), .A3(G651), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n521), .B1(new_n505), .B2(G651), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n571), .A2(new_n572), .A3(new_n520), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n523), .A2(KEYINPUT77), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G303));
  NAND2_X1  g150(.A1(new_n558), .A2(new_n559), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n516), .A2(G49), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  AND3_X1   g155(.A1(new_n525), .A2(KEYINPUT76), .A3(new_n517), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT76), .B1(new_n525), .B2(new_n517), .ZN(new_n582));
  OAI21_X1  g157(.A(G86), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT78), .B1(new_n584), .B2(new_n509), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n542), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n588), .A2(new_n589), .A3(G651), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n516), .A2(G48), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n583), .A2(new_n591), .A3(new_n592), .ZN(G305));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n594), .A2(new_n515), .B1(new_n518), .B2(new_n595), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(KEYINPUT79), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(KEYINPUT79), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n542), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n576), .A2(G92), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n542), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n516), .A2(G54), .B1(G651), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n576), .A2(new_n612), .A3(G92), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n607), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n605), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n605), .B1(new_n614), .B2(G868), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT80), .B1(G168), .B2(new_n617), .ZN(new_n618));
  OR3_X1    g193(.A1(G168), .A2(KEYINPUT80), .A3(new_n617), .ZN(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(G868), .ZN(G297));
  OAI211_X1 g196(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n614), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n614), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n483), .A2(new_n466), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n478), .A2(G123), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n465), .A2(G135), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n475), .A2(G111), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n632), .A2(new_n638), .ZN(G156));
  XOR2_X1   g214(.A(KEYINPUT15), .B(G2435), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2438), .ZN(new_n641));
  XOR2_X1   g216(.A(G2427), .B(G2430), .Z(new_n642));
  OAI21_X1  g217(.A(KEYINPUT14), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT81), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n651), .B(new_n652), .Z(new_n653));
  AND2_X1   g228(.A1(new_n653), .A2(G14), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2067), .B(G2678), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT17), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n658), .B2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT82), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT83), .ZN(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n670), .A2(new_n671), .ZN(new_n677));
  AOI22_X1  g252(.A1(new_n675), .A2(new_n676), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  OR3_X1    g253(.A1(new_n672), .A2(new_n677), .A3(new_n674), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n678), .B(new_n679), .C1(new_n676), .C2(new_n675), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  INV_X1    g258(.A(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n682), .B(new_n686), .ZN(G229));
  NOR2_X1   g262(.A1(G16), .A2(G23), .ZN(new_n688));
  INV_X1    g263(.A(G288), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(G16), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT33), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G22), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G166), .B2(new_n693), .ZN(new_n695));
  INV_X1    g270(.A(G1971), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(G6), .B(G305), .S(G16), .Z(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n692), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT34), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n478), .A2(G119), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n465), .A2(G131), .ZN(new_n707));
  OAI21_X1  g282(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n475), .A2(G107), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n706), .B(new_n707), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G29), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G25), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT35), .B(G1991), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(G290), .A2(KEYINPUT84), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n597), .A2(new_n598), .B1(G651), .B2(new_n602), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT84), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n693), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G16), .A2(G24), .ZN(new_n722));
  OR3_X1    g297(.A1(new_n721), .A2(G1986), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(G1986), .B1(new_n721), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n714), .A2(new_n715), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n705), .A2(new_n716), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(KEYINPUT85), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n730), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n705), .A2(new_n727), .A3(new_n732), .A4(new_n716), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g309(.A1(KEYINPUT24), .A2(G34), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT24), .A2(G34), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n735), .A2(new_n712), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G160), .B2(new_n712), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G27), .A2(G29), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G164), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2078), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT29), .B(G2090), .ZN(new_n746));
  NAND2_X1  g321(.A1(G162), .A2(G29), .ZN(new_n747));
  OR2_X1    g322(.A1(G29), .A2(G35), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AND3_X1   g324(.A1(new_n747), .A2(new_n748), .A3(new_n746), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n745), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G5), .A2(G16), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G171), .B2(G16), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(G1961), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n693), .A2(G21), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G168), .B2(new_n693), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n712), .B1(new_n759), .B2(G28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(G28), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT94), .Z(new_n762));
  OAI21_X1  g337(.A(new_n758), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n712), .A2(G32), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n478), .A2(G129), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT91), .Z(new_n766));
  AND2_X1   g341(.A1(new_n466), .A2(G105), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT26), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n767), .B(new_n769), .C1(G141), .C2(new_n465), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(G29), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT27), .B(G1996), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n772), .A2(new_n773), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G2084), .B2(new_n738), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n753), .A2(G1961), .ZN(new_n780));
  OR3_X1    g355(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n754), .B(new_n763), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n734), .A2(new_n742), .A3(new_n751), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n693), .A2(G19), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n549), .B2(new_n693), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1341), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n614), .A2(G16), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G4), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT87), .B(G1348), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT86), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n693), .A2(KEYINPUT23), .A3(G20), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT23), .ZN(new_n795));
  INV_X1    g370(.A(G20), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(G16), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n794), .B(new_n797), .C1(new_n620), .C2(new_n693), .ZN(new_n798));
  INV_X1    g373(.A(G1956), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n789), .A2(new_n792), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n793), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n637), .A2(new_n712), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT93), .Z(new_n805));
  XOR2_X1   g380(.A(KEYINPUT31), .B(G11), .Z(new_n806));
  NOR4_X1   g381(.A1(new_n802), .A2(new_n803), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n712), .A2(G33), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n466), .A2(G103), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT89), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT25), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n465), .A2(G139), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n483), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n475), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT90), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n809), .B1(new_n818), .B2(new_n712), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(G2072), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n478), .A2(G128), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n465), .A2(G140), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n475), .A2(G116), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n821), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G29), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n712), .A2(G26), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(G2067), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n820), .A2(new_n832), .ZN(new_n833));
  NOR4_X1   g408(.A1(new_n784), .A2(new_n787), .A3(new_n808), .A4(new_n833), .ZN(G311));
  INV_X1    g409(.A(new_n784), .ZN(new_n835));
  INV_X1    g410(.A(new_n787), .ZN(new_n836));
  INV_X1    g411(.A(new_n833), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n835), .A2(new_n836), .A3(new_n807), .A4(new_n837), .ZN(G150));
  NAND2_X1  g413(.A1(G80), .A2(G543), .ZN(new_n839));
  INV_X1    g414(.A(G67), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n542), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n516), .A2(G55), .B1(G651), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n519), .A2(G93), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n614), .A2(G559), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT39), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n844), .A2(new_n549), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n548), .A2(new_n842), .A3(new_n843), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n850), .B(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n846), .B1(new_n854), .B2(G860), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT97), .ZN(G145));
  NAND2_X1  g431(.A1(new_n478), .A2(G130), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n465), .A2(G142), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n475), .A2(G118), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n857), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n710), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n818), .B(new_n825), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n482), .A2(new_n485), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n482), .B2(new_n485), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n490), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n630), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n864), .A2(new_n870), .ZN(new_n872));
  XNOR2_X1  g447(.A(G160), .B(new_n637), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(G162), .Z(new_n874));
  INV_X1    g449(.A(new_n771), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n871), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n871), .B2(new_n872), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n863), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n871), .A2(new_n872), .ZN(new_n880));
  INV_X1    g455(.A(new_n876), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n871), .A2(new_n872), .A3(new_n876), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n862), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n879), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n625), .B(new_n853), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n607), .A2(new_n611), .A3(new_n613), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n620), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g466(.A1(G299), .A2(new_n611), .A3(new_n607), .A4(new_n613), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n892), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT41), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(KEYINPUT99), .A3(new_n898), .ZN(new_n899));
  OR3_X1    g474(.A1(new_n895), .A2(KEYINPUT99), .A3(new_n896), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(new_n900), .A3(new_n889), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n888), .B1(new_n894), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(G290), .A2(new_n689), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n718), .A2(G288), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n523), .B(G305), .ZN(new_n907));
  OR3_X1    g482(.A1(new_n906), .A2(KEYINPUT100), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n905), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n718), .A2(G288), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT100), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n904), .A2(new_n905), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n913), .A3(new_n907), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n894), .A2(new_n901), .A3(new_n888), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n903), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n903), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n844), .A2(new_n617), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(G295));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n920), .ZN(G331));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  NAND2_X1  g499(.A1(G168), .A2(KEYINPUT101), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n926));
  NAND2_X1  g501(.A1(G286), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(G301), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n534), .A2(new_n535), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT75), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n932), .A2(KEYINPUT101), .A3(G168), .A4(new_n533), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n853), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n853), .A2(new_n928), .A3(new_n933), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(KEYINPUT103), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n895), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT104), .ZN(new_n943));
  OR3_X1    g518(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT102), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n936), .A2(KEYINPUT102), .A3(new_n937), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n899), .A2(new_n900), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(new_n947), .A3(new_n895), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n943), .A2(new_n915), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n885), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n947), .B1(new_n941), .B2(new_n895), .ZN(new_n951));
  AOI211_X1 g526(.A(KEYINPUT104), .B(new_n893), .C1(new_n938), .C2(new_n940), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n915), .B1(new_n953), .B2(new_n946), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n924), .B1(new_n950), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n915), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n897), .B(KEYINPUT105), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n941), .B1(new_n957), .B2(new_n898), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n893), .B1(new_n944), .B2(new_n945), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(new_n949), .A3(KEYINPUT43), .A4(new_n885), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n923), .B1(new_n955), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT43), .B1(new_n950), .B2(new_n954), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(new_n949), .A3(new_n924), .A4(new_n885), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n923), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n963), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT44), .B1(new_n964), .B2(new_n965), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT106), .B1(new_n962), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(G397));
  INV_X1    g547(.A(KEYINPUT61), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT57), .ZN(new_n974));
  INV_X1    g549(.A(new_n566), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT117), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n560), .B2(new_n563), .ZN(new_n977));
  OAI21_X1  g552(.A(G91), .B1(new_n581), .B2(new_n582), .ZN(new_n978));
  INV_X1    g553(.A(new_n563), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(KEYINPUT117), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n975), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n974), .B1(new_n981), .B2(KEYINPUT116), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n974), .B1(new_n564), .B2(new_n566), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n490), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n486), .A2(KEYINPUT98), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n482), .A2(new_n485), .A3(new_n865), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT50), .B1(new_n989), .B2(G1384), .ZN(new_n990));
  AND2_X1   g565(.A1(G160), .A2(G40), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n493), .A2(new_n992), .A3(new_n993), .A4(new_n494), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n990), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n799), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n493), .A2(new_n993), .A3(new_n494), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n868), .A2(KEYINPUT45), .A3(new_n993), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT56), .B(G2072), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n999), .A2(new_n991), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  AND4_X1   g577(.A1(new_n982), .A2(new_n985), .A3(new_n996), .A4(new_n1002), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n982), .A2(new_n985), .B1(new_n996), .B2(new_n1002), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n973), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n868), .A2(new_n993), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G160), .A2(G40), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1006), .A2(new_n1007), .A3(G2067), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n868), .A2(new_n992), .A3(new_n993), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n486), .A2(KEYINPUT71), .A3(new_n490), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT71), .B1(new_n486), .B2(new_n490), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1010), .A2(new_n1011), .A3(G1384), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1009), .B(new_n991), .C1(new_n1012), .C2(new_n992), .ZN(new_n1013));
  INV_X1    g588(.A(new_n790), .ZN(new_n1014));
  AOI211_X1 g589(.A(new_n614), .B(new_n1008), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1008), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n890), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT60), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n982), .A2(new_n985), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n996), .A2(new_n1002), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n982), .A2(new_n985), .A3(new_n996), .A4(new_n1002), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(KEYINPUT61), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1005), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1996), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n999), .A2(new_n1026), .A3(new_n991), .A4(new_n1000), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n987), .A2(new_n988), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n1030), .B2(new_n490), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1007), .B1(new_n1031), .B2(KEYINPUT45), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1032), .A2(KEYINPUT118), .A3(new_n1026), .A4(new_n999), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT58), .B(G1341), .Z(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1029), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n549), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n1036), .B2(new_n549), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1041), .A2(KEYINPUT60), .A3(new_n890), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1025), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1023), .B1(new_n1004), .B2(new_n1018), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT119), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n998), .B1(new_n989), .B2(G1384), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n493), .A2(KEYINPUT45), .A3(new_n993), .A4(new_n494), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n991), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n757), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1007), .B1(new_n997), .B2(KEYINPUT50), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(new_n740), .A3(new_n1009), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  NOR2_X1   g629(.A1(G168), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n1057));
  OAI211_X1 g632(.A(G8), .B(new_n1057), .C1(new_n1053), .C2(G286), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1054), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1061));
  OAI211_X1 g636(.A(KEYINPUT121), .B(new_n1057), .C1(new_n1061), .C2(new_n1055), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1053), .A2(new_n1064), .A3(G8), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI22_X1  g642(.A1(new_n1061), .A2(new_n1064), .B1(new_n1054), .B2(G168), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1056), .B1(new_n1063), .B2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1071));
  NAND2_X1  g646(.A1(G171), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(KEYINPUT54), .B2(G171), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n1074));
  INV_X1    g649(.A(G2078), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1047), .A2(KEYINPUT53), .A3(new_n1075), .A4(new_n991), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1048), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1961), .B1(new_n1051), .B2(new_n1009), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1074), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1961), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1013), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(KEYINPUT124), .C1(new_n1077), .C2(new_n1076), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1032), .A2(new_n1075), .A3(new_n999), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1073), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1089));
  NOR2_X1   g664(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n572), .B1(new_n571), .B2(new_n520), .ZN(new_n1093));
  AND4_X1   g668(.A1(new_n572), .A2(new_n507), .A3(new_n520), .A4(new_n522), .ZN(new_n1094));
  OAI211_X1 g669(.A(G8), .B(new_n1092), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1054), .B1(new_n573), .B2(new_n574), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(new_n1089), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n990), .A2(new_n991), .A3(new_n994), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT110), .B(G2090), .Z(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1000), .B(new_n991), .C1(new_n1012), .C2(KEYINPUT45), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT109), .B(G1971), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1098), .A2(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1054), .B1(new_n1103), .B2(KEYINPUT114), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1099), .B2(new_n995), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1097), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1051), .A2(new_n1009), .A3(new_n1100), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1054), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1097), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n519), .A2(G86), .B1(G651), .B2(new_n588), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n592), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G1981), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT112), .B(G1981), .Z(new_n1116));
  NAND4_X1  g691(.A1(new_n583), .A2(new_n591), .A3(new_n592), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT113), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1115), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT49), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1124), .A2(new_n1054), .ZN(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT49), .B(new_n1115), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(G1976), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1125), .B1(new_n1128), .B2(G288), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT52), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT52), .B1(G288), .B2(new_n1128), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1125), .B(new_n1131), .C1(new_n1128), .C2(G288), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1112), .A2(new_n1127), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1088), .A2(new_n1109), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1087), .B1(KEYINPUT54), .B2(G301), .ZN(new_n1135));
  AND2_X1   g710(.A1(G301), .A2(new_n1071), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1076), .B1(KEYINPUT45), .B2(new_n1031), .ZN(new_n1137));
  OR4_X1    g712(.A1(new_n1079), .A2(new_n1135), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1070), .A2(new_n1134), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1036), .A2(new_n549), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1036), .A2(new_n1037), .A3(new_n549), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1144), .A2(new_n1005), .A3(new_n1024), .A4(new_n1019), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1140), .B(new_n1044), .C1(new_n1145), .C2(new_n1042), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1046), .A2(new_n1139), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1133), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1061), .A2(G168), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1097), .ZN(new_n1150));
  OAI21_X1  g725(.A(G8), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1103), .A2(KEYINPUT114), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1148), .A2(new_n1149), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT115), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT115), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1148), .A2(new_n1153), .A3(new_n1157), .A4(new_n1149), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1111), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1156), .B1(new_n1160), .B2(new_n1150), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1148), .A2(new_n1161), .A3(new_n1149), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1165));
  NOR4_X1   g740(.A1(new_n1165), .A2(new_n1109), .A3(new_n1133), .A4(G301), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1167), .B(new_n1056), .C1(new_n1063), .C2(new_n1069), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1164), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1127), .A2(new_n1128), .A3(new_n689), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1112), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1127), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1171), .A2(new_n1125), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1147), .A2(new_n1163), .A3(new_n1169), .A4(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1047), .A2(new_n1007), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1176), .A2(G1996), .A3(new_n771), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1177), .A2(KEYINPUT108), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(KEYINPUT108), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n825), .B(new_n831), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1180), .B1(new_n771), .B2(G1996), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1181), .A2(new_n1176), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1178), .A2(new_n1179), .A3(new_n1182), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n710), .A2(new_n715), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n710), .A2(new_n715), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1176), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1176), .ZN(new_n1189));
  INV_X1    g764(.A(G1986), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n718), .A2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT107), .Z(new_n1192));
  NAND2_X1  g767(.A1(G290), .A2(G1986), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1189), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1188), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1175), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1180), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1176), .B1(new_n771), .B2(new_n1197), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1189), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT46), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1200), .B1(new_n1176), .B2(new_n1026), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1198), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT47), .Z(new_n1203));
  NOR2_X1   g778(.A1(new_n1192), .A2(new_n1189), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT48), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1205), .A2(new_n1188), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1185), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1183), .B1(KEYINPUT126), .B2(new_n1207), .ZN(new_n1208));
  AND2_X1   g783(.A1(new_n1207), .A2(KEYINPUT126), .ZN(new_n1209));
  OAI22_X1  g784(.A1(new_n1208), .A2(new_n1209), .B1(G2067), .B2(new_n825), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1210), .B(new_n1211), .ZN(new_n1212));
  AOI211_X1 g787(.A(new_n1203), .B(new_n1206), .C1(new_n1212), .C2(new_n1176), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1196), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g789(.A1(G401), .A2(G227), .ZN(new_n1216));
  AND2_X1   g790(.A1(new_n886), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g791(.A(G229), .ZN(new_n1218));
  AND4_X1   g792(.A1(G319), .A2(new_n1217), .A3(new_n1218), .A4(new_n966), .ZN(G308));
  NAND4_X1  g793(.A1(new_n1217), .A2(G319), .A3(new_n1218), .A4(new_n966), .ZN(G225));
endmodule


