//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n211), .B(new_n217), .C1(G97), .C2(G257), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G1), .B2(G20), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT0), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n228), .A2(G50), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n231));
  OAI22_X1  g0031(.A1(new_n230), .A2(new_n231), .B1(new_n225), .B2(new_n226), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(new_n220), .B2(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n222), .A2(new_n227), .A3(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G116), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n205), .A2(G97), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n204), .A2(G107), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G97), .B(G107), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n250), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n246), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G223), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n214), .A2(G1698), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n255), .A2(new_n258), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G87), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  OAI211_X1 g0065(.A(G1), .B(G13), .C1(new_n254), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G232), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(KEYINPUT68), .A2(G179), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT68), .A2(G179), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n268), .A2(new_n272), .A3(new_n274), .A4(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n266), .A2(new_n270), .ZN(new_n280));
  INV_X1    g0080(.A(G232), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n274), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n266), .B1(new_n262), .B2(new_n263), .ZN(new_n283));
  OAI21_X1  g0083(.A(G169), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n279), .A2(KEYINPUT73), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT73), .B1(new_n279), .B2(new_n284), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT66), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G1), .A2(G13), .ZN(new_n290));
  AND3_X1   g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G58), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(new_n215), .ZN(new_n295));
  OAI21_X1  g0095(.A(G20), .B1(new_n295), .B2(new_n201), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G159), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT7), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT3), .B(G33), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(G20), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n255), .A2(new_n260), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n300), .A2(G20), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n299), .B1(new_n306), .B2(G68), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n293), .B1(new_n307), .B2(KEYINPUT16), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT16), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT72), .B1(new_n259), .B2(G33), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT72), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(new_n254), .A3(KEYINPUT3), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n312), .A3(new_n260), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n304), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n215), .B1(new_n314), .B2(new_n302), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n309), .B1(new_n315), .B2(new_n299), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT67), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n291), .B2(new_n292), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n288), .A2(new_n290), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT66), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(KEYINPUT67), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT8), .B(G58), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G20), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(G1), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n324), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n308), .A2(new_n316), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT18), .B1(new_n287), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n279), .A2(new_n284), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT73), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n279), .A2(KEYINPUT73), .A3(new_n284), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n328), .A2(new_n331), .ZN(new_n339));
  INV_X1    g0139(.A(new_n293), .ZN(new_n340));
  INV_X1    g0140(.A(new_n299), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n303), .A2(new_n329), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n343));
  OAI211_X1 g0143(.A(KEYINPUT16), .B(new_n341), .C1(new_n343), .C2(new_n215), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n316), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT18), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n338), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n282), .A2(new_n283), .ZN(new_n349));
  INV_X1    g0149(.A(G190), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(G200), .B2(new_n349), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n339), .A2(new_n352), .A3(new_n345), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT17), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n332), .A2(KEYINPUT17), .A3(new_n352), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n333), .A2(new_n348), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  XOR2_X1   g0157(.A(new_n357), .B(KEYINPUT74), .Z(new_n358));
  INV_X1    g0158(.A(new_n324), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n318), .B2(new_n322), .ZN(new_n360));
  INV_X1    g0160(.A(new_n330), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(G50), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n323), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n364));
  INV_X1    g0164(.A(G150), .ZN(new_n365));
  INV_X1    g0165(.A(new_n297), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n329), .A2(G33), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n364), .B1(new_n365), .B2(new_n366), .C1(new_n326), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n359), .A2(new_n213), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n362), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT9), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n257), .A2(G222), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n301), .B(new_n374), .C1(new_n256), .C2(new_n257), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(new_n267), .C1(G77), .C2(new_n301), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n376), .B(new_n274), .C1(new_n214), .C2(new_n280), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G200), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n362), .A2(new_n369), .A3(KEYINPUT9), .A4(new_n370), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n377), .A2(new_n350), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n373), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT10), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n266), .A2(G238), .A3(new_n270), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G97), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(G226), .A2(G1698), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n281), .B2(G1698), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n385), .B1(new_n387), .B2(new_n301), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n274), .B(new_n383), .C1(new_n388), .C2(new_n266), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT13), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT71), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n281), .A2(G1698), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(G226), .B2(G1698), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n384), .B1(new_n393), .B2(new_n303), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n267), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n395), .A2(new_n396), .A3(new_n274), .A4(new_n383), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n390), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n389), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(G169), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT14), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n398), .A2(KEYINPUT14), .A3(G169), .A4(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n390), .A2(G179), .A3(new_n397), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n215), .A2(G20), .ZN(new_n407));
  INV_X1    g0207(.A(G77), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n407), .B1(new_n367), .B2(new_n408), .C1(new_n366), .C2(new_n213), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n363), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT11), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G13), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n407), .A2(G1), .A3(new_n413), .ZN(new_n414));
  XOR2_X1   g0214(.A(new_n414), .B(KEYINPUT12), .Z(new_n415));
  NAND3_X1  g0215(.A1(new_n363), .A2(KEYINPUT11), .A3(new_n409), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n293), .A2(G68), .A3(new_n361), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n412), .A2(new_n415), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n406), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(G169), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n377), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n371), .B(new_n421), .C1(new_n377), .C2(new_n278), .ZN(new_n422));
  INV_X1    g0222(.A(new_n418), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n390), .A2(G190), .A3(new_n397), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n398), .A2(G200), .A3(new_n399), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AND4_X1   g0226(.A1(new_n382), .A2(new_n419), .A3(new_n422), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n326), .A2(KEYINPUT69), .ZN(new_n428));
  OR2_X1    g0228(.A1(KEYINPUT8), .A2(G58), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT69), .ZN(new_n430));
  NAND2_X1  g0230(.A1(KEYINPUT8), .A2(G58), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n297), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G20), .A2(G77), .ZN(new_n434));
  XOR2_X1   g0234(.A(KEYINPUT15), .B(G87), .Z(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(new_n329), .A3(G33), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n340), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n359), .A2(new_n408), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n293), .A2(G77), .A3(new_n361), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G238), .A2(G1698), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n301), .B(new_n442), .C1(new_n281), .C2(G1698), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(new_n267), .C1(G107), .C2(new_n301), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n271), .A2(G244), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n274), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n420), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT70), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n446), .A2(new_n278), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT70), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n441), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n441), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n446), .A2(G200), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n454), .B(new_n455), .C1(new_n350), .C2(new_n446), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n358), .A2(new_n427), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n384), .A2(new_n329), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT76), .B(G87), .ZN(new_n461));
  OAI211_X1 g0261(.A(KEYINPUT19), .B(new_n460), .C1(new_n461), .C2(new_n206), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n301), .A2(new_n329), .A3(G68), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n384), .A2(G20), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n462), .B(new_n463), .C1(KEYINPUT19), .C2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n435), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n465), .A2(new_n340), .B1(new_n359), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n254), .A2(G1), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n360), .A2(G87), .A3(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n216), .A2(new_n257), .ZN(new_n472));
  INV_X1    g0272(.A(G244), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G1698), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n255), .A2(new_n472), .A3(new_n260), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G116), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n266), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n269), .A2(G45), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(new_n273), .ZN(new_n479));
  AND2_X1   g0279(.A1(G33), .A2(G41), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n478), .B(G250), .C1(new_n480), .C2(new_n290), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n477), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n350), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(G200), .B2(new_n483), .ZN(new_n485));
  NOR4_X1   g0285(.A1(new_n477), .A2(new_n278), .A3(new_n482), .A4(new_n479), .ZN(new_n486));
  INV_X1    g0286(.A(new_n479), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n475), .A2(new_n476), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n481), .C1(new_n488), .C2(new_n266), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n486), .B1(new_n420), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n360), .A2(new_n435), .A3(new_n469), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n467), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n471), .A2(new_n485), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n205), .B1(new_n314), .B2(new_n302), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n297), .A2(G77), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT6), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n496), .A2(new_n204), .A3(G107), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n497), .B1(new_n496), .B2(new_n251), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n495), .B1(new_n498), .B2(new_n329), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n340), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n360), .A2(G97), .A3(new_n469), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n359), .A2(new_n204), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n265), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G41), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n479), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G45), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(G1), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(new_n504), .A3(new_n506), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n266), .ZN(new_n511));
  INV_X1    g0311(.A(G257), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n255), .A2(new_n260), .A3(G250), .ZN(new_n514));
  NOR2_X1   g0314(.A1(KEYINPUT75), .A2(KEYINPUT4), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G1698), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n255), .A2(new_n260), .A3(G244), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n515), .B1(G33), .B2(G283), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n255), .A2(new_n260), .A3(G244), .A4(new_n257), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT75), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n518), .B(new_n520), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  AOI211_X1 g0325(.A(G190), .B(new_n513), .C1(new_n525), .C2(new_n267), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n518), .A2(new_n520), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n524), .B1(new_n521), .B2(new_n522), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n267), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n513), .ZN(new_n530));
  AOI21_X1  g0330(.A(G200), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n503), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n529), .A2(new_n277), .A3(new_n530), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n513), .B1(new_n525), .B2(new_n267), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n533), .B(new_n534), .C1(G169), .C2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n493), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT24), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT23), .B1(new_n329), .B2(G107), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(new_n205), .A3(G20), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n329), .A2(G33), .A3(G116), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT84), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT84), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n539), .A2(new_n541), .A3(new_n542), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n255), .A2(new_n260), .A3(new_n329), .A4(G87), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT22), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT22), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n301), .A2(new_n550), .A3(new_n329), .A4(G87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT83), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n547), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n547), .B2(new_n552), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n538), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n547), .A2(new_n552), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT83), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n547), .A2(new_n552), .A3(new_n553), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(KEYINPUT24), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n556), .A2(new_n560), .A3(new_n340), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n269), .A2(new_n205), .A3(G13), .A4(G20), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n562), .B(KEYINPUT25), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n325), .A2(new_n468), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n563), .B1(new_n564), .B2(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n301), .A2(G257), .A3(G1698), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G294), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n566), .B(new_n567), .C1(G1698), .C2(new_n514), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n267), .ZN(new_n569));
  INV_X1    g0369(.A(new_n511), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G264), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n507), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G200), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n568), .A2(new_n267), .B1(G264), .B2(new_n570), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(new_n350), .A3(new_n507), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n561), .A2(new_n565), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n537), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(G264), .A2(G1698), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n255), .A2(new_n260), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT77), .ZN(new_n582));
  XNOR2_X1  g0382(.A(KEYINPUT78), .B(G303), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n303), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n255), .A2(new_n260), .A3(G257), .A4(new_n257), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT77), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n255), .A2(new_n260), .A3(new_n580), .A4(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n582), .A2(new_n584), .A3(new_n585), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n267), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n507), .B1(new_n511), .B2(new_n210), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n420), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n468), .A2(new_n209), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n320), .A2(new_n593), .A3(new_n324), .A4(new_n321), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n359), .A2(new_n209), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n288), .A2(new_n290), .B1(G20), .B2(new_n209), .ZN(new_n596));
  NAND2_X1  g0396(.A1(G33), .A2(G283), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n597), .B(new_n329), .C1(G33), .C2(new_n204), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n596), .A2(KEYINPUT20), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT20), .B1(new_n596), .B2(new_n598), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n594), .B(new_n595), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(KEYINPUT79), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT79), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n359), .A2(new_n209), .A3(new_n468), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n293), .A2(new_n604), .B1(new_n209), .B2(new_n359), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n596), .A2(new_n598), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT20), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n596), .A2(KEYINPUT20), .A3(new_n598), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n603), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n592), .B1(new_n602), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT81), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT21), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT81), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT80), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n590), .B1(new_n588), .B2(new_n267), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n592), .A2(KEYINPUT21), .B1(G179), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n602), .A2(new_n611), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n589), .A2(new_n591), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(KEYINPUT21), .A3(G169), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n619), .A2(G179), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n602), .A2(new_n611), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(KEYINPUT80), .A3(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n615), .A2(new_n617), .B1(new_n622), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n561), .A2(new_n565), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n572), .A2(new_n420), .ZN(new_n631));
  INV_X1    g0431(.A(G179), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n575), .A2(new_n632), .A3(new_n507), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT82), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n619), .A2(new_n573), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n627), .B2(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n621), .B(KEYINPUT82), .C1(new_n573), .C2(new_n619), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n637), .B(new_n638), .C1(new_n350), .C2(new_n623), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n579), .A2(new_n629), .A3(new_n634), .A4(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n459), .A2(new_n640), .ZN(G372));
  INV_X1    g0441(.A(new_n422), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n355), .A2(new_n356), .ZN(new_n643));
  INV_X1    g0443(.A(new_n419), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n426), .A2(new_n450), .A3(new_n449), .A4(new_n452), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n346), .A2(new_n334), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(new_n347), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n642), .B1(new_n649), .B2(new_n382), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n561), .A2(new_n565), .A3(new_n577), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT85), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n483), .B2(G169), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n489), .A2(KEYINPUT85), .A3(new_n420), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n486), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n655), .A2(new_n492), .B1(new_n471), .B2(new_n485), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n651), .A2(new_n656), .A3(new_n536), .A4(new_n532), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n617), .A2(new_n615), .B1(new_n627), .B2(new_n626), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n634), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n493), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT26), .B1(new_n663), .B2(new_n536), .ZN(new_n664));
  INV_X1    g0464(.A(new_n536), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n656), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n655), .A2(new_n492), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n664), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n650), .B1(new_n459), .B2(new_n672), .ZN(G369));
  NOR2_X1   g0473(.A1(new_n413), .A2(G20), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n269), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n621), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n629), .A2(new_n639), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n659), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n661), .A2(new_n681), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n630), .A2(new_n680), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n651), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n634), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n634), .A2(new_n680), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n629), .A2(new_n680), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n690), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(G399));
  NOR2_X1   g0497(.A1(new_n461), .A2(new_n206), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n209), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n224), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n700), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n230), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n629), .A2(new_n634), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n658), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n665), .A2(new_n656), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT26), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n711), .A2(new_n668), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n665), .A2(new_n666), .A3(new_n493), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n707), .B1(new_n714), .B2(new_n681), .ZN(new_n715));
  AOI211_X1 g0515(.A(KEYINPUT29), .B(new_n680), .C1(new_n662), .C2(new_n670), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n623), .A2(new_n632), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n575), .A3(new_n483), .A4(new_n535), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n625), .A2(new_n489), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(KEYINPUT30), .A3(new_n575), .A4(new_n535), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n529), .A2(new_n530), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n483), .A2(new_n278), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n623), .A3(new_n572), .A4(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT86), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n619), .B1(new_n507), .B2(new_n575), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(KEYINPUT86), .A3(new_n725), .A4(new_n726), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n680), .B1(new_n724), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n727), .ZN(new_n736));
  OAI211_X1 g0536(.A(KEYINPUT31), .B(new_n680), .C1(new_n724), .C2(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n735), .B(new_n737), .C1(new_n640), .C2(new_n680), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n717), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n706), .B1(new_n741), .B2(G1), .ZN(G364));
  INV_X1    g0542(.A(new_n686), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n674), .A2(G45), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n703), .A2(G1), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G330), .B2(new_n685), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n632), .A2(G200), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT90), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G190), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n350), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G107), .A2(new_n752), .B1(new_n753), .B2(new_n461), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n277), .A2(new_n329), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n350), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n756), .A2(G190), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n754), .B1(new_n213), .B2(new_n758), .C1(new_n215), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n350), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n632), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n301), .B1(new_n765), .B2(new_n204), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT89), .B(G159), .Z(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n329), .A2(G190), .A3(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n632), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT32), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n278), .A2(new_n769), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n755), .A2(new_n762), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n774), .A2(KEYINPUT88), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(KEYINPUT88), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n772), .B1(new_n408), .B2(new_n773), .C1(new_n777), .C2(new_n294), .ZN(new_n778));
  OR3_X1    g0578(.A1(new_n761), .A2(new_n766), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n777), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n780), .A2(G322), .B1(new_n759), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT92), .ZN(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  INV_X1    g0584(.A(new_n753), .ZN(new_n785));
  INV_X1    g0585(.A(G303), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n303), .B1(new_n784), .B2(new_n773), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G283), .B2(new_n752), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n757), .A2(G326), .ZN(new_n789));
  INV_X1    g0589(.A(G294), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n790), .B2(new_n765), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(KEYINPUT91), .ZN(new_n792));
  INV_X1    g0592(.A(new_n770), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G329), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n791), .A2(KEYINPUT91), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n788), .A2(new_n792), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n779), .B1(new_n783), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n290), .B1(G20), .B2(new_n420), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n798), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n246), .A2(G45), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n701), .A2(new_n301), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n803), .B(new_n804), .C1(G45), .C2(new_n230), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n301), .A2(new_n224), .ZN(new_n806));
  XNOR2_X1  g0606(.A(G355), .B(KEYINPUT87), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(G116), .B2(new_n224), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n797), .A2(new_n798), .B1(new_n802), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n801), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n685), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n748), .B1(new_n745), .B2(new_n811), .ZN(G396));
  NAND2_X1  g0612(.A1(new_n671), .A2(new_n681), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n454), .A2(new_n681), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n453), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n457), .B2(new_n814), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n453), .A2(new_n814), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n453), .A2(new_n456), .ZN(new_n819));
  INV_X1    g0619(.A(new_n814), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n657), .B1(new_n634), .B2(new_n659), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n821), .B(new_n681), .C1(new_n822), .C2(new_n669), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n817), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n739), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n817), .A2(G330), .A3(new_n738), .A4(new_n823), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n745), .A3(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G137), .A2(new_n757), .B1(new_n759), .B2(G150), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT93), .B(G143), .Z(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n768), .B2(new_n773), .C1(new_n777), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT34), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n793), .A2(G132), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(new_n832), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n301), .B1(new_n294), .B2(new_n765), .C1(new_n785), .C2(new_n213), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G68), .B2(new_n752), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n785), .A2(new_n205), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n765), .A2(new_n204), .B1(new_n773), .B2(new_n209), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n780), .B2(G294), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G87), .A2(new_n752), .B1(new_n759), .B2(G283), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n303), .B1(new_n770), .B2(new_n784), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n757), .B2(G303), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n838), .B1(new_n839), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n798), .A2(new_n799), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n846), .A2(new_n798), .B1(new_n408), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n848), .B(new_n746), .C1(new_n800), .C2(new_n821), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n827), .A2(new_n849), .ZN(G384));
  INV_X1    g0650(.A(KEYINPUT40), .ZN(new_n851));
  INV_X1    g0651(.A(new_n678), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n346), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n853), .A2(new_n854), .A3(new_n353), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n338), .A2(new_n346), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n307), .A2(KEYINPUT16), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(new_n363), .A3(new_n344), .ZN(new_n859));
  INV_X1    g0659(.A(new_n334), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n859), .A2(new_n339), .B1(new_n860), .B2(new_n678), .ZN(new_n861));
  INV_X1    g0661(.A(new_n353), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT37), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n857), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT97), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n678), .B1(new_n859), .B2(new_n339), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n357), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n865), .B1(new_n357), .B2(new_n866), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(KEYINPUT38), .B(new_n864), .C1(new_n867), .C2(new_n868), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(KEYINPUT31), .B(new_n680), .C1(new_n724), .C2(new_n732), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n735), .B(new_n874), .C1(new_n640), .C2(new_n680), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n418), .A2(new_n680), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n406), .A2(KEYINPUT96), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT96), .ZN(new_n879));
  INV_X1    g0679(.A(new_n405), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n402), .B2(new_n403), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n879), .B1(new_n881), .B2(new_n876), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n426), .B(new_n876), .C1(new_n881), .C2(new_n423), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n816), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n875), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n851), .B1(new_n873), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n853), .B1(new_n648), .B2(new_n643), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n647), .A2(new_n853), .A3(new_n353), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n855), .A2(new_n856), .B1(new_n889), .B2(KEYINPUT37), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n870), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n872), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n892), .A2(KEYINPUT40), .A3(new_n875), .A4(new_n885), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n458), .A2(new_n875), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n894), .B(new_n895), .Z(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(G330), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n648), .A2(new_n852), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n871), .A2(new_n872), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n453), .A2(new_n680), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT95), .Z(new_n901));
  NAND2_X1  g0701(.A1(new_n823), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n883), .A2(new_n884), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n899), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n871), .A2(KEYINPUT39), .A3(new_n872), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n892), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n644), .A2(new_n681), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n898), .B(new_n904), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n458), .B1(new_n715), .B2(new_n716), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n650), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n910), .B(new_n912), .Z(new_n913));
  XNOR2_X1  g0713(.A(new_n897), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n269), .B2(new_n674), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n230), .A2(new_n408), .A3(new_n295), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n215), .A2(G50), .ZN(new_n917));
  OAI211_X1 g0717(.A(G1), .B(new_n413), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT35), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n231), .B1(new_n498), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(G116), .C1(new_n919), .C2(new_n498), .ZN(new_n921));
  XOR2_X1   g0721(.A(KEYINPUT94), .B(KEYINPUT36), .Z(new_n922));
  XNOR2_X1  g0722(.A(new_n921), .B(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n915), .A2(new_n918), .A3(new_n923), .ZN(G367));
  INV_X1    g0724(.A(G283), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n303), .B1(new_n773), .B2(new_n925), .C1(new_n205), .C2(new_n765), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(G294), .B2(new_n759), .ZN(new_n927));
  AOI22_X1  g0727(.A1(G97), .A2(new_n752), .B1(new_n757), .B2(G311), .ZN(new_n928));
  INV_X1    g0728(.A(new_n583), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n927), .B(new_n928), .C1(new_n929), .C2(new_n777), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT103), .B1(new_n753), .B2(G116), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT46), .Z(new_n932));
  AOI211_X1 g0732(.A(new_n930), .B(new_n932), .C1(G317), .C2(new_n793), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n753), .A2(G58), .B1(G137), .B2(new_n793), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT104), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n765), .A2(new_n215), .ZN(new_n936));
  AOI22_X1  g0736(.A1(G77), .A2(new_n752), .B1(new_n757), .B2(new_n829), .ZN(new_n937));
  INV_X1    g0737(.A(new_n773), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n759), .A2(new_n767), .B1(G50), .B2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n937), .B(new_n939), .C1(new_n365), .C2(new_n777), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n935), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n933), .B1(new_n301), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT47), .Z(new_n943));
  AOI21_X1  g0743(.A(new_n745), .B1(new_n943), .B2(new_n798), .ZN(new_n944));
  INV_X1    g0744(.A(new_n804), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n802), .B1(new_n224), .B2(new_n466), .C1(new_n242), .C2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n656), .B1(new_n471), .B2(new_n681), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT98), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n668), .A2(new_n471), .A3(new_n681), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(KEYINPUT98), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n944), .B(new_n946), .C1(new_n810), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n744), .A2(G1), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n691), .B1(new_n629), .B2(new_n680), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n695), .A2(new_n687), .A3(new_n690), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n743), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n686), .A2(new_n955), .A3(new_n954), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n740), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n725), .A2(new_n420), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n961), .A2(new_n534), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n503), .A2(new_n681), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT99), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n532), .A2(new_n536), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n964), .B(new_n965), .C1(new_n966), .C2(new_n963), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n962), .A2(KEYINPUT99), .A3(new_n963), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n696), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT45), .ZN(new_n972));
  XOR2_X1   g0772(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OR3_X1    g0774(.A1(new_n696), .A2(new_n970), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n696), .B2(new_n970), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g0777(.A(KEYINPUT102), .B(new_n692), .C1(new_n972), .C2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n692), .A2(KEYINPUT102), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT45), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n971), .B(new_n980), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n981), .A2(new_n693), .A3(new_n975), .A4(new_n976), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n960), .A2(new_n978), .A3(new_n979), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n741), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n702), .B(KEYINPUT41), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n953), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n955), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT100), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n987), .A2(new_n988), .A3(new_n970), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT100), .B1(new_n955), .B2(new_n969), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT42), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n536), .B1(new_n969), .B2(new_n634), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n681), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT42), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n693), .A2(new_n969), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n999), .B1(new_n997), .B2(new_n1000), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n1001), .A2(new_n1002), .B1(KEYINPUT43), .B2(new_n951), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n997), .A2(new_n1000), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n998), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n952), .B1(new_n986), .B2(new_n1009), .ZN(G387));
  INV_X1    g0810(.A(new_n953), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n959), .A2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G311), .A2(new_n759), .B1(new_n757), .B2(G322), .ZN(new_n1013));
  INV_X1    g0813(.A(G317), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(new_n929), .B2(new_n773), .C1(new_n1014), .C2(new_n777), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT48), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n925), .B2(new_n765), .C1(new_n790), .C2(new_n785), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT49), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n301), .B1(new_n752), .B2(G116), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1019), .B(new_n1022), .C1(G326), .C2(new_n793), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n764), .A2(new_n435), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n301), .C1(new_n365), .C2(new_n770), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n752), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1026), .A2(new_n204), .B1(new_n215), .B2(new_n773), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(G50), .C2(new_n780), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G159), .A2(new_n757), .B1(new_n759), .B2(new_n327), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(new_n408), .C2(new_n785), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT106), .Z(new_n1031));
  OAI21_X1  g0831(.A(new_n798), .B1(new_n1023), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n428), .A2(new_n432), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1033), .A2(G50), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n1035));
  AOI21_X1  g0835(.A(new_n699), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1036), .B(new_n508), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G68), .B2(G77), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n804), .B1(new_n239), .B2(new_n508), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1038), .A2(new_n1039), .B1(G107), .B2(new_n224), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n700), .A2(new_n806), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n802), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n691), .A2(new_n801), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1032), .A2(new_n746), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n960), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n959), .A2(new_n740), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT107), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n702), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1012), .B(new_n1044), .C1(new_n1049), .C2(new_n1050), .ZN(G393));
  OAI21_X1  g0851(.A(new_n692), .B1(new_n972), .B2(new_n977), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1052), .A2(new_n982), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n983), .B(new_n702), .C1(new_n960), .C2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n759), .A2(new_n583), .B1(G116), .B2(new_n764), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT108), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n777), .A2(new_n784), .B1(new_n1014), .B2(new_n758), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  OAI22_X1  g0858(.A1(new_n1026), .A2(new_n205), .B1(new_n790), .B2(new_n773), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n301), .B1(new_n793), .B2(G322), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n785), .B2(new_n925), .ZN(new_n1061));
  OR4_X1    g0861(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT109), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n760), .A2(new_n213), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n780), .A2(G159), .B1(G150), .B2(new_n757), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1065), .A2(KEYINPUT51), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n764), .A2(G77), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n301), .C1(new_n770), .C2(new_n830), .ZN(new_n1068));
  INV_X1    g0868(.A(G87), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1026), .A2(new_n1069), .B1(new_n1033), .B2(new_n773), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1068), .B(new_n1070), .C1(G68), .C2(new_n753), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1065), .A2(KEYINPUT51), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1066), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1063), .B1(new_n1064), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n745), .B1(new_n1074), .B2(new_n798), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n252), .A2(new_n804), .B1(G97), .B2(new_n701), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n802), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1075), .B(new_n1077), .C1(new_n810), .C2(new_n970), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1052), .A2(new_n982), .A3(new_n953), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1054), .A2(new_n1080), .ZN(G390));
  NAND4_X1  g0881(.A1(new_n875), .A2(G330), .A3(new_n821), .A4(new_n903), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n902), .A2(new_n903), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n907), .A2(new_n905), .B1(new_n1084), .B2(new_n909), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n892), .A2(new_n909), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n714), .A2(new_n681), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n901), .B1(new_n1087), .B2(new_n816), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n903), .B(KEYINPUT110), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1083), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1084), .A2(new_n909), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n908), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1086), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n901), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n711), .A2(new_n668), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n708), .B2(new_n658), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n680), .B1(new_n1097), .B2(new_n713), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1098), .B2(new_n821), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT110), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n903), .B(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1094), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n738), .A2(G330), .A3(new_n821), .A4(new_n903), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1093), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1091), .A2(new_n1104), .A3(new_n953), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT112), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1091), .A2(new_n1104), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT111), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n738), .A2(G330), .A3(new_n821), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n903), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n902), .B1(new_n1112), .B2(new_n1083), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n875), .A2(G330), .A3(new_n821), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1099), .B(new_n1103), .C1(new_n1089), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n458), .A2(G330), .A3(new_n875), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n911), .A2(new_n650), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1108), .A2(new_n1109), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1118), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1104), .B(new_n1091), .C1(new_n1122), .C2(KEYINPUT111), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n702), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n908), .A2(new_n799), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n785), .A2(new_n1069), .B1(new_n758), .B2(new_n925), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(G107), .B2(new_n759), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n752), .A2(G68), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n303), .B1(new_n790), .B2(new_n770), .C1(new_n773), .C2(new_n204), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n780), .B2(G116), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1127), .A2(new_n1128), .A3(new_n1067), .A4(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT53), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n753), .B2(G150), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n785), .A2(KEYINPUT53), .A3(new_n365), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(G132), .C2(new_n780), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT54), .B(G143), .Z(new_n1136));
  AOI22_X1  g0936(.A1(new_n938), .A2(new_n1136), .B1(G159), .B2(new_n764), .ZN(new_n1137));
  INV_X1    g0937(.A(G128), .ZN(new_n1138));
  INV_X1    g0938(.A(G137), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1137), .B1(new_n758), .B2(new_n1138), .C1(new_n1139), .C2(new_n760), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n301), .B1(new_n1026), .B2(new_n213), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(KEYINPUT113), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1135), .B(new_n1142), .C1(KEYINPUT113), .C2(new_n1141), .ZN(new_n1143));
  INV_X1    g0943(.A(G125), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n770), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1131), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1146), .A2(new_n798), .B1(new_n326), .B2(new_n847), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1125), .A2(new_n746), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1107), .A2(new_n1124), .A3(new_n1148), .ZN(G378));
  NAND3_X1  g0949(.A1(new_n1091), .A2(new_n1104), .A3(new_n1116), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1119), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n886), .B1(new_n872), .B2(new_n871), .ZN(new_n1152));
  OAI211_X1 g0952(.A(G330), .B(new_n893), .C1(new_n1152), .C2(KEYINPUT40), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n371), .A2(new_n852), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT56), .Z(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n382), .A2(new_n422), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT55), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1157), .A2(KEYINPUT55), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1156), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1160), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n1158), .A3(new_n1155), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1153), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n887), .A2(G330), .A3(new_n1166), .A4(new_n893), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n910), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1165), .A2(new_n910), .A3(new_n1167), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1151), .B(KEYINPUT57), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT116), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1165), .A2(new_n1171), .A3(new_n1167), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n910), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1165), .A2(new_n1167), .A3(new_n1171), .A4(new_n910), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1174), .A2(new_n1175), .B1(new_n1119), .B2(new_n1150), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1170), .B(new_n702), .C1(new_n1176), .C2(KEYINPUT57), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n953), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1166), .A2(new_n799), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n753), .A2(new_n1136), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n758), .A2(new_n1144), .B1(new_n365), .B2(new_n765), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(G132), .C2(new_n759), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n1138), .B2(new_n777), .C1(new_n1139), .C2(new_n773), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1186));
  XOR2_X1   g0986(.A(KEYINPUT115), .B(G124), .Z(new_n1187));
  AOI21_X1  g0987(.A(G33), .B1(new_n793), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(G41), .B1(new_n752), .B2(new_n767), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n265), .B1(new_n259), .B2(new_n254), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(KEYINPUT114), .A3(new_n213), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n204), .A2(new_n760), .B1(new_n758), .B2(new_n209), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n936), .B(new_n1193), .C1(G58), .C2(new_n752), .ZN(new_n1194));
  AOI21_X1  g0994(.A(G41), .B1(new_n793), .B2(G283), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n466), .B2(new_n773), .C1(new_n785), .C2(new_n408), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G107), .B2(new_n780), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1194), .A2(new_n303), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT58), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT114), .B1(new_n1191), .B2(new_n213), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1190), .A2(new_n1192), .A3(new_n1200), .A4(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1203), .A2(new_n798), .B1(new_n213), .B2(new_n847), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1180), .A2(new_n746), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT117), .B1(new_n1179), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1011), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT117), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1205), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1177), .B1(new_n1206), .B2(new_n1210), .ZN(G375));
  NAND2_X1  g1011(.A1(new_n1116), .A2(new_n953), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n301), .B1(new_n773), .B2(new_n365), .C1(new_n213), .C2(new_n765), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G58), .B2(new_n752), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G159), .A2(new_n753), .B1(new_n759), .B2(new_n1136), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n1138), .B2(new_n770), .C1(new_n1139), .C2(new_n777), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n757), .A2(G132), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT118), .Z(new_n1219));
  AOI22_X1  g1019(.A1(G116), .A2(new_n759), .B1(new_n757), .B2(G294), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n1024), .C1(new_n204), .C2(new_n785), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n303), .B1(new_n770), .B2(new_n786), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n938), .B2(G107), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n1026), .B2(new_n408), .C1(new_n777), .C2(new_n925), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n1217), .A2(new_n1219), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1225), .A2(new_n798), .B1(new_n215), .B2(new_n847), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n746), .B(new_n1226), .C1(new_n1089), .C2(new_n800), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1212), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1113), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1120), .A2(new_n985), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(G381));
  OR2_X1    g1031(.A1(G375), .A2(G378), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1232), .A2(G384), .A3(G381), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1054), .A2(new_n1080), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(new_n952), .C1(new_n986), .C2(new_n1009), .ZN(new_n1235));
  OR2_X1    g1035(.A1(G393), .A2(G396), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1237), .ZN(G407));
  NAND2_X1  g1038(.A1(new_n679), .A2(G213), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT119), .ZN(new_n1240));
  OAI211_X1 g1040(.A(G407), .B(G213), .C1(new_n1232), .C2(new_n1240), .ZN(G409));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1229), .A2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1113), .A2(new_n1115), .A3(new_n1118), .A4(KEYINPUT60), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1243), .A2(new_n1120), .A3(new_n702), .A4(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1228), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT120), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G384), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n827), .A2(KEYINPUT120), .A3(new_n849), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1245), .A2(new_n1228), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G378), .B(new_n1177), .C1(new_n1206), .C2(new_n1210), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1107), .A2(new_n1124), .A3(new_n1148), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n953), .B1(new_n1169), .B2(new_n1168), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1178), .A2(new_n1151), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n985), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1256), .B1(new_n1260), .B2(new_n1209), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1255), .A2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT126), .B1(new_n1262), .B2(new_n1240), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT126), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1240), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n1255), .C2(new_n1261), .ZN(new_n1266));
  OAI211_X1 g1066(.A(KEYINPUT63), .B(new_n1254), .C1(new_n1263), .C2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1239), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n1269), .B(new_n1253), .C1(new_n1255), .C2(new_n1261), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(G2897), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1212), .A2(new_n1227), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1122), .B1(new_n1242), .B2(new_n1229), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1244), .A2(new_n702), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1272), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1248), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1252), .B(new_n1271), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT121), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1249), .A2(KEYINPUT121), .A3(new_n1252), .A4(new_n1271), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1253), .A2(G2897), .A3(new_n1265), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT122), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1262), .A2(new_n1239), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT122), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1281), .A2(new_n1286), .A3(new_n1282), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1284), .A2(new_n1285), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1270), .B1(new_n1288), .B2(KEYINPUT63), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT124), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G393), .A2(G396), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(G387), .A2(new_n1291), .B1(new_n1236), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G387), .A2(G390), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1293), .A2(KEYINPUT123), .A3(new_n1235), .A4(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1236), .A2(new_n1292), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1235), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1291), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT123), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1290), .B(new_n1295), .C1(new_n1298), .C2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT124), .B1(new_n1294), .B2(new_n1235), .ZN(new_n1304));
  OAI22_X1  g1104(.A1(new_n1304), .A2(new_n1296), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1305), .A2(KEYINPUT125), .A3(new_n1290), .A4(new_n1295), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1303), .A2(new_n1306), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1268), .A2(new_n1289), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1305), .A2(new_n1295), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1262), .A2(new_n1311), .A3(new_n1239), .A4(new_n1254), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1290), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1283), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1313), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1254), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT62), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1310), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(KEYINPUT127), .B1(new_n1308), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1262), .A2(new_n1240), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1264), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1262), .A2(KEYINPUT126), .A3(new_n1240), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1311), .B1(new_n1324), .B2(new_n1254), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1322), .A2(new_n1323), .A3(new_n1315), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1313), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1309), .B1(new_n1325), .B2(new_n1328), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1303), .A2(new_n1306), .ZN(new_n1330));
  AND2_X1   g1130(.A1(new_n1288), .A2(KEYINPUT63), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1330), .B(new_n1267), .C1(new_n1331), .C2(new_n1270), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1329), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1320), .A2(new_n1334), .ZN(G405));
  NAND2_X1  g1135(.A1(G375), .A2(new_n1256), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1336), .A2(new_n1255), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1310), .B(new_n1337), .ZN(new_n1338));
  XNOR2_X1  g1138(.A(new_n1338), .B(new_n1254), .ZN(G402));
endmodule


