

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U319 ( .A(n377), .B(KEYINPUT41), .ZN(n554) );
  NOR2_X1 U320 ( .A1(n416), .A2(n415), .ZN(n417) );
  XNOR2_X1 U321 ( .A(n383), .B(n360), .ZN(n362) );
  XNOR2_X1 U322 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U323 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U324 ( .A(n370), .B(n369), .ZN(n374) );
  OR2_X1 U325 ( .A1(n571), .A2(KEYINPUT64), .ZN(n375) );
  INV_X1 U326 ( .A(G190GAT), .ZN(n446) );
  XNOR2_X1 U327 ( .A(n446), .B(KEYINPUT58), .ZN(n447) );
  XNOR2_X1 U328 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  XOR2_X1 U329 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n288) );
  XNOR2_X1 U330 ( .A(KEYINPUT67), .B(KEYINPUT72), .ZN(n287) );
  XNOR2_X1 U331 ( .A(n288), .B(n287), .ZN(n306) );
  XOR2_X1 U332 ( .A(G197GAT), .B(G36GAT), .Z(n290) );
  XNOR2_X1 U333 ( .A(G29GAT), .B(G141GAT), .ZN(n289) );
  XNOR2_X1 U334 ( .A(n290), .B(n289), .ZN(n294) );
  XOR2_X1 U335 ( .A(KEYINPUT29), .B(G169GAT), .Z(n292) );
  XNOR2_X1 U336 ( .A(G113GAT), .B(G1GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U338 ( .A(n294), .B(n293), .Z(n304) );
  XOR2_X1 U339 ( .A(KEYINPUT7), .B(KEYINPUT70), .Z(n296) );
  XNOR2_X1 U340 ( .A(G50GAT), .B(G43GAT), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U342 ( .A(KEYINPUT8), .B(n297), .Z(n395) );
  XOR2_X1 U343 ( .A(G8GAT), .B(KEYINPUT71), .Z(n299) );
  XNOR2_X1 U344 ( .A(G22GAT), .B(G15GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n402) );
  XOR2_X1 U346 ( .A(n402), .B(KEYINPUT68), .Z(n301) );
  NAND2_X1 U347 ( .A1(G229GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n395), .B(n302), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(n306), .B(n305), .Z(n565) );
  XOR2_X1 U352 ( .A(KEYINPUT76), .B(G204GAT), .Z(n308) );
  XNOR2_X1 U353 ( .A(G106GAT), .B(G78GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n364) );
  XOR2_X1 U355 ( .A(n364), .B(G22GAT), .Z(n310) );
  NAND2_X1 U356 ( .A1(G228GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U358 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n312) );
  XNOR2_X1 U359 ( .A(G148GAT), .B(KEYINPUT22), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U361 ( .A(n314), .B(n313), .Z(n319) );
  XOR2_X1 U362 ( .A(KEYINPUT21), .B(G197GAT), .Z(n316) );
  XNOR2_X1 U363 ( .A(G218GAT), .B(KEYINPUT89), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U365 ( .A(G211GAT), .B(n317), .Z(n347) );
  XNOR2_X1 U366 ( .A(G50GAT), .B(n347), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n324) );
  XOR2_X1 U368 ( .A(KEYINPUT3), .B(KEYINPUT90), .Z(n321) );
  XNOR2_X1 U369 ( .A(G141GAT), .B(G155GAT), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n323) );
  XOR2_X1 U371 ( .A(G162GAT), .B(KEYINPUT2), .Z(n322) );
  XNOR2_X1 U372 ( .A(n323), .B(n322), .ZN(n340) );
  XNOR2_X1 U373 ( .A(n324), .B(n340), .ZN(n460) );
  XNOR2_X1 U374 ( .A(G148GAT), .B(G120GAT), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n325), .B(G57GAT), .ZN(n361) );
  XOR2_X1 U376 ( .A(G127GAT), .B(G1GAT), .Z(n399) );
  XOR2_X1 U377 ( .A(n361), .B(n399), .Z(n327) );
  NAND2_X1 U378 ( .A1(G225GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n339) );
  XOR2_X1 U380 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n329) );
  XNOR2_X1 U381 ( .A(G85GAT), .B(KEYINPUT93), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U383 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n331) );
  XNOR2_X1 U384 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U386 ( .A(n333), .B(n332), .Z(n337) );
  XNOR2_X1 U387 ( .A(G29GAT), .B(KEYINPUT82), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n334), .B(G134GAT), .ZN(n387) );
  XNOR2_X1 U389 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n335) );
  XNOR2_X1 U390 ( .A(n335), .B(KEYINPUT86), .ZN(n428) );
  XNOR2_X1 U391 ( .A(n387), .B(n428), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n341) );
  XOR2_X1 U394 ( .A(n341), .B(n340), .Z(n457) );
  XNOR2_X1 U395 ( .A(KEYINPUT94), .B(n457), .ZN(n496) );
  XOR2_X1 U396 ( .A(KEYINPUT88), .B(G169GAT), .Z(n343) );
  XNOR2_X1 U397 ( .A(KEYINPUT87), .B(KEYINPUT18), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U399 ( .A(n344), .B(KEYINPUT19), .Z(n346) );
  XNOR2_X1 U400 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n441) );
  XNOR2_X1 U402 ( .A(n441), .B(n347), .ZN(n359) );
  XOR2_X1 U403 ( .A(G190GAT), .B(G36GAT), .Z(n386) );
  XOR2_X1 U404 ( .A(KEYINPUT96), .B(KEYINPUT98), .Z(n349) );
  XNOR2_X1 U405 ( .A(G8GAT), .B(G204GAT), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U407 ( .A(n386), .B(n350), .Z(n352) );
  NAND2_X1 U408 ( .A1(G226GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U410 ( .A(n353), .B(KEYINPUT97), .Z(n357) );
  XOR2_X1 U411 ( .A(KEYINPUT77), .B(G176GAT), .Z(n355) );
  XNOR2_X1 U412 ( .A(G92GAT), .B(G64GAT), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n372) );
  XNOR2_X1 U414 ( .A(n372), .B(KEYINPUT95), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n359), .B(n358), .ZN(n499) );
  INV_X1 U417 ( .A(n499), .ZN(n512) );
  XNOR2_X1 U418 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n379) );
  XOR2_X1 U419 ( .A(G85GAT), .B(G99GAT), .Z(n383) );
  AND2_X1 U420 ( .A1(G230GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n363), .B(KEYINPUT75), .ZN(n370) );
  XOR2_X1 U422 ( .A(n364), .B(KEYINPUT78), .Z(n368) );
  XOR2_X1 U423 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n366) );
  XNOR2_X1 U424 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U426 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n371), .B(KEYINPUT73), .ZN(n398) );
  XOR2_X1 U428 ( .A(n398), .B(n372), .Z(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n571) );
  NAND2_X1 U430 ( .A1(n571), .A2(KEYINPUT64), .ZN(n376) );
  NAND2_X1 U431 ( .A1(n376), .A2(n375), .ZN(n377) );
  NOR2_X1 U432 ( .A1(n565), .A2(n554), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n416) );
  XOR2_X1 U434 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n381) );
  XNOR2_X1 U435 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U437 ( .A(n382), .B(G106GAT), .Z(n385) );
  XNOR2_X1 U438 ( .A(n383), .B(G218GAT), .ZN(n384) );
  XNOR2_X1 U439 ( .A(n385), .B(n384), .ZN(n391) );
  XOR2_X1 U440 ( .A(n387), .B(n386), .Z(n389) );
  NAND2_X1 U441 ( .A1(G232GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U442 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U443 ( .A(n391), .B(n390), .Z(n397) );
  XOR2_X1 U444 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n393) );
  XNOR2_X1 U445 ( .A(G162GAT), .B(KEYINPUT80), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U448 ( .A(n397), .B(n396), .ZN(n465) );
  XOR2_X1 U449 ( .A(n398), .B(G78GAT), .Z(n401) );
  XNOR2_X1 U450 ( .A(G155GAT), .B(n399), .ZN(n400) );
  XNOR2_X1 U451 ( .A(n401), .B(n400), .ZN(n406) );
  XOR2_X1 U452 ( .A(KEYINPUT12), .B(n402), .Z(n404) );
  NAND2_X1 U453 ( .A1(G231GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U454 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U455 ( .A(n406), .B(n405), .Z(n414) );
  XOR2_X1 U456 ( .A(G64GAT), .B(G183GAT), .Z(n408) );
  XNOR2_X1 U457 ( .A(G57GAT), .B(G211GAT), .ZN(n407) );
  XNOR2_X1 U458 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U459 ( .A(KEYINPUT15), .B(KEYINPUT83), .Z(n410) );
  XNOR2_X1 U460 ( .A(KEYINPUT14), .B(KEYINPUT84), .ZN(n409) );
  XNOR2_X1 U461 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U462 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U463 ( .A(n414), .B(n413), .ZN(n561) );
  NAND2_X1 U464 ( .A1(n465), .A2(n561), .ZN(n415) );
  XNOR2_X1 U465 ( .A(KEYINPUT47), .B(n417), .ZN(n423) );
  XOR2_X1 U466 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n419) );
  XOR2_X1 U467 ( .A(KEYINPUT36), .B(n465), .Z(n577) );
  INV_X1 U468 ( .A(n561), .ZN(n575) );
  NAND2_X1 U469 ( .A1(n577), .A2(n575), .ZN(n418) );
  XNOR2_X1 U470 ( .A(n419), .B(n418), .ZN(n420) );
  NOR2_X1 U471 ( .A1(n571), .A2(n420), .ZN(n421) );
  NAND2_X1 U472 ( .A1(n565), .A2(n421), .ZN(n422) );
  NAND2_X1 U473 ( .A1(n423), .A2(n422), .ZN(n424) );
  XOR2_X1 U474 ( .A(KEYINPUT48), .B(n424), .Z(n523) );
  NOR2_X1 U475 ( .A1(n512), .A2(n523), .ZN(n425) );
  XOR2_X1 U476 ( .A(n425), .B(KEYINPUT54), .Z(n426) );
  NOR2_X1 U477 ( .A1(n496), .A2(n426), .ZN(n564) );
  NAND2_X1 U478 ( .A1(n460), .A2(n564), .ZN(n427) );
  XNOR2_X1 U479 ( .A(n427), .B(KEYINPUT55), .ZN(n442) );
  XOR2_X1 U480 ( .A(G190GAT), .B(n428), .Z(n430) );
  NAND2_X1 U481 ( .A1(G227GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U483 ( .A(G176GAT), .B(KEYINPUT20), .Z(n432) );
  XNOR2_X1 U484 ( .A(G15GAT), .B(G71GAT), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U486 ( .A(n434), .B(n433), .Z(n439) );
  XOR2_X1 U487 ( .A(G99GAT), .B(G43GAT), .Z(n436) );
  XNOR2_X1 U488 ( .A(G120GAT), .B(G127GAT), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U490 ( .A(G134GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n525) );
  NAND2_X1 U493 ( .A1(n442), .A2(n525), .ZN(n560) );
  NOR2_X1 U494 ( .A1(n565), .A2(n560), .ZN(n445) );
  INV_X1 U495 ( .A(KEYINPUT122), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n443), .B(G169GAT), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(G1348GAT) );
  NOR2_X1 U498 ( .A1(n465), .A2(n560), .ZN(n448) );
  INV_X1 U499 ( .A(n496), .ZN(n510) );
  NOR2_X1 U500 ( .A1(n565), .A2(n571), .ZN(n482) );
  NAND2_X1 U501 ( .A1(n499), .A2(n525), .ZN(n449) );
  XNOR2_X1 U502 ( .A(KEYINPUT100), .B(n449), .ZN(n450) );
  NAND2_X1 U503 ( .A1(n450), .A2(n460), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n451), .B(KEYINPUT25), .ZN(n455) );
  XNOR2_X1 U505 ( .A(n499), .B(KEYINPUT27), .ZN(n452) );
  XOR2_X1 U506 ( .A(n452), .B(KEYINPUT99), .Z(n459) );
  OR2_X1 U507 ( .A1(n460), .A2(n525), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n453), .B(KEYINPUT26), .ZN(n540) );
  INV_X1 U509 ( .A(n540), .ZN(n563) );
  AND2_X1 U510 ( .A1(n459), .A2(n563), .ZN(n454) );
  NOR2_X1 U511 ( .A1(n455), .A2(n454), .ZN(n456) );
  NOR2_X1 U512 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n458), .B(KEYINPUT101), .ZN(n464) );
  NAND2_X1 U514 ( .A1(n496), .A2(n459), .ZN(n522) );
  XNOR2_X1 U515 ( .A(KEYINPUT28), .B(KEYINPUT66), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n461), .B(n460), .ZN(n526) );
  INV_X1 U517 ( .A(n526), .ZN(n503) );
  NOR2_X1 U518 ( .A1(n522), .A2(n503), .ZN(n462) );
  INV_X1 U519 ( .A(n525), .ZN(n515) );
  NAND2_X1 U520 ( .A1(n462), .A2(n515), .ZN(n463) );
  NAND2_X1 U521 ( .A1(n464), .A2(n463), .ZN(n478) );
  INV_X1 U522 ( .A(n465), .ZN(n551) );
  NOR2_X1 U523 ( .A1(n551), .A2(n561), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(KEYINPUT85), .ZN(n467) );
  XOR2_X1 U525 ( .A(KEYINPUT16), .B(n467), .Z(n468) );
  AND2_X1 U526 ( .A1(n478), .A2(n468), .ZN(n494) );
  NAND2_X1 U527 ( .A1(n482), .A2(n494), .ZN(n476) );
  NOR2_X1 U528 ( .A1(n510), .A2(n476), .ZN(n469) );
  XOR2_X1 U529 ( .A(G1GAT), .B(n469), .Z(n470) );
  XNOR2_X1 U530 ( .A(KEYINPUT34), .B(n470), .ZN(G1324GAT) );
  NOR2_X1 U531 ( .A1(n512), .A2(n476), .ZN(n471) );
  XOR2_X1 U532 ( .A(G8GAT), .B(n471), .Z(G1325GAT) );
  NOR2_X1 U533 ( .A1(n476), .A2(n515), .ZN(n475) );
  XOR2_X1 U534 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n473) );
  XNOR2_X1 U535 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n472) );
  XNOR2_X1 U536 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U537 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  NOR2_X1 U538 ( .A1(n526), .A2(n476), .ZN(n477) );
  XOR2_X1 U539 ( .A(G22GAT), .B(n477), .Z(G1327GAT) );
  NAND2_X1 U540 ( .A1(n561), .A2(n478), .ZN(n479) );
  XOR2_X1 U541 ( .A(KEYINPUT104), .B(n479), .Z(n480) );
  NAND2_X1 U542 ( .A1(n480), .A2(n577), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n481), .B(KEYINPUT37), .ZN(n509) );
  NAND2_X1 U544 ( .A1(n482), .A2(n509), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n483), .B(KEYINPUT38), .ZN(n491) );
  NOR2_X1 U546 ( .A1(n510), .A2(n491), .ZN(n486) );
  XOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT105), .Z(n484) );
  XNOR2_X1 U548 ( .A(KEYINPUT39), .B(n484), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  NOR2_X1 U550 ( .A1(n491), .A2(n512), .ZN(n487) );
  XOR2_X1 U551 ( .A(G36GAT), .B(n487), .Z(G1329GAT) );
  XNOR2_X1 U552 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n489) );
  NOR2_X1 U553 ( .A1(n515), .A2(n491), .ZN(n488) );
  XNOR2_X1 U554 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U555 ( .A(G43GAT), .B(n490), .Z(G1330GAT) );
  XNOR2_X1 U556 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n493) );
  NOR2_X1 U557 ( .A1(n526), .A2(n491), .ZN(n492) );
  XNOR2_X1 U558 ( .A(n493), .B(n492), .ZN(G1331GAT) );
  XNOR2_X1 U559 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n498) );
  INV_X1 U560 ( .A(n565), .ZN(n542) );
  NOR2_X1 U561 ( .A1(n554), .A2(n542), .ZN(n508) );
  NAND2_X1 U562 ( .A1(n508), .A2(n494), .ZN(n495) );
  XOR2_X1 U563 ( .A(KEYINPUT108), .B(n495), .Z(n504) );
  NAND2_X1 U564 ( .A1(n496), .A2(n504), .ZN(n497) );
  XNOR2_X1 U565 ( .A(n498), .B(n497), .ZN(G1332GAT) );
  XOR2_X1 U566 ( .A(G64GAT), .B(KEYINPUT109), .Z(n501) );
  NAND2_X1 U567 ( .A1(n499), .A2(n504), .ZN(n500) );
  XNOR2_X1 U568 ( .A(n501), .B(n500), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n504), .A2(n525), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n502), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n506) );
  NAND2_X1 U572 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(n507), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n509), .A2(n508), .ZN(n519) );
  NOR2_X1 U576 ( .A1(n510), .A2(n519), .ZN(n511) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n511), .Z(G1336GAT) );
  NOR2_X1 U578 ( .A1(n512), .A2(n519), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1337GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n519), .ZN(n516) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n516), .Z(G1338GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n518) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(KEYINPUT113), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n521) );
  NOR2_X1 U586 ( .A1(n526), .A2(n519), .ZN(n520) );
  XOR2_X1 U587 ( .A(n521), .B(n520), .Z(G1339GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n529) );
  NOR2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(KEYINPUT115), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U592 ( .A1(n539), .A2(n527), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n536), .A2(n542), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n532) );
  INV_X1 U597 ( .A(n554), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n536), .A2(n545), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G120GAT), .B(n533), .ZN(G1341GAT) );
  NAND2_X1 U601 ( .A1(n575), .A2(n536), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U605 ( .A1(n536), .A2(n551), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U608 ( .A(KEYINPUT119), .B(n541), .Z(n552) );
  NAND2_X1 U609 ( .A1(n542), .A2(n552), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n543), .B(KEYINPUT120), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n547) );
  NAND2_X1 U613 ( .A1(n552), .A2(n545), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n548), .ZN(G1345GAT) );
  XOR2_X1 U616 ( .A(G155GAT), .B(KEYINPUT121), .Z(n550) );
  NAND2_X1 U617 ( .A1(n552), .A2(n575), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n553), .ZN(G1347GAT) );
  NOR2_X1 U621 ( .A1(n554), .A2(n560), .ZN(n559) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(KEYINPUT56), .B(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(G183GAT), .B(n562), .Z(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n570) );
  NOR2_X1 U630 ( .A1(n565), .A2(n570), .ZN(n567) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n573) );
  INV_X1 U636 ( .A(n570), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n578), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(n574), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n578), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n580) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

