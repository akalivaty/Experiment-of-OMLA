//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n599, new_n600, new_n601,
    new_n603, new_n604, new_n605, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n643, new_n646,
    new_n647, new_n649, new_n650, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1240, new_n1241, new_n1242;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n460), .A2(new_n461), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n459), .A2(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(KEYINPUT67), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n459), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n479), .A2(KEYINPUT68), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT69), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2105), .B1(new_n476), .B2(new_n478), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n489), .B1(new_n491), .B2(G124), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  OAI21_X1  g072(.A(G2105), .B1(new_n497), .B2(G114), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(KEYINPUT70), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n460), .B2(new_n461), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n506), .B1(new_n460), .B2(new_n461), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n506), .B(new_n509), .C1(new_n461), .C2(new_n460), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n504), .B1(new_n508), .B2(new_n510), .ZN(G164));
  AND2_X1   g086(.A1(KEYINPUT72), .A2(KEYINPUT6), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT72), .A2(KEYINPUT6), .ZN(new_n513));
  OAI21_X1  g088(.A(G651), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g091(.A(KEYINPUT73), .B(G651), .C1(new_n512), .C2(new_n513), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT71), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n520), .A2(new_n522), .A3(KEYINPUT6), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n518), .A2(G50), .A3(G543), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT74), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n523), .B1(new_n516), .B2(new_n517), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n527), .A2(new_n528), .A3(G50), .A4(G543), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n520), .A2(new_n522), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G62), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT75), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT5), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n537), .A2(KEYINPUT76), .ZN(new_n538));
  NAND2_X1  g113(.A1(G75), .A2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n539), .B1(new_n537), .B2(KEYINPUT76), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n531), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n535), .A2(new_n536), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n527), .A2(G88), .A3(new_n542), .ZN(new_n543));
  AND4_X1   g118(.A1(new_n526), .A2(new_n529), .A3(new_n541), .A4(new_n543), .ZN(G166));
  NAND3_X1  g119(.A1(new_n527), .A2(G51), .A3(G543), .ZN(new_n545));
  AND3_X1   g120(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n546));
  AOI21_X1  g121(.A(KEYINPUT5), .B1(KEYINPUT75), .B2(G543), .ZN(new_n547));
  OAI21_X1  g122(.A(KEYINPUT77), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n535), .A2(new_n549), .A3(new_n536), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n551), .A2(G63), .A3(G651), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n518), .A2(G89), .A3(new_n524), .A4(new_n542), .ZN(new_n554));
  NAND3_X1  g129(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT7), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT78), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n554), .A2(new_n559), .A3(new_n556), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n553), .B1(new_n558), .B2(new_n560), .ZN(G168));
  NAND2_X1  g136(.A1(new_n551), .A2(G64), .ZN(new_n562));
  NAND2_X1  g137(.A1(G77), .A2(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n530), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n518), .A2(G52), .A3(G543), .A4(new_n524), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n518), .A2(G90), .A3(new_n524), .A4(new_n542), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT79), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n565), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n564), .B1(new_n568), .B2(new_n570), .ZN(G171));
  NAND3_X1  g146(.A1(new_n548), .A2(new_n550), .A3(G56), .ZN(new_n572));
  INV_X1    g147(.A(G68), .ZN(new_n573));
  INV_X1    g148(.A(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(new_n531), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n527), .A2(G81), .A3(new_n542), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n527), .A2(G43), .A3(G543), .ZN(new_n578));
  AND3_X1   g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G860), .ZN(G153));
  NAND4_X1  g155(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g156(.A1(G1), .A2(G3), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT8), .ZN(new_n583));
  NAND4_X1  g158(.A1(G319), .A2(G483), .A3(G661), .A4(new_n583), .ZN(G188));
  INV_X1    g159(.A(G53), .ZN(new_n585));
  NOR3_X1   g160(.A1(new_n585), .A2(new_n574), .A3(KEYINPUT80), .ZN(new_n586));
  XNOR2_X1  g161(.A(KEYINPUT72), .B(KEYINPUT6), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT73), .B1(new_n587), .B2(G651), .ZN(new_n588));
  INV_X1    g163(.A(new_n517), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n524), .B(new_n586), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT9), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n542), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n519), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n518), .A2(G91), .A3(new_n524), .A4(new_n542), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n518), .A2(KEYINPUT9), .A3(new_n524), .A4(new_n586), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n592), .A2(new_n595), .A3(new_n596), .A4(new_n597), .ZN(G299));
  INV_X1    g173(.A(new_n564), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n565), .A2(new_n566), .A3(new_n569), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n569), .B1(new_n565), .B2(new_n566), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(G301));
  INV_X1    g177(.A(new_n553), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n554), .A2(new_n559), .A3(new_n556), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n559), .B1(new_n554), .B2(new_n556), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(G286));
  NAND4_X1  g181(.A1(new_n526), .A2(new_n529), .A3(new_n541), .A4(new_n543), .ZN(G303));
  NAND3_X1  g182(.A1(new_n527), .A2(G87), .A3(new_n542), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n518), .A2(G49), .A3(G543), .A4(new_n524), .ZN(new_n609));
  OAI21_X1  g184(.A(G651), .B1(new_n551), .B2(G74), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(G288));
  NAND4_X1  g186(.A1(new_n518), .A2(G86), .A3(new_n524), .A4(new_n542), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n518), .A2(G48), .A3(G543), .A4(new_n524), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n542), .A2(G61), .ZN(new_n614));
  AND2_X1   g189(.A1(G73), .A2(G543), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n531), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n612), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT81), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n612), .A2(new_n613), .A3(new_n619), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(G305));
  XOR2_X1   g197(.A(KEYINPUT82), .B(G47), .Z(new_n623));
  NAND3_X1  g198(.A1(new_n527), .A2(G543), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n548), .A2(new_n550), .A3(G60), .ZN(new_n625));
  NAND2_X1  g200(.A1(G72), .A2(G543), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n531), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n518), .A2(G85), .A3(new_n524), .A4(new_n542), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n624), .A2(new_n628), .A3(new_n629), .ZN(G290));
  NAND4_X1  g205(.A1(new_n518), .A2(G92), .A3(new_n524), .A4(new_n542), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT10), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n633));
  NAND4_X1  g208(.A1(new_n527), .A2(new_n633), .A3(G92), .A4(new_n542), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n542), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(new_n519), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n527), .A2(G54), .A3(G543), .ZN(new_n637));
  NAND4_X1  g212(.A1(new_n632), .A2(new_n634), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(G868), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G171), .B2(new_n639), .ZN(G284));
  OAI21_X1  g216(.A(new_n640), .B1(G171), .B2(new_n639), .ZN(G321));
  NAND2_X1  g217(.A1(G299), .A2(new_n639), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(G168), .B2(new_n639), .ZN(G297));
  OAI21_X1  g219(.A(new_n643), .B1(G168), .B2(new_n639), .ZN(G280));
  INV_X1    g220(.A(new_n638), .ZN(new_n646));
  INV_X1    g221(.A(G559), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n647), .B2(G860), .ZN(G148));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G868), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(G868), .B2(new_n579), .ZN(G323));
  XNOR2_X1  g226(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g227(.A1(new_n477), .A2(new_n467), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT84), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT13), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n658), .A2(G2100), .ZN(new_n659));
  INV_X1    g234(.A(G123), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n459), .A2(G111), .ZN(new_n661));
  OAI21_X1  g236(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n662));
  OAI22_X1  g237(.A1(new_n490), .A2(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n484), .B2(G135), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n665), .A2(G2096), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n658), .A2(G2100), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(G2096), .ZN(new_n668));
  NAND4_X1  g243(.A1(new_n659), .A2(new_n666), .A3(new_n667), .A4(new_n668), .ZN(G156));
  XNOR2_X1  g244(.A(G2427), .B(G2438), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2430), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT15), .B(G2435), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(KEYINPUT14), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2443), .B(G2446), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1341), .B(G1348), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT86), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2451), .B(G2454), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT16), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT85), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n680), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(G14), .A3(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G401));
  INV_X1    g262(.A(KEYINPUT18), .ZN(new_n688));
  XOR2_X1   g263(.A(G2084), .B(G2090), .Z(new_n689));
  XNOR2_X1  g264(.A(G2067), .B(G2678), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(KEYINPUT17), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n689), .A2(new_n690), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n688), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G2096), .B(G2100), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G2072), .B(G2078), .Z(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n691), .B2(KEYINPUT18), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT87), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n696), .B(new_n699), .ZN(G227));
  XOR2_X1   g275(.A(G1971), .B(G1976), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT19), .ZN(new_n702));
  XOR2_X1   g277(.A(G1956), .B(G2474), .Z(new_n703));
  XOR2_X1   g278(.A(G1961), .B(G1966), .Z(new_n704));
  AND2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT20), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n703), .A2(new_n704), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n702), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n702), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n711), .B(new_n712), .Z(new_n713));
  XNOR2_X1  g288(.A(G1991), .B(G1996), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT88), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1981), .B(G1986), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n713), .A2(new_n715), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n713), .A2(new_n715), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n720), .A2(new_n717), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n722), .ZN(G229));
  NOR2_X1   g298(.A1(G16), .A2(G22), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G166), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1971), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT33), .B(G1976), .Z(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G23), .ZN(new_n729));
  AND3_X1   g304(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n728), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT89), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n726), .B1(new_n727), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n728), .A2(G6), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n621), .B2(new_n728), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT32), .B(G1981), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n732), .A2(new_n727), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n733), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(KEYINPUT34), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(KEYINPUT34), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n484), .A2(G131), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(G107), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G2105), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n491), .B2(G119), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  MUX2_X1   g322(.A(G25), .B(new_n747), .S(G29), .Z(new_n748));
  XOR2_X1   g323(.A(KEYINPUT35), .B(G1991), .Z(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n748), .B(new_n750), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n728), .A2(G24), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G290), .B2(G16), .ZN(new_n753));
  INV_X1    g328(.A(G1986), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n751), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n740), .A2(new_n741), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(KEYINPUT90), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(KEYINPUT90), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n758), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n740), .A2(new_n760), .A3(new_n741), .A4(new_n757), .ZN(new_n764));
  INV_X1    g339(.A(G29), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n765), .A2(G35), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n493), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT29), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n767), .A2(new_n768), .ZN(new_n771));
  OAI21_X1  g346(.A(G2090), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n771), .ZN(new_n773));
  INV_X1    g348(.A(G2090), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n773), .A2(new_n774), .A3(new_n769), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT26), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n467), .A2(G105), .ZN(new_n779));
  INV_X1    g354(.A(G129), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n778), .B(new_n779), .C1(new_n490), .C2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n484), .B2(G141), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(new_n765), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n765), .B2(G32), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT27), .B(G1996), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n765), .A2(G27), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT94), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n497), .A2(G114), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n499), .A2(KEYINPUT70), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n789), .A2(new_n790), .A3(G2105), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n791), .A2(new_n496), .B1(new_n477), .B2(new_n502), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n509), .B1(new_n477), .B2(new_n506), .ZN(new_n793));
  INV_X1    g368(.A(new_n510), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n788), .B1(new_n795), .B2(G29), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT95), .Z(new_n797));
  INV_X1    g372(.A(G2078), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  INV_X1    g375(.A(G28), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT30), .ZN(new_n802));
  AOI21_X1  g377(.A(G29), .B1(new_n801), .B2(KEYINPUT30), .ZN(new_n803));
  OR2_X1    g378(.A1(KEYINPUT31), .A2(G11), .ZN(new_n804));
  NAND2_X1  g379(.A1(KEYINPUT31), .A2(G11), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n802), .A2(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G34), .ZN(new_n807));
  AOI21_X1  g382(.A(G29), .B1(new_n807), .B2(KEYINPUT24), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(KEYINPUT24), .B2(new_n807), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n473), .B2(new_n765), .ZN(new_n810));
  INV_X1    g385(.A(G2084), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n664), .B2(G29), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n786), .A2(new_n799), .A3(new_n800), .A4(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G2072), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n765), .A2(G33), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n484), .A2(G139), .ZN(new_n817));
  NAND2_X1  g392(.A1(G115), .A2(G2104), .ZN(new_n818));
  INV_X1    g393(.A(G127), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n469), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT25), .ZN(new_n821));
  NAND2_X1  g396(.A1(G103), .A2(G2104), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(G2105), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n459), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n820), .A2(G2105), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT91), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n816), .B1(new_n827), .B2(G29), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n814), .B1(new_n815), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n728), .A2(G21), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G168), .B2(new_n728), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(G1966), .Z(new_n832));
  OR2_X1    g407(.A1(new_n828), .A2(new_n815), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n728), .A2(G20), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT23), .Z(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G299), .B2(G16), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1956), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n829), .A2(new_n832), .A3(new_n833), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n810), .A2(new_n811), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT92), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n728), .A2(G5), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G171), .B2(new_n728), .ZN(new_n842));
  OAI221_X1 g417(.A(new_n840), .B1(G1961), .B2(new_n842), .C1(new_n784), .C2(new_n785), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT93), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n765), .A2(G26), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT28), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n484), .A2(G140), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n850));
  INV_X1    g425(.A(G116), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n851), .B2(G2105), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n491), .B2(G128), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n848), .B1(new_n854), .B2(G29), .ZN(new_n855));
  INV_X1    g430(.A(G2067), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n728), .A2(G4), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n646), .B2(new_n728), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(G1348), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n579), .A2(G16), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(G16), .B2(G19), .ZN(new_n862));
  INV_X1    g437(.A(G1341), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  NOR4_X1   g440(.A1(new_n857), .A2(new_n860), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n842), .A2(G1961), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n845), .A2(new_n846), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n776), .A2(new_n838), .A3(new_n868), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n763), .A2(new_n764), .A3(new_n869), .ZN(G311));
  NAND3_X1  g445(.A1(new_n763), .A2(new_n869), .A3(new_n764), .ZN(G150));
  NAND3_X1  g446(.A1(new_n548), .A2(new_n550), .A3(G67), .ZN(new_n872));
  NAND2_X1  g447(.A1(G80), .A2(G543), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n531), .ZN(new_n875));
  XOR2_X1   g450(.A(KEYINPUT97), .B(G93), .Z(new_n876));
  NAND4_X1  g451(.A1(new_n518), .A2(new_n524), .A3(new_n542), .A4(new_n876), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n518), .A2(G55), .A3(G543), .A4(new_n524), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(KEYINPUT99), .B(G860), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT37), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n638), .A2(new_n647), .ZN(new_n884));
  XOR2_X1   g459(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n879), .A2(KEYINPUT98), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n875), .A2(new_n877), .A3(new_n878), .A4(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n579), .A2(new_n880), .A3(new_n889), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n886), .B(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT39), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n895), .A2(new_n896), .A3(new_n881), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n896), .B1(new_n895), .B2(new_n881), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n883), .B1(new_n897), .B2(new_n898), .ZN(G145));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n747), .B(new_n656), .ZN(new_n901));
  OR2_X1    g476(.A1(G106), .A2(G2105), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n902), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n903));
  INV_X1    g478(.A(G130), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(new_n490), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n905), .B1(new_n484), .B2(G142), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n901), .B(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n849), .A2(KEYINPUT101), .A3(new_n853), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n910));
  INV_X1    g485(.A(G140), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(new_n482), .B2(new_n483), .ZN(new_n912));
  INV_X1    g487(.A(new_n853), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n909), .A2(new_n914), .A3(new_n795), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n795), .B1(new_n909), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n782), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n909), .A2(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(G164), .ZN(new_n919));
  INV_X1    g494(.A(new_n782), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n909), .A2(new_n914), .A3(new_n795), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n917), .A2(new_n922), .A3(new_n827), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n826), .B1(new_n917), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n908), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n826), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n915), .A2(new_n916), .A3(new_n782), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n901), .B(new_n906), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n917), .A2(new_n922), .A3(new_n827), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n664), .B(new_n473), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n493), .B(new_n933), .Z(new_n934));
  NAND3_X1  g509(.A1(new_n925), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G37), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n934), .B1(new_n925), .B2(new_n932), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n900), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n938), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n940), .A2(KEYINPUT40), .A3(new_n936), .A4(new_n935), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n939), .A2(new_n941), .ZN(G395));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(new_n879), .B2(new_n639), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n893), .B(new_n649), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n638), .A2(G299), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT41), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n638), .A2(G299), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n947), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n950), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n638), .A2(G299), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT41), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n955), .A3(KEYINPUT103), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n946), .A2(new_n951), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n947), .A2(new_n950), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n891), .A2(new_n892), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(new_n649), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n621), .A2(G166), .ZN(new_n965));
  NAND3_X1  g540(.A1(G303), .A2(new_n618), .A3(new_n620), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(G290), .A2(G288), .ZN(new_n968));
  NOR2_X1   g543(.A1(G290), .A2(G288), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT104), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT104), .B1(new_n968), .B2(new_n969), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n628), .A2(new_n629), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n730), .A2(new_n624), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n975));
  NAND2_X1  g550(.A1(G290), .A2(G288), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n972), .A2(new_n977), .A3(new_n965), .A4(new_n966), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n971), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT42), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n639), .B1(new_n964), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n957), .A2(new_n963), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n979), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n945), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n980), .A2(new_n963), .A3(new_n957), .ZN(new_n987));
  AND4_X1   g562(.A1(new_n943), .A2(new_n987), .A3(new_n985), .A4(G868), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n986), .A2(new_n988), .ZN(G295));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n985), .A3(G868), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n944), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT106), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n991), .B(new_n992), .C1(KEYINPUT105), .C2(new_n990), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT106), .B1(new_n986), .B2(new_n988), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(G331));
  NAND2_X1  g570(.A1(G171), .A2(G168), .ZN(new_n996));
  NAND2_X1  g571(.A1(G301), .A2(G286), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(new_n961), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n996), .A2(new_n997), .B1(new_n892), .B2(new_n891), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n956), .B(new_n951), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT107), .B1(new_n998), .B2(new_n961), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n958), .B1(new_n998), .B2(new_n961), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n893), .A2(new_n1004), .A3(new_n997), .A4(new_n996), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n979), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1001), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n998), .A2(new_n961), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1002), .A2(new_n1009), .A3(new_n1005), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n954), .A2(new_n955), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n999), .A2(new_n1000), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1010), .A2(new_n1011), .B1(new_n1012), .B2(new_n960), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n979), .A2(KEYINPUT108), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n971), .A2(new_n978), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n936), .B(new_n1008), .C1(new_n1013), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT43), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1008), .A2(new_n936), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1012), .A2(new_n960), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1017), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT110), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1020), .A2(new_n1027), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n936), .B(new_n1008), .C1(new_n1029), .C2(new_n1017), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT44), .B1(new_n1030), .B2(KEYINPUT43), .ZN(new_n1031));
  NOR2_X1   g606(.A1(KEYINPUT43), .A2(G37), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1026), .A2(KEYINPUT109), .A3(new_n1008), .A4(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1017), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1008), .A2(new_n1032), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1033), .A2(new_n1037), .B1(KEYINPUT43), .B2(new_n1030), .ZN(new_n1038));
  OAI22_X1  g613(.A1(new_n1028), .A2(new_n1031), .B1(new_n1038), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g614(.A1(new_n920), .A2(G1996), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n854), .A2(G2067), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n849), .A2(new_n856), .A3(new_n853), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1384), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n795), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(KEYINPUT111), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT45), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n508), .A2(new_n510), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1384), .B1(new_n1049), .B2(new_n792), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G40), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n464), .A2(new_n471), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1044), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(G1996), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT113), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(new_n920), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT114), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n1062));
  OAI221_X1 g637(.A(new_n1062), .B1(new_n1059), .B2(new_n920), .C1(new_n1056), .C2(new_n1044), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1056), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n747), .A2(new_n750), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n749), .B1(new_n742), .B2(new_n746), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n973), .A2(new_n754), .A3(new_n624), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G290), .A2(G1986), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(KEYINPUT112), .A3(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1064), .B(new_n1070), .C1(KEYINPUT112), .C2(new_n1069), .ZN(new_n1071));
  AND4_X1   g646(.A1(new_n1061), .A2(new_n1063), .A3(new_n1067), .A4(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1055), .B1(new_n1050), .B2(KEYINPUT45), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n795), .A2(KEYINPUT45), .A3(new_n1045), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1046), .A2(KEYINPUT50), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT50), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1050), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1079), .A3(new_n1055), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1076), .A2(G1966), .B1(new_n1080), .B2(G2084), .ZN(new_n1081));
  OAI21_X1  g656(.A(G8), .B1(new_n1081), .B2(G286), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1081), .A2(G286), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT51), .B1(new_n1084), .B2(new_n1082), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT53), .B1(new_n1076), .B2(new_n798), .ZN(new_n1087));
  INV_X1    g662(.A(G1961), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n1080), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1076), .A2(KEYINPUT53), .A3(new_n798), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(G301), .B(KEYINPUT54), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1092), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT125), .B(G2078), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1055), .A2(KEYINPUT53), .A3(new_n1095), .ZN(new_n1096));
  OR3_X1    g671(.A1(new_n1053), .A2(new_n1075), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(new_n1089), .A3(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1086), .A2(new_n1093), .A3(new_n1098), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n617), .A2(G1981), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n617), .A2(G1981), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT49), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1100), .A2(KEYINPUT49), .A3(new_n1101), .ZN(new_n1105));
  INV_X1    g680(.A(G8), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n730), .A2(G1976), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT117), .B(G1976), .Z(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT52), .B1(G288), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(new_n1111), .A3(new_n1107), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1109), .A2(new_n1107), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1108), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(G303), .A2(G8), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT115), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(KEYINPUT55), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1120));
  NAND3_X1  g695(.A1(G303), .A2(G8), .A3(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1076), .A2(G1971), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1055), .B1(new_n1050), .B2(new_n1078), .ZN(new_n1124));
  AOI211_X1 g699(.A(KEYINPUT50), .B(G1384), .C1(new_n1049), .C2(new_n792), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n774), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1106), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1122), .A2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1119), .A2(KEYINPUT116), .A3(new_n1121), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT116), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1128), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1116), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1122), .A2(new_n1128), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1136), .A2(new_n1108), .A3(new_n1115), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(KEYINPUT126), .A3(new_n1132), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1099), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT118), .B(G1956), .Z(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1048), .B1(G164), .B2(G1384), .ZN(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT56), .B(G2072), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1142), .A2(new_n1055), .A3(new_n1074), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n546), .A2(new_n547), .ZN(new_n1147));
  AOI211_X1 g722(.A(new_n1147), .B(new_n523), .C1(new_n516), .C2(new_n517), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n594), .B1(new_n1148), .B2(G91), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(new_n592), .A4(new_n597), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1146), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1145), .A2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1146), .A2(new_n1151), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT119), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1141), .A2(new_n1146), .A3(new_n1151), .A4(new_n1144), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT119), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1153), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(KEYINPUT123), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1145), .A2(new_n1152), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1154), .A2(new_n1155), .A3(KEYINPUT119), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1163), .B1(new_n1167), .B2(KEYINPUT61), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n465), .A2(G40), .A3(new_n472), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1169), .B1(new_n1046), .B2(KEYINPUT50), .ZN(new_n1170));
  AOI21_X1  g745(.A(G1348), .B1(new_n1170), .B2(new_n1079), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1055), .A2(new_n1045), .A3(new_n795), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1172), .A2(G2067), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1174), .A2(KEYINPUT60), .A3(new_n638), .ZN(new_n1175));
  XNOR2_X1  g750(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(G1341), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT122), .ZN(new_n1179));
  INV_X1    g754(.A(G1996), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1142), .A2(new_n1180), .A3(new_n1055), .A4(new_n1074), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1172), .A2(new_n1182), .A3(new_n1177), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1179), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT59), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1184), .A2(new_n1185), .A3(new_n579), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1185), .B1(new_n1184), .B2(new_n579), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1175), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1153), .A2(KEYINPUT61), .A3(new_n1157), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT60), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1190), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1173), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1192), .B(KEYINPUT60), .C1(new_n1126), .C2(G1348), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1191), .A2(new_n1193), .A3(new_n646), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1189), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1188), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1162), .A2(new_n1168), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1153), .B1(new_n638), .B2(new_n1174), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1198), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(KEYINPUT120), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT120), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1198), .B(new_n1201), .C1(new_n1156), .C2(new_n1159), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1197), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1197), .A2(KEYINPUT124), .A3(new_n1203), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1139), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  AND3_X1   g783(.A1(new_n1081), .A2(G8), .A3(G168), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1116), .A2(new_n1129), .A3(new_n1132), .A4(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT63), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1137), .A2(KEYINPUT63), .A3(new_n1132), .A4(new_n1209), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NOR3_X1   g789(.A1(new_n1132), .A2(new_n1108), .A3(new_n1115), .ZN(new_n1215));
  OR2_X1    g790(.A1(G288), .A2(G1976), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1100), .B1(new_n1108), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1215), .B1(new_n1107), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1138), .A2(new_n1135), .ZN(new_n1219));
  AND3_X1   g794(.A1(new_n1083), .A2(new_n1085), .A3(KEYINPUT62), .ZN(new_n1220));
  AOI21_X1  g795(.A(KEYINPUT62), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1221));
  OAI211_X1 g796(.A(G171), .B(new_n1091), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g797(.A(new_n1214), .B(new_n1218), .C1(new_n1219), .C2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1072), .B1(new_n1208), .B2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1056), .A2(new_n1068), .ZN(new_n1225));
  XOR2_X1   g800(.A(new_n1225), .B(KEYINPUT48), .Z(new_n1226));
  NAND4_X1  g801(.A1(new_n1061), .A2(new_n1063), .A3(new_n1067), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1056), .B1(new_n1043), .B2(new_n782), .ZN(new_n1228));
  XNOR2_X1  g803(.A(new_n1228), .B(KEYINPUT127), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n1059), .B(KEYINPUT46), .ZN(new_n1230));
  INV_X1    g805(.A(KEYINPUT47), .ZN(new_n1231));
  AND3_X1   g806(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1231), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1227), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g809(.A1(new_n1061), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1056), .B1(new_n1235), .B2(new_n1042), .ZN(new_n1236));
  NOR2_X1   g811(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1224), .A2(new_n1237), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g813(.A1(G227), .A2(new_n457), .ZN(new_n1240));
  NOR3_X1   g814(.A1(G229), .A2(G401), .A3(new_n1240), .ZN(new_n1241));
  OAI21_X1  g815(.A(new_n1241), .B1(new_n937), .B2(new_n938), .ZN(new_n1242));
  NOR2_X1   g816(.A1(new_n1242), .A2(new_n1038), .ZN(G308));
  OR2_X1    g817(.A1(new_n1242), .A2(new_n1038), .ZN(G225));
endmodule


