

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U322 ( .A(G8GAT), .B(G92GAT), .Z(n290) );
  XOR2_X1 U323 ( .A(n394), .B(KEYINPUT90), .Z(n291) );
  INV_X1 U324 ( .A(KEYINPUT25), .ZN(n413) );
  XNOR2_X1 U325 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U326 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U327 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U328 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U329 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U330 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U331 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n465) );
  XNOR2_X1 U332 ( .A(n466), .B(n465), .ZN(n534) );
  XNOR2_X1 U333 ( .A(n342), .B(n290), .ZN(n300) );
  XNOR2_X1 U334 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U335 ( .A(n453), .B(KEYINPUT41), .Z(n554) );
  INV_X1 U336 ( .A(G36GAT), .ZN(n444) );
  XNOR2_X1 U337 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U338 ( .A(n444), .B(KEYINPUT102), .ZN(n445) );
  XNOR2_X1 U339 ( .A(n475), .B(n474), .ZN(G1349GAT) );
  XNOR2_X1 U340 ( .A(n446), .B(n445), .ZN(G1329GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n293) );
  XNOR2_X1 U342 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U344 ( .A(G169GAT), .B(n294), .Z(n356) );
  XOR2_X1 U345 ( .A(KEYINPUT74), .B(G64GAT), .Z(n296) );
  XNOR2_X1 U346 ( .A(G176GAT), .B(G204GAT), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n329) );
  XNOR2_X1 U348 ( .A(n356), .B(n329), .ZN(n303) );
  XOR2_X1 U349 ( .A(G211GAT), .B(KEYINPUT21), .Z(n298) );
  XNOR2_X1 U350 ( .A(G197GAT), .B(G218GAT), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n394) );
  NAND2_X1 U352 ( .A1(G226GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n291), .B(n299), .ZN(n301) );
  XOR2_X1 U354 ( .A(G36GAT), .B(G190GAT), .Z(n342) );
  XOR2_X1 U355 ( .A(n303), .B(n302), .Z(n526) );
  INV_X1 U356 ( .A(n526), .ZN(n493) );
  XNOR2_X1 U357 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n304), .B(G8GAT), .ZN(n435) );
  XOR2_X1 U359 ( .A(G141GAT), .B(G22GAT), .Z(n401) );
  XOR2_X1 U360 ( .A(n435), .B(n401), .Z(n306) );
  XNOR2_X1 U361 ( .A(G36GAT), .B(G50GAT), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n312) );
  XOR2_X1 U363 ( .A(G29GAT), .B(G43GAT), .Z(n308) );
  XNOR2_X1 U364 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n308), .B(n307), .ZN(n343) );
  XOR2_X1 U366 ( .A(n343), .B(KEYINPUT30), .Z(n310) );
  NAND2_X1 U367 ( .A1(G229GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U369 ( .A(n312), .B(n311), .Z(n320) );
  XOR2_X1 U370 ( .A(G113GAT), .B(G15GAT), .Z(n314) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(G197GAT), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U373 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n316) );
  XNOR2_X1 U374 ( .A(KEYINPUT68), .B(KEYINPUT66), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U377 ( .A(n320), .B(n319), .Z(n512) );
  INV_X1 U378 ( .A(n512), .ZN(n572) );
  XOR2_X1 U379 ( .A(KEYINPUT72), .B(G92GAT), .Z(n322) );
  XNOR2_X1 U380 ( .A(G99GAT), .B(KEYINPUT71), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U382 ( .A(G85GAT), .B(n323), .Z(n350) );
  XOR2_X1 U383 ( .A(KEYINPUT32), .B(KEYINPUT77), .Z(n325) );
  NAND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U386 ( .A(n326), .B(KEYINPUT33), .Z(n331) );
  XOR2_X1 U387 ( .A(G78GAT), .B(G148GAT), .Z(n328) );
  XNOR2_X1 U388 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n398) );
  XNOR2_X1 U390 ( .A(n398), .B(n329), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n337) );
  XOR2_X1 U392 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n333) );
  XNOR2_X1 U393 ( .A(KEYINPUT31), .B(KEYINPUT76), .ZN(n332) );
  XOR2_X1 U394 ( .A(n333), .B(n332), .Z(n335) );
  XOR2_X1 U395 ( .A(G120GAT), .B(G71GAT), .Z(n359) );
  XOR2_X1 U396 ( .A(G57GAT), .B(KEYINPUT13), .Z(n426) );
  XNOR2_X1 U397 ( .A(n359), .B(n426), .ZN(n334) );
  XOR2_X1 U398 ( .A(n350), .B(n338), .Z(n447) );
  NAND2_X1 U399 ( .A1(n572), .A2(n447), .ZN(n489) );
  XOR2_X1 U400 ( .A(KEYINPUT64), .B(G106GAT), .Z(n340) );
  XNOR2_X1 U401 ( .A(G134GAT), .B(G218GAT), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U403 ( .A(n342), .B(n341), .Z(n345) );
  XOR2_X1 U404 ( .A(G50GAT), .B(G162GAT), .Z(n400) );
  XNOR2_X1 U405 ( .A(n343), .B(n400), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U407 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n347) );
  NAND2_X1 U408 ( .A1(G232GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U410 ( .A(n349), .B(n348), .Z(n352) );
  XNOR2_X1 U411 ( .A(n350), .B(KEYINPUT9), .ZN(n351) );
  XOR2_X1 U412 ( .A(n352), .B(n351), .Z(n483) );
  XNOR2_X1 U413 ( .A(KEYINPUT36), .B(n483), .ZN(n479) );
  XOR2_X1 U414 ( .A(KEYINPUT81), .B(G134GAT), .Z(n354) );
  XNOR2_X1 U415 ( .A(KEYINPUT80), .B(KEYINPUT0), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U417 ( .A(G113GAT), .B(n355), .Z(n384) );
  XNOR2_X1 U418 ( .A(n384), .B(n356), .ZN(n367) );
  XOR2_X1 U419 ( .A(G176GAT), .B(KEYINPUT20), .Z(n358) );
  XNOR2_X1 U420 ( .A(G43GAT), .B(KEYINPUT82), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n363) );
  XOR2_X1 U422 ( .A(G190GAT), .B(G99GAT), .Z(n361) );
  XOR2_X1 U423 ( .A(G15GAT), .B(G127GAT), .Z(n427) );
  XNOR2_X1 U424 ( .A(n427), .B(n359), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U426 ( .A(n363), .B(n362), .Z(n365) );
  NAND2_X1 U427 ( .A1(G227GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U429 ( .A(n367), .B(n366), .Z(n535) );
  INV_X1 U430 ( .A(n535), .ZN(n504) );
  XOR2_X1 U431 ( .A(G148GAT), .B(G120GAT), .Z(n369) );
  XNOR2_X1 U432 ( .A(G1GAT), .B(G127GAT), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U434 ( .A(G85GAT), .B(G162GAT), .Z(n371) );
  XNOR2_X1 U435 ( .A(G29GAT), .B(G141GAT), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U437 ( .A(n373), .B(n372), .ZN(n388) );
  XOR2_X1 U438 ( .A(KEYINPUT89), .B(KEYINPUT5), .Z(n375) );
  XNOR2_X1 U439 ( .A(G57GAT), .B(KEYINPUT88), .ZN(n374) );
  XNOR2_X1 U440 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U441 ( .A(KEYINPUT6), .B(KEYINPUT86), .Z(n377) );
  XNOR2_X1 U442 ( .A(KEYINPUT4), .B(KEYINPUT87), .ZN(n376) );
  XNOR2_X1 U443 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U444 ( .A(n379), .B(n378), .Z(n386) );
  XNOR2_X1 U445 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n380), .B(KEYINPUT2), .ZN(n395) );
  XOR2_X1 U447 ( .A(n395), .B(KEYINPUT1), .Z(n382) );
  NAND2_X1 U448 ( .A1(G225GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U449 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U452 ( .A(n388), .B(n387), .Z(n550) );
  INV_X1 U453 ( .A(n550), .ZN(n500) );
  XOR2_X1 U454 ( .A(n526), .B(KEYINPUT27), .Z(n410) );
  XOR2_X1 U455 ( .A(G204GAT), .B(KEYINPUT83), .Z(n390) );
  XNOR2_X1 U456 ( .A(KEYINPUT23), .B(KEYINPUT85), .ZN(n389) );
  XNOR2_X1 U457 ( .A(n390), .B(n389), .ZN(n405) );
  XOR2_X1 U458 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n392) );
  NAND2_X1 U459 ( .A1(G228GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U461 ( .A(n393), .B(KEYINPUT84), .Z(n397) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n397), .B(n396), .ZN(n399) );
  XOR2_X1 U464 ( .A(n399), .B(n398), .Z(n403) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U466 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n469) );
  XNOR2_X1 U468 ( .A(KEYINPUT28), .B(n469), .ZN(n530) );
  OR2_X1 U469 ( .A1(n410), .A2(n530), .ZN(n406) );
  NOR2_X1 U470 ( .A1(n500), .A2(n406), .ZN(n536) );
  NAND2_X1 U471 ( .A1(n504), .A2(n536), .ZN(n407) );
  XNOR2_X1 U472 ( .A(n407), .B(KEYINPUT91), .ZN(n420) );
  NAND2_X1 U473 ( .A1(n469), .A2(n504), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n408), .B(KEYINPUT26), .ZN(n409) );
  XNOR2_X1 U475 ( .A(KEYINPUT92), .B(n409), .ZN(n476) );
  NOR2_X1 U476 ( .A1(n476), .A2(n410), .ZN(n551) );
  NOR2_X1 U477 ( .A1(n504), .A2(n493), .ZN(n411) );
  XOR2_X1 U478 ( .A(KEYINPUT93), .B(n411), .Z(n412) );
  NOR2_X1 U479 ( .A1(n469), .A2(n412), .ZN(n416) );
  XOR2_X1 U480 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n414) );
  NOR2_X1 U481 ( .A1(n551), .A2(n417), .ZN(n418) );
  NOR2_X1 U482 ( .A1(n550), .A2(n418), .ZN(n419) );
  NOR2_X1 U483 ( .A1(n420), .A2(n419), .ZN(n421) );
  XNOR2_X1 U484 ( .A(KEYINPUT96), .B(n421), .ZN(n487) );
  NOR2_X1 U485 ( .A1(n479), .A2(n487), .ZN(n440) );
  XOR2_X1 U486 ( .A(G78GAT), .B(G71GAT), .Z(n423) );
  XNOR2_X1 U487 ( .A(G22GAT), .B(G183GAT), .ZN(n422) );
  XNOR2_X1 U488 ( .A(n423), .B(n422), .ZN(n439) );
  XOR2_X1 U489 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n425) );
  XNOR2_X1 U490 ( .A(KEYINPUT12), .B(KEYINPUT79), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n431) );
  XOR2_X1 U492 ( .A(n426), .B(G211GAT), .Z(n429) );
  XNOR2_X1 U493 ( .A(n427), .B(G155GAT), .ZN(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U495 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U496 ( .A1(G231GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U498 ( .A(n434), .B(G64GAT), .Z(n437) );
  XNOR2_X1 U499 ( .A(n435), .B(KEYINPUT14), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n582) );
  INV_X1 U502 ( .A(n582), .ZN(n484) );
  NAND2_X1 U503 ( .A1(n440), .A2(n484), .ZN(n441) );
  XOR2_X1 U504 ( .A(KEYINPUT37), .B(n441), .Z(n524) );
  NOR2_X1 U505 ( .A1(n489), .A2(n524), .ZN(n443) );
  XNOR2_X1 U506 ( .A(KEYINPUT101), .B(KEYINPUT38), .ZN(n442) );
  XNOR2_X1 U507 ( .A(n443), .B(n442), .ZN(n509) );
  NOR2_X1 U508 ( .A1(n493), .A2(n509), .ZN(n446) );
  INV_X1 U509 ( .A(n447), .ZN(n453) );
  XOR2_X1 U510 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n449) );
  NOR2_X1 U511 ( .A1(n479), .A2(n484), .ZN(n448) );
  XOR2_X1 U512 ( .A(n449), .B(n448), .Z(n450) );
  NOR2_X1 U513 ( .A1(n453), .A2(n450), .ZN(n451) );
  XNOR2_X1 U514 ( .A(n451), .B(KEYINPUT111), .ZN(n452) );
  NOR2_X1 U515 ( .A1(n572), .A2(n452), .ZN(n464) );
  NAND2_X1 U516 ( .A1(n572), .A2(n554), .ZN(n455) );
  INV_X1 U517 ( .A(KEYINPUT46), .ZN(n454) );
  XNOR2_X1 U518 ( .A(n455), .B(n454), .ZN(n456) );
  NOR2_X1 U519 ( .A1(n582), .A2(n456), .ZN(n457) );
  XNOR2_X1 U520 ( .A(n457), .B(KEYINPUT108), .ZN(n458) );
  AND2_X1 U521 ( .A1(n458), .A2(n483), .ZN(n462) );
  XOR2_X1 U522 ( .A(KEYINPUT47), .B(KEYINPUT109), .Z(n460) );
  INV_X1 U523 ( .A(KEYINPUT110), .ZN(n459) );
  NOR2_X1 U524 ( .A1(n464), .A2(n463), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n534), .A2(n493), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n467), .B(KEYINPUT54), .ZN(n468) );
  NAND2_X1 U527 ( .A1(n468), .A2(n500), .ZN(n477) );
  NOR2_X1 U528 ( .A1(n477), .A2(n469), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(KEYINPUT55), .ZN(n471) );
  NOR2_X2 U530 ( .A1(n504), .A2(n471), .ZN(n567) );
  NAND2_X1 U531 ( .A1(n567), .A2(n554), .ZN(n475) );
  XOR2_X1 U532 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n473) );
  XNOR2_X1 U533 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n472) );
  INV_X1 U534 ( .A(G218GAT), .ZN(n482) );
  NOR2_X1 U535 ( .A1(n477), .A2(n476), .ZN(n583) );
  INV_X1 U536 ( .A(n583), .ZN(n478) );
  NOR2_X1 U537 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U538 ( .A(KEYINPUT62), .B(n480), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(G1355GAT) );
  INV_X1 U540 ( .A(n483), .ZN(n566) );
  NOR2_X1 U541 ( .A1(n566), .A2(n484), .ZN(n485) );
  XOR2_X1 U542 ( .A(KEYINPUT16), .B(n485), .Z(n486) );
  NOR2_X1 U543 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U544 ( .A(KEYINPUT97), .B(n488), .ZN(n513) );
  NOR2_X1 U545 ( .A1(n513), .A2(n489), .ZN(n490) );
  XOR2_X1 U546 ( .A(KEYINPUT98), .B(n490), .Z(n497) );
  NOR2_X1 U547 ( .A1(n500), .A2(n497), .ZN(n491) );
  XOR2_X1 U548 ( .A(n491), .B(KEYINPUT34), .Z(n492) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n492), .ZN(G1324GAT) );
  NOR2_X1 U550 ( .A1(n493), .A2(n497), .ZN(n494) );
  XOR2_X1 U551 ( .A(G8GAT), .B(n494), .Z(G1325GAT) );
  XNOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n496) );
  NOR2_X1 U553 ( .A1(n504), .A2(n497), .ZN(n495) );
  XNOR2_X1 U554 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  INV_X1 U555 ( .A(n530), .ZN(n508) );
  NOR2_X1 U556 ( .A1(n497), .A2(n508), .ZN(n499) );
  XNOR2_X1 U557 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(G1327GAT) );
  XNOR2_X1 U559 ( .A(KEYINPUT100), .B(KEYINPUT39), .ZN(n502) );
  NOR2_X1 U560 ( .A1(n500), .A2(n509), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(n503), .ZN(G1328GAT) );
  XNOR2_X1 U563 ( .A(KEYINPUT103), .B(KEYINPUT40), .ZN(n506) );
  NOR2_X1 U564 ( .A1(n504), .A2(n509), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NOR2_X1 U567 ( .A1(n509), .A2(n508), .ZN(n510) );
  XOR2_X1 U568 ( .A(KEYINPUT104), .B(n510), .Z(n511) );
  XNOR2_X1 U569 ( .A(G50GAT), .B(n511), .ZN(G1331GAT) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n515) );
  NAND2_X1 U571 ( .A1(n512), .A2(n554), .ZN(n523) );
  NOR2_X1 U572 ( .A1(n513), .A2(n523), .ZN(n519) );
  NAND2_X1 U573 ( .A1(n519), .A2(n550), .ZN(n514) );
  XNOR2_X1 U574 ( .A(n515), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n519), .A2(n526), .ZN(n516) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n516), .ZN(G1333GAT) );
  XOR2_X1 U577 ( .A(G71GAT), .B(KEYINPUT105), .Z(n518) );
  NAND2_X1 U578 ( .A1(n519), .A2(n535), .ZN(n517) );
  XNOR2_X1 U579 ( .A(n518), .B(n517), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U581 ( .A1(n519), .A2(n530), .ZN(n520) );
  XNOR2_X1 U582 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(n522), .ZN(G1335GAT) );
  NOR2_X1 U584 ( .A1(n524), .A2(n523), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n531), .A2(n550), .ZN(n525) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n526), .A2(n531), .ZN(n527) );
  XNOR2_X1 U588 ( .A(n527), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U589 ( .A(G99GAT), .B(KEYINPUT107), .Z(n529) );
  NAND2_X1 U590 ( .A1(n531), .A2(n535), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n529), .B(n528), .ZN(G1338GAT) );
  NAND2_X1 U592 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U593 ( .A(n532), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NAND2_X1 U595 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n534), .A2(n537), .ZN(n546) );
  NAND2_X1 U597 ( .A1(n546), .A2(n572), .ZN(n538) );
  XNOR2_X1 U598 ( .A(n538), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U600 ( .A1(n546), .A2(n554), .ZN(n539) );
  XNOR2_X1 U601 ( .A(n540), .B(n539), .ZN(n542) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT113), .Z(n541) );
  XNOR2_X1 U603 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n544) );
  NAND2_X1 U605 ( .A1(n546), .A2(n582), .ZN(n543) );
  XNOR2_X1 U606 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n548) );
  NAND2_X1 U609 ( .A1(n546), .A2(n566), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U613 ( .A1(n534), .A2(n552), .ZN(n560) );
  NAND2_X1 U614 ( .A1(n560), .A2(n572), .ZN(n553) );
  XNOR2_X1 U615 ( .A(n553), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n556) );
  NAND2_X1 U617 ( .A1(n560), .A2(n554), .ZN(n555) );
  XNOR2_X1 U618 ( .A(n556), .B(n555), .ZN(n558) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .Z(n557) );
  XNOR2_X1 U620 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n582), .A2(n560), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n560), .A2(n566), .ZN(n561) );
  XNOR2_X1 U624 ( .A(n561), .B(KEYINPUT118), .ZN(n562) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n562), .ZN(G1347GAT) );
  XOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT119), .Z(n564) );
  NAND2_X1 U627 ( .A1(n567), .A2(n572), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n564), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n582), .A2(n567), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n568) );
  XNOR2_X1 U633 ( .A(n569), .B(n568), .ZN(n571) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(G1351GAT) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n583), .A2(n572), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n583), .A2(n453), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  XOR2_X1 U647 ( .A(G211GAT), .B(KEYINPUT127), .Z(n585) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1354GAT) );
endmodule

