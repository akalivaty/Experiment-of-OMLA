

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760;

  XNOR2_X1 U375 ( .A(n421), .B(n419), .ZN(n675) );
  NAND2_X1 U376 ( .A1(n385), .A2(n384), .ZN(n524) );
  NOR2_X1 U377 ( .A1(n756), .A2(n758), .ZN(n546) );
  AND2_X1 U378 ( .A1(n374), .A2(n599), .ZN(n355) );
  XNOR2_X1 U379 ( .A(n355), .B(KEYINPUT33), .ZN(n672) );
  INV_X1 U380 ( .A(G953), .ZN(n748) );
  XNOR2_X2 U381 ( .A(n544), .B(KEYINPUT115), .ZN(n556) );
  XNOR2_X2 U382 ( .A(G116), .B(G119), .ZN(n370) );
  NOR2_X2 U383 ( .A1(n692), .A2(n691), .ZN(n698) );
  OR2_X2 U384 ( .A1(n605), .A2(n606), .ZN(n428) );
  NOR2_X2 U385 ( .A1(n631), .A2(G902), .ZN(n503) );
  XNOR2_X2 U386 ( .A(n378), .B(KEYINPUT101), .ZN(n650) );
  XNOR2_X2 U387 ( .A(n503), .B(n502), .ZN(n567) );
  AND2_X1 U388 ( .A1(n376), .A2(n375), .ZN(n641) );
  NAND2_X1 U389 ( .A1(n401), .A2(n404), .ZN(n624) );
  OR2_X1 U390 ( .A1(n601), .A2(n600), .ZN(n432) );
  XNOR2_X1 U391 ( .A(n536), .B(n417), .ZN(n577) );
  INV_X1 U392 ( .A(n563), .ZN(n611) );
  NOR2_X1 U393 ( .A1(n552), .A2(n692), .ZN(n429) );
  XNOR2_X1 U394 ( .A(n524), .B(n440), .ZN(n631) );
  XNOR2_X1 U395 ( .A(n479), .B(n478), .ZN(n527) );
  XNOR2_X1 U396 ( .A(n500), .B(G125), .ZN(n485) );
  XNOR2_X1 U397 ( .A(G101), .B(KEYINPUT3), .ZN(n478) );
  INV_X1 U398 ( .A(G146), .ZN(n500) );
  XNOR2_X2 U399 ( .A(n540), .B(KEYINPUT41), .ZN(n688) );
  AND2_X1 U400 ( .A1(n759), .A2(KEYINPUT44), .ZN(n400) );
  NOR2_X1 U401 ( .A1(n650), .A2(n666), .ZN(n616) );
  AND2_X1 U402 ( .A1(n676), .A2(n675), .ZN(n680) );
  INV_X1 U403 ( .A(G134), .ZN(n462) );
  NAND2_X1 U404 ( .A1(n598), .A2(n354), .ZN(n408) );
  NOR2_X1 U405 ( .A1(n562), .A2(n561), .ZN(n570) );
  AND2_X1 U406 ( .A1(n403), .A2(n402), .ZN(n401) );
  OR2_X1 U407 ( .A1(G237), .A2(G902), .ZN(n522) );
  XOR2_X1 U408 ( .A(KEYINPUT94), .B(G140), .Z(n491) );
  XNOR2_X1 U409 ( .A(G101), .B(G104), .ZN(n490) );
  INV_X1 U410 ( .A(n372), .ZN(n423) );
  XNOR2_X1 U411 ( .A(G902), .B(KEYINPUT15), .ZN(n626) );
  OR2_X1 U412 ( .A1(n598), .A2(KEYINPUT113), .ZN(n405) );
  XNOR2_X1 U413 ( .A(n457), .B(n456), .ZN(n549) );
  NOR2_X1 U414 ( .A1(G902), .A2(n722), .ZN(n457) );
  XOR2_X1 U415 ( .A(G110), .B(G137), .Z(n515) );
  XNOR2_X1 U416 ( .A(G119), .B(G128), .ZN(n514) );
  XNOR2_X1 U417 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U418 ( .A(KEYINPUT70), .B(KEYINPUT24), .Z(n510) );
  XNOR2_X1 U419 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n508) );
  XNOR2_X1 U420 ( .A(n485), .B(n422), .ZN(n744) );
  XNOR2_X1 U421 ( .A(KEYINPUT10), .B(G140), .ZN(n422) );
  XNOR2_X1 U422 ( .A(n734), .B(n433), .ZN(n637) );
  XNOR2_X1 U423 ( .A(n434), .B(n484), .ZN(n433) );
  XNOR2_X1 U424 ( .A(n371), .B(n486), .ZN(n434) );
  XNOR2_X1 U425 ( .A(n418), .B(KEYINPUT39), .ZN(n417) );
  INV_X1 U426 ( .A(KEYINPUT71), .ZN(n418) );
  INV_X1 U427 ( .A(KEYINPUT36), .ZN(n398) );
  XNOR2_X1 U428 ( .A(n380), .B(n597), .ZN(n601) );
  NAND2_X1 U429 ( .A1(n613), .A2(n595), .ZN(n380) );
  XNOR2_X1 U430 ( .A(n411), .B(n410), .ZN(n600) );
  INV_X1 U431 ( .A(KEYINPUT79), .ZN(n410) );
  NAND2_X1 U432 ( .A1(n406), .A2(n405), .ZN(n411) );
  AND2_X1 U433 ( .A1(n408), .A2(n407), .ZN(n406) );
  INV_X1 U434 ( .A(n549), .ZN(n558) );
  NOR2_X1 U435 ( .A1(n609), .A2(n608), .ZN(n365) );
  XNOR2_X1 U436 ( .A(n563), .B(KEYINPUT6), .ZN(n599) );
  XNOR2_X1 U437 ( .A(n521), .B(n420), .ZN(n419) );
  OR2_X1 U438 ( .A1(n730), .A2(G902), .ZN(n421) );
  INV_X1 U439 ( .A(KEYINPUT25), .ZN(n420) );
  NAND2_X1 U440 ( .A1(n622), .A2(KEYINPUT86), .ZN(n381) );
  XNOR2_X1 U441 ( .A(G131), .B(KEYINPUT4), .ZN(n495) );
  XNOR2_X1 U442 ( .A(KEYINPUT48), .B(KEYINPUT85), .ZN(n576) );
  XOR2_X1 U443 ( .A(KEYINPUT97), .B(KEYINPUT23), .Z(n509) );
  XNOR2_X1 U444 ( .A(n485), .B(n435), .ZN(n371) );
  XNOR2_X1 U445 ( .A(n487), .B(n436), .ZN(n435) );
  INV_X1 U446 ( .A(KEYINPUT4), .ZN(n436) );
  AND2_X1 U447 ( .A1(n428), .A2(n607), .ZN(n404) );
  NAND2_X1 U448 ( .A1(G234), .A2(G237), .ZN(n473) );
  NAND2_X1 U449 ( .A1(n399), .A2(n395), .ZN(n394) );
  NOR2_X1 U450 ( .A1(n409), .A2(n599), .ZN(n407) );
  XNOR2_X1 U451 ( .A(n488), .B(n489), .ZN(n552) );
  XNOR2_X1 U452 ( .A(G116), .B(G107), .ZN(n463) );
  XOR2_X1 U453 ( .A(KEYINPUT7), .B(G122), .Z(n464) );
  XOR2_X1 U454 ( .A(n494), .B(n493), .Z(n440) );
  XNOR2_X1 U455 ( .A(n492), .B(n439), .ZN(n493) );
  XNOR2_X1 U456 ( .A(n679), .B(n568), .ZN(n598) );
  AND2_X1 U457 ( .A1(n599), .A2(n390), .ZN(n565) );
  INV_X1 U458 ( .A(n564), .ZN(n390) );
  INV_X1 U459 ( .A(KEYINPUT0), .ZN(n373) );
  BUF_X1 U460 ( .A(n552), .Z(n580) );
  AND2_X1 U461 ( .A1(n533), .A2(n534), .ZN(n547) );
  XNOR2_X1 U462 ( .A(n437), .B(n481), .ZN(n734) );
  XNOR2_X1 U463 ( .A(n527), .B(n480), .ZN(n437) );
  XNOR2_X1 U464 ( .A(n519), .B(n518), .ZN(n730) );
  XNOR2_X1 U465 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U466 ( .A(n744), .B(n512), .ZN(n519) );
  BUF_X1 U467 ( .A(n720), .Z(n728) );
  XNOR2_X1 U468 ( .A(n538), .B(KEYINPUT116), .ZN(n756) );
  XNOR2_X1 U469 ( .A(n416), .B(n537), .ZN(n538) );
  XNOR2_X1 U470 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n424) );
  INV_X1 U471 ( .A(n593), .ZN(n426) );
  XNOR2_X1 U472 ( .A(n431), .B(KEYINPUT78), .ZN(n430) );
  INV_X1 U473 ( .A(KEYINPUT32), .ZN(n431) );
  BUF_X1 U474 ( .A(G146), .Z(n372) );
  NOR2_X1 U475 ( .A1(n611), .A2(n602), .ZN(n655) );
  NOR2_X1 U476 ( .A1(n558), .A2(n557), .ZN(n663) );
  OR2_X1 U477 ( .A1(n610), .A2(n611), .ZN(n378) );
  XNOR2_X1 U478 ( .A(n365), .B(n364), .ZN(n610) );
  INV_X1 U479 ( .A(KEYINPUT100), .ZN(n364) );
  AND2_X1 U480 ( .A1(n619), .A2(n360), .ZN(n621) );
  INV_X1 U481 ( .A(KEYINPUT60), .ZN(n368) );
  OR2_X1 U482 ( .A1(n661), .A2(n692), .ZN(n353) );
  AND2_X1 U483 ( .A1(n620), .A2(KEYINPUT113), .ZN(n354) );
  AND2_X1 U484 ( .A1(n759), .A2(n604), .ZN(n356) );
  NOR2_X1 U485 ( .A1(n661), .A2(n394), .ZN(n393) );
  AND2_X1 U486 ( .A1(n460), .A2(G134), .ZN(n357) );
  AND2_X1 U487 ( .A1(n582), .A2(n671), .ZN(n358) );
  NAND2_X1 U488 ( .A1(n393), .A2(KEYINPUT36), .ZN(n359) );
  AND2_X1 U489 ( .A1(n618), .A2(n675), .ZN(n360) );
  XOR2_X1 U490 ( .A(n591), .B(KEYINPUT34), .Z(n361) );
  XOR2_X1 U491 ( .A(n639), .B(n638), .Z(n362) );
  XOR2_X1 U492 ( .A(n722), .B(n721), .Z(n363) );
  INV_X1 U493 ( .A(n732), .ZN(n375) );
  NAND2_X2 U494 ( .A1(n414), .A2(n358), .ZN(n747) );
  NAND2_X1 U495 ( .A1(n547), .A2(n535), .ZN(n536) );
  NOR2_X1 U496 ( .A1(n392), .A2(n391), .ZN(n397) );
  NOR2_X1 U497 ( .A1(n709), .A2(n625), .ZN(n627) );
  NOR2_X2 U498 ( .A1(n712), .A2(n747), .ZN(n709) );
  XNOR2_X2 U499 ( .A(n366), .B(n530), .ZN(n643) );
  XNOR2_X2 U500 ( .A(n524), .B(G113), .ZN(n366) );
  NAND2_X1 U501 ( .A1(n367), .A2(n567), .ZN(n544) );
  XNOR2_X1 U502 ( .A(n543), .B(KEYINPUT28), .ZN(n367) );
  XNOR2_X1 U503 ( .A(n369), .B(n368), .ZN(G60) );
  NAND2_X1 U504 ( .A1(n724), .A2(n375), .ZN(n369) );
  NAND2_X1 U505 ( .A1(n577), .A2(n663), .ZN(n416) );
  INV_X1 U506 ( .A(n370), .ZN(n479) );
  XNOR2_X1 U507 ( .A(n429), .B(n555), .ZN(n588) );
  INV_X1 U508 ( .A(n613), .ZN(n609) );
  XNOR2_X2 U509 ( .A(n590), .B(n373), .ZN(n613) );
  INV_X1 U510 ( .A(n599), .ZN(n618) );
  INV_X1 U511 ( .A(n612), .ZN(n374) );
  XNOR2_X1 U512 ( .A(n640), .B(n362), .ZN(n376) );
  NOR2_X2 U513 ( .A1(n377), .A2(n574), .ZN(n575) );
  NAND2_X1 U514 ( .A1(n573), .A2(n572), .ZN(n377) );
  INV_X1 U515 ( .A(n611), .ZN(n379) );
  XNOR2_X1 U516 ( .A(n592), .B(n361), .ZN(n427) );
  NAND2_X1 U517 ( .A1(n382), .A2(n381), .ZN(n403) );
  NAND2_X1 U518 ( .A1(n588), .A2(n589), .ZN(n590) );
  NAND2_X1 U519 ( .A1(n400), .A2(n622), .ZN(n382) );
  NOR2_X2 U520 ( .A1(n643), .A2(G902), .ZN(n531) );
  XNOR2_X1 U521 ( .A(n383), .B(n648), .ZN(G57) );
  NOR2_X2 U522 ( .A1(n646), .A2(n732), .ZN(n383) );
  NAND2_X1 U523 ( .A1(n427), .A2(n426), .ZN(n425) );
  NAND2_X1 U524 ( .A1(n746), .A2(n372), .ZN(n384) );
  NAND2_X1 U525 ( .A1(n386), .A2(n423), .ZN(n385) );
  INV_X1 U526 ( .A(n746), .ZN(n386) );
  XNOR2_X2 U527 ( .A(n499), .B(n498), .ZN(n746) );
  XNOR2_X2 U528 ( .A(n387), .B(n576), .ZN(n414) );
  NAND2_X1 U529 ( .A1(n388), .A2(n415), .ZN(n387) );
  XNOR2_X1 U530 ( .A(n575), .B(n389), .ZN(n388) );
  INV_X1 U531 ( .A(KEYINPUT67), .ZN(n389) );
  XNOR2_X2 U532 ( .A(n531), .B(G472), .ZN(n563) );
  NOR2_X1 U533 ( .A1(n393), .A2(KEYINPUT36), .ZN(n391) );
  AND2_X1 U534 ( .A1(n566), .A2(n398), .ZN(n392) );
  INV_X1 U535 ( .A(n692), .ZN(n395) );
  NAND2_X1 U536 ( .A1(n397), .A2(n396), .ZN(n569) );
  OR2_X1 U537 ( .A1(n359), .A2(n566), .ZN(n396) );
  OR2_X1 U538 ( .A1(n566), .A2(n353), .ZN(n578) );
  INV_X1 U539 ( .A(n580), .ZN(n399) );
  NOR2_X1 U540 ( .A1(n356), .A2(n617), .ZN(n402) );
  NOR2_X1 U541 ( .A1(n620), .A2(KEYINPUT113), .ZN(n409) );
  NAND2_X1 U542 ( .A1(n461), .A2(n460), .ZN(n482) );
  NAND2_X1 U543 ( .A1(n357), .A2(n461), .ZN(n413) );
  NAND2_X2 U544 ( .A1(n413), .A2(n412), .ZN(n498) );
  NAND2_X1 U545 ( .A1(n482), .A2(n462), .ZN(n412) );
  XNOR2_X1 U546 ( .A(n546), .B(KEYINPUT46), .ZN(n415) );
  XNOR2_X2 U547 ( .A(n425), .B(n424), .ZN(n759) );
  XNOR2_X2 U548 ( .A(n432), .B(n430), .ZN(n757) );
  XNOR2_X1 U549 ( .A(n635), .B(n634), .ZN(n636) );
  AND2_X1 U550 ( .A1(n636), .A2(n375), .ZN(G54) );
  AND2_X1 U551 ( .A1(G227), .A2(n748), .ZN(n439) );
  NOR2_X1 U552 ( .A1(G952), .A2(n748), .ZN(n732) );
  INV_X1 U553 ( .A(n480), .ZN(n443) );
  XNOR2_X1 U554 ( .A(n443), .B(n444), .ZN(n445) );
  XNOR2_X1 U555 ( .A(n744), .B(n445), .ZN(n453) );
  XNOR2_X1 U556 ( .A(n527), .B(n526), .ZN(n529) );
  XNOR2_X1 U557 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U558 ( .A(n501), .B(G469), .ZN(n502) );
  INV_X1 U559 ( .A(KEYINPUT77), .ZN(n553) );
  XNOR2_X1 U560 ( .A(n554), .B(n553), .ZN(n555) );
  INV_X1 U561 ( .A(KEYINPUT89), .ZN(n568) );
  XNOR2_X1 U562 ( .A(n647), .B(KEYINPUT63), .ZN(n648) );
  INV_X1 U563 ( .A(KEYINPUT40), .ZN(n537) );
  NOR2_X1 U564 ( .A1(G237), .A2(G953), .ZN(n441) );
  XNOR2_X1 U565 ( .A(n441), .B(KEYINPUT76), .ZN(n525) );
  NAND2_X1 U566 ( .A1(G214), .A2(n525), .ZN(n444) );
  XNOR2_X1 U567 ( .A(G113), .B(G122), .ZN(n442) );
  XNOR2_X1 U568 ( .A(n442), .B(G104), .ZN(n480) );
  XOR2_X1 U569 ( .A(KEYINPUT103), .B(KEYINPUT11), .Z(n447) );
  XNOR2_X1 U570 ( .A(G143), .B(KEYINPUT12), .ZN(n446) );
  XNOR2_X1 U571 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U572 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n449) );
  XNOR2_X1 U573 ( .A(G131), .B(KEYINPUT106), .ZN(n448) );
  XNOR2_X1 U574 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U575 ( .A(n451), .B(n450), .Z(n452) );
  XNOR2_X1 U576 ( .A(n453), .B(n452), .ZN(n722) );
  XOR2_X1 U577 ( .A(KEYINPUT108), .B(KEYINPUT13), .Z(n455) );
  XNOR2_X1 U578 ( .A(KEYINPUT107), .B(G475), .ZN(n454) );
  XNOR2_X1 U579 ( .A(n455), .B(n454), .ZN(n456) );
  INV_X1 U580 ( .A(G128), .ZN(n458) );
  NAND2_X1 U581 ( .A1(G143), .A2(n458), .ZN(n461) );
  INV_X1 U582 ( .A(G143), .ZN(n459) );
  NAND2_X1 U583 ( .A1(n459), .A2(G128), .ZN(n460) );
  XNOR2_X1 U584 ( .A(n464), .B(n463), .ZN(n465) );
  XOR2_X1 U585 ( .A(n498), .B(n465), .Z(n468) );
  NAND2_X1 U586 ( .A1(G234), .A2(n748), .ZN(n466) );
  XOR2_X1 U587 ( .A(KEYINPUT8), .B(n466), .Z(n513) );
  NAND2_X1 U588 ( .A1(G217), .A2(n513), .ZN(n467) );
  XNOR2_X1 U589 ( .A(n468), .B(n467), .ZN(n470) );
  XOR2_X1 U590 ( .A(KEYINPUT9), .B(KEYINPUT109), .Z(n469) );
  XNOR2_X1 U591 ( .A(n470), .B(n469), .ZN(n726) );
  NOR2_X1 U592 ( .A1(G902), .A2(n726), .ZN(n472) );
  XOR2_X1 U593 ( .A(KEYINPUT110), .B(G478), .Z(n471) );
  XNOR2_X1 U594 ( .A(n472), .B(n471), .ZN(n557) );
  XNOR2_X1 U595 ( .A(n473), .B(KEYINPUT14), .ZN(n474) );
  NAND2_X1 U596 ( .A1(G952), .A2(n474), .ZN(n707) );
  NOR2_X1 U597 ( .A1(G953), .A2(n707), .ZN(n583) );
  NAND2_X1 U598 ( .A1(n474), .A2(G902), .ZN(n475) );
  XOR2_X1 U599 ( .A(KEYINPUT92), .B(n475), .Z(n584) );
  NAND2_X1 U600 ( .A1(n584), .A2(G953), .ZN(n476) );
  NOR2_X1 U601 ( .A1(G900), .A2(n476), .ZN(n477) );
  NOR2_X1 U602 ( .A1(n583), .A2(n477), .ZN(n541) );
  INV_X1 U603 ( .A(n541), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n522), .A2(G210), .ZN(n489) );
  XOR2_X1 U605 ( .A(G107), .B(G110), .Z(n492) );
  XNOR2_X1 U606 ( .A(n492), .B(KEYINPUT16), .ZN(n481) );
  XNOR2_X1 U607 ( .A(n482), .B(KEYINPUT88), .ZN(n483) );
  XNOR2_X1 U608 ( .A(n483), .B(KEYINPUT17), .ZN(n484) );
  AND2_X1 U609 ( .A1(G224), .A2(n748), .ZN(n486) );
  INV_X1 U610 ( .A(KEYINPUT18), .ZN(n487) );
  NAND2_X1 U611 ( .A1(n637), .A2(n626), .ZN(n488) );
  XNOR2_X1 U612 ( .A(KEYINPUT38), .B(n580), .ZN(n539) );
  AND2_X1 U613 ( .A1(n548), .A2(n539), .ZN(n535) );
  XNOR2_X1 U614 ( .A(n491), .B(n490), .ZN(n494) );
  INV_X1 U615 ( .A(n495), .ZN(n497) );
  XNOR2_X1 U616 ( .A(KEYINPUT66), .B(G137), .ZN(n496) );
  XNOR2_X1 U617 ( .A(n497), .B(n496), .ZN(n499) );
  XNOR2_X1 U618 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n501) );
  XOR2_X1 U619 ( .A(KEYINPUT21), .B(KEYINPUT98), .Z(n506) );
  NAND2_X1 U620 ( .A1(n626), .A2(G234), .ZN(n504) );
  XNOR2_X1 U621 ( .A(n504), .B(KEYINPUT20), .ZN(n520) );
  NAND2_X1 U622 ( .A1(G221), .A2(n520), .ZN(n505) );
  XNOR2_X1 U623 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U624 ( .A(KEYINPUT99), .B(n507), .Z(n676) );
  XNOR2_X1 U625 ( .A(n509), .B(n508), .ZN(n511) );
  NAND2_X1 U626 ( .A1(n513), .A2(G221), .ZN(n517) );
  XNOR2_X1 U627 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U628 ( .A1(G217), .A2(n520), .ZN(n521) );
  NAND2_X1 U629 ( .A1(n567), .A2(n680), .ZN(n608) );
  INV_X1 U630 ( .A(n608), .ZN(n534) );
  NAND2_X1 U631 ( .A1(G214), .A2(n522), .ZN(n523) );
  XNOR2_X1 U632 ( .A(KEYINPUT91), .B(n523), .ZN(n692) );
  NAND2_X1 U633 ( .A1(G210), .A2(n525), .ZN(n526) );
  XOR2_X1 U634 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n528) );
  NOR2_X1 U635 ( .A1(n692), .A2(n563), .ZN(n532) );
  XNOR2_X1 U636 ( .A(n532), .B(KEYINPUT30), .ZN(n533) );
  INV_X1 U637 ( .A(n539), .ZN(n691) );
  NOR2_X1 U638 ( .A1(n557), .A2(n549), .ZN(n694) );
  NAND2_X1 U639 ( .A1(n698), .A2(n694), .ZN(n540) );
  NOR2_X1 U640 ( .A1(n541), .A2(n675), .ZN(n542) );
  NAND2_X1 U641 ( .A1(n676), .A2(n542), .ZN(n564) );
  NOR2_X1 U642 ( .A1(n379), .A2(n564), .ZN(n543) );
  NAND2_X1 U643 ( .A1(n688), .A2(n556), .ZN(n545) );
  XOR2_X1 U644 ( .A(KEYINPUT42), .B(n545), .Z(n758) );
  AND2_X1 U645 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U646 ( .A1(n557), .A2(n549), .ZN(n593) );
  NOR2_X1 U647 ( .A1(n580), .A2(n593), .ZN(n550) );
  NAND2_X1 U648 ( .A1(n551), .A2(n550), .ZN(n659) );
  XNOR2_X1 U649 ( .A(n659), .B(KEYINPUT81), .ZN(n562) );
  XNOR2_X1 U650 ( .A(KEYINPUT19), .B(KEYINPUT65), .ZN(n554) );
  NAND2_X1 U651 ( .A1(n556), .A2(n588), .ZN(n660) );
  NAND2_X1 U652 ( .A1(n558), .A2(n557), .ZN(n656) );
  INV_X1 U653 ( .A(n656), .ZN(n665) );
  NOR2_X1 U654 ( .A1(n663), .A2(n665), .ZN(n696) );
  NOR2_X1 U655 ( .A1(KEYINPUT47), .A2(n696), .ZN(n559) );
  XOR2_X1 U656 ( .A(KEYINPUT74), .B(n559), .Z(n560) );
  NOR2_X1 U657 ( .A1(n660), .A2(n560), .ZN(n561) );
  INV_X1 U658 ( .A(n663), .ZN(n661) );
  XOR2_X1 U659 ( .A(KEYINPUT114), .B(n565), .Z(n566) );
  XNOR2_X2 U660 ( .A(n567), .B(KEYINPUT1), .ZN(n679) );
  NAND2_X1 U661 ( .A1(n569), .A2(n598), .ZN(n669) );
  NAND2_X1 U662 ( .A1(n570), .A2(n669), .ZN(n574) );
  NAND2_X1 U663 ( .A1(n660), .A2(KEYINPUT47), .ZN(n571) );
  XNOR2_X1 U664 ( .A(n571), .B(KEYINPUT80), .ZN(n573) );
  NAND2_X1 U665 ( .A1(n696), .A2(KEYINPUT47), .ZN(n572) );
  AND2_X1 U666 ( .A1(n577), .A2(n665), .ZN(n670) );
  INV_X1 U667 ( .A(n670), .ZN(n582) );
  OR2_X1 U668 ( .A1(n578), .A2(n679), .ZN(n579) );
  XNOR2_X1 U669 ( .A(n579), .B(KEYINPUT43), .ZN(n581) );
  NAND2_X1 U670 ( .A1(n581), .A2(n580), .ZN(n671) );
  NAND2_X1 U671 ( .A1(n680), .A2(n679), .ZN(n612) );
  INV_X1 U672 ( .A(n583), .ZN(n586) );
  NOR2_X1 U673 ( .A1(G898), .A2(n748), .ZN(n733) );
  NAND2_X1 U674 ( .A1(n733), .A2(n584), .ZN(n585) );
  NAND2_X1 U675 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U676 ( .A(KEYINPUT93), .B(n587), .Z(n589) );
  NOR2_X1 U677 ( .A1(n672), .A2(n609), .ZN(n592) );
  INV_X1 U678 ( .A(KEYINPUT72), .ZN(n591) );
  NOR2_X1 U679 ( .A1(KEYINPUT44), .A2(n759), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n694), .A2(n676), .ZN(n594) );
  XNOR2_X1 U681 ( .A(n594), .B(KEYINPUT111), .ZN(n595) );
  XOR2_X1 U682 ( .A(KEYINPUT22), .B(KEYINPUT64), .Z(n596) );
  XNOR2_X1 U683 ( .A(KEYINPUT73), .B(n596), .ZN(n597) );
  INV_X1 U684 ( .A(n675), .ZN(n620) );
  NOR2_X2 U685 ( .A1(n679), .A2(n601), .ZN(n619) );
  NAND2_X1 U686 ( .A1(n620), .A2(n619), .ZN(n602) );
  NOR2_X1 U687 ( .A1(n757), .A2(n655), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n603), .A2(n605), .ZN(n607) );
  AND2_X1 U689 ( .A1(KEYINPUT86), .A2(KEYINPUT44), .ZN(n604) );
  INV_X1 U690 ( .A(KEYINPUT44), .ZN(n606) );
  NOR2_X1 U691 ( .A1(n379), .A2(n612), .ZN(n685) );
  NAND2_X1 U692 ( .A1(n613), .A2(n685), .ZN(n614) );
  XNOR2_X1 U693 ( .A(n614), .B(KEYINPUT102), .ZN(n615) );
  XNOR2_X1 U694 ( .A(KEYINPUT31), .B(n615), .ZN(n666) );
  NOR2_X1 U695 ( .A1(n696), .A2(n616), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n621), .B(KEYINPUT112), .ZN(n760) );
  INV_X1 U697 ( .A(n760), .ZN(n622) );
  INV_X1 U698 ( .A(KEYINPUT45), .ZN(n623) );
  XNOR2_X2 U699 ( .A(n624), .B(n623), .ZN(n712) );
  INV_X1 U700 ( .A(KEYINPUT83), .ZN(n625) );
  XNOR2_X1 U701 ( .A(n627), .B(n626), .ZN(n630) );
  INV_X1 U702 ( .A(KEYINPUT2), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n709), .B(n628), .ZN(n629) );
  AND2_X2 U704 ( .A1(n630), .A2(n629), .ZN(n720) );
  NAND2_X1 U705 ( .A1(n728), .A2(G469), .ZN(n635) );
  XOR2_X1 U706 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n633) );
  XNOR2_X1 U707 ( .A(n631), .B(KEYINPUT123), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n633), .B(n632), .ZN(n634) );
  XOR2_X1 U709 ( .A(KEYINPUT87), .B(KEYINPUT55), .Z(n639) );
  XNOR2_X1 U710 ( .A(n637), .B(KEYINPUT54), .ZN(n638) );
  NAND2_X1 U711 ( .A1(n720), .A2(G210), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n641), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U713 ( .A1(n720), .A2(G472), .ZN(n645) );
  XOR2_X1 U714 ( .A(KEYINPUT62), .B(KEYINPUT117), .Z(n642) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(n646) );
  INV_X1 U717 ( .A(KEYINPUT90), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n650), .A2(n663), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n649), .B(G104), .ZN(G6) );
  XNOR2_X1 U720 ( .A(G107), .B(KEYINPUT27), .ZN(n654) );
  XOR2_X1 U721 ( .A(KEYINPUT118), .B(KEYINPUT26), .Z(n652) );
  NAND2_X1 U722 ( .A1(n650), .A2(n665), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U724 ( .A(n654), .B(n653), .ZN(G9) );
  XOR2_X1 U725 ( .A(G110), .B(n655), .Z(G12) );
  NOR2_X1 U726 ( .A1(n660), .A2(n656), .ZN(n658) );
  XNOR2_X1 U727 ( .A(G128), .B(KEYINPUT29), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n658), .B(n657), .ZN(G30) );
  XNOR2_X1 U729 ( .A(G143), .B(n659), .ZN(G45) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U731 ( .A(n372), .B(n662), .Z(G48) );
  NAND2_X1 U732 ( .A1(n666), .A2(n663), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n664), .B(G113), .ZN(G15) );
  NAND2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n667), .B(G116), .ZN(G18) );
  XOR2_X1 U736 ( .A(G125), .B(KEYINPUT37), .Z(n668) );
  XNOR2_X1 U737 ( .A(n669), .B(n668), .ZN(G27) );
  XOR2_X1 U738 ( .A(G134), .B(n670), .Z(G36) );
  XNOR2_X1 U739 ( .A(G140), .B(n671), .ZN(G42) );
  INV_X1 U740 ( .A(n688), .ZN(n673) );
  NOR2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U742 ( .A1(G953), .A2(n674), .ZN(n718) );
  NOR2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U744 ( .A(n677), .B(KEYINPUT49), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n379), .A2(n678), .ZN(n683) );
  NOR2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n681), .B(KEYINPUT50), .ZN(n682) );
  NOR2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U750 ( .A(KEYINPUT119), .B(n686), .Z(n687) );
  XNOR2_X1 U751 ( .A(KEYINPUT51), .B(n687), .ZN(n689) );
  NAND2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U753 ( .A(KEYINPUT120), .B(n690), .Z(n704) );
  NAND2_X1 U754 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U755 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U756 ( .A(KEYINPUT121), .B(n695), .ZN(n701) );
  INV_X1 U757 ( .A(n696), .ZN(n697) );
  NAND2_X1 U758 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U759 ( .A(KEYINPUT122), .B(n699), .Z(n700) );
  NOR2_X1 U760 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U761 ( .A1(n702), .A2(n672), .ZN(n703) );
  NOR2_X1 U762 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U763 ( .A(n705), .B(KEYINPUT52), .ZN(n706) );
  NOR2_X1 U764 ( .A1(n707), .A2(n706), .ZN(n716) );
  NAND2_X1 U765 ( .A1(n628), .A2(n747), .ZN(n708) );
  XNOR2_X1 U766 ( .A(n708), .B(KEYINPUT82), .ZN(n711) );
  NAND2_X1 U767 ( .A1(KEYINPUT2), .A2(n709), .ZN(n710) );
  NAND2_X1 U768 ( .A1(n711), .A2(n710), .ZN(n714) );
  INV_X1 U769 ( .A(n712), .ZN(n739) );
  NOR2_X1 U770 ( .A1(n739), .A2(KEYINPUT2), .ZN(n713) );
  NOR2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U772 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U773 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U774 ( .A(KEYINPUT53), .B(n719), .Z(G75) );
  NAND2_X1 U775 ( .A1(n720), .A2(G475), .ZN(n723) );
  XOR2_X1 U776 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n721) );
  XNOR2_X1 U777 ( .A(n723), .B(n363), .ZN(n724) );
  NAND2_X1 U778 ( .A1(G478), .A2(n728), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n732), .A2(n727), .ZN(G63) );
  NAND2_X1 U781 ( .A1(G217), .A2(n728), .ZN(n729) );
  XNOR2_X1 U782 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n732), .A2(n731), .ZN(G66) );
  NOR2_X1 U784 ( .A1(n734), .A2(n733), .ZN(n743) );
  XOR2_X1 U785 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n736) );
  NAND2_X1 U786 ( .A1(G224), .A2(G953), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U788 ( .A(KEYINPUT125), .B(n737), .ZN(n738) );
  NAND2_X1 U789 ( .A1(n738), .A2(G898), .ZN(n741) );
  NAND2_X1 U790 ( .A1(n739), .A2(n748), .ZN(n740) );
  NAND2_X1 U791 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n743), .B(n742), .ZN(G69) );
  XOR2_X1 U793 ( .A(n744), .B(KEYINPUT94), .Z(n745) );
  XNOR2_X1 U794 ( .A(n746), .B(n745), .ZN(n750) );
  XNOR2_X1 U795 ( .A(n747), .B(n750), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(n755) );
  XNOR2_X1 U797 ( .A(G227), .B(n750), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n751), .A2(G900), .ZN(n752) );
  XOR2_X1 U799 ( .A(KEYINPUT127), .B(n752), .Z(n753) );
  NAND2_X1 U800 ( .A1(G953), .A2(n753), .ZN(n754) );
  NAND2_X1 U801 ( .A1(n755), .A2(n754), .ZN(G72) );
  XOR2_X1 U802 ( .A(G131), .B(n756), .Z(G33) );
  XOR2_X1 U803 ( .A(G119), .B(n757), .Z(G21) );
  XOR2_X1 U804 ( .A(G137), .B(n758), .Z(G39) );
  XOR2_X1 U805 ( .A(n759), .B(G122), .Z(G24) );
  XOR2_X1 U806 ( .A(n760), .B(G101), .Z(G3) );
endmodule

