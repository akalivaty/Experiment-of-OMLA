

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770;

  AND2_X2 U376 ( .A1(n369), .A2(n360), .ZN(n724) );
  XNOR2_X1 U377 ( .A(n382), .B(G119), .ZN(n466) );
  XNOR2_X1 U378 ( .A(n742), .B(n518), .ZN(n725) );
  XNOR2_X2 U379 ( .A(n517), .B(n516), .ZN(n742) );
  XNOR2_X2 U380 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n642) );
  XOR2_X2 U381 ( .A(KEYINPUT66), .B(KEYINPUT22), .Z(n363) );
  NOR2_X2 U382 ( .A1(n716), .A2(n732), .ZN(n718) );
  NOR2_X2 U383 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U384 ( .A1(n607), .A2(n666), .ZN(n663) );
  XNOR2_X1 U385 ( .A(n402), .B(n401), .ZN(n518) );
  NAND2_X1 U386 ( .A1(n357), .A2(n356), .ZN(n354) );
  AND2_X2 U387 ( .A1(n411), .A2(n354), .ZN(n410) );
  NOR2_X2 U388 ( .A1(n652), .A2(n732), .ZN(n654) );
  INV_X2 U389 ( .A(G146), .ZN(n376) );
  NAND2_X1 U390 ( .A1(n385), .A2(n383), .ZN(n704) );
  AND2_X1 U391 ( .A1(n390), .A2(n386), .ZN(n385) );
  XNOR2_X1 U392 ( .A(n403), .B(KEYINPUT82), .ZN(n392) );
  NAND2_X1 U393 ( .A1(n404), .A2(n360), .ZN(n403) );
  NAND2_X1 U394 ( .A1(n366), .A2(n408), .ZN(n407) );
  NOR2_X1 U395 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U396 ( .A(n455), .B(G104), .ZN(n515) );
  XNOR2_X1 U397 ( .A(n579), .B(KEYINPUT19), .ZN(n574) );
  NAND2_X1 U398 ( .A1(n410), .A2(n407), .ZN(n579) );
  OR2_X1 U399 ( .A1(n725), .A2(n406), .ZN(n355) );
  OR2_X1 U400 ( .A1(n725), .A2(n406), .ZN(n413) );
  XNOR2_X1 U401 ( .A(n378), .B(n377), .ZN(n622) );
  NOR2_X2 U402 ( .A1(n698), .A2(n618), .ZN(n619) );
  XNOR2_X2 U403 ( .A(n617), .B(n616), .ZN(n698) );
  NOR2_X1 U404 ( .A1(n522), .A2(n525), .ZN(n356) );
  XNOR2_X1 U405 ( .A(n518), .B(n742), .ZN(n357) );
  BUF_X1 U406 ( .A(n658), .Z(n746) );
  NAND2_X1 U407 ( .A1(n622), .A2(n358), .ZN(n639) );
  INV_X1 U408 ( .A(KEYINPUT70), .ZN(n464) );
  INV_X1 U409 ( .A(KEYINPUT121), .ZN(n388) );
  NAND2_X1 U410 ( .A1(G234), .A2(G237), .ZN(n420) );
  NOR2_X1 U411 ( .A1(n770), .A2(n766), .ZN(n375) );
  INV_X1 U412 ( .A(KEYINPUT88), .ZN(n380) );
  OR2_X1 U413 ( .A1(n521), .A2(n520), .ZN(n381) );
  NOR2_X1 U414 ( .A1(n409), .A2(KEYINPUT85), .ZN(n408) );
  XNOR2_X1 U415 ( .A(n643), .B(n642), .ZN(n658) );
  XNOR2_X1 U416 ( .A(n452), .B(G131), .ZN(n453) );
  XNOR2_X1 U417 ( .A(KEYINPUT4), .B(G137), .ZN(n452) );
  XNOR2_X1 U418 ( .A(n515), .B(n514), .ZN(n517) );
  AND2_X1 U419 ( .A1(n644), .A2(KEYINPUT65), .ZN(n400) );
  NAND2_X1 U420 ( .A1(n397), .A2(n395), .ZN(n394) );
  NAND2_X1 U421 ( .A1(n646), .A2(n396), .ZN(n395) );
  NAND2_X1 U422 ( .A1(n414), .A2(n398), .ZN(n397) );
  NAND2_X1 U423 ( .A1(KEYINPUT2), .A2(n398), .ZN(n396) );
  AND2_X1 U424 ( .A1(n387), .A2(n762), .ZN(n386) );
  NAND2_X1 U425 ( .A1(n389), .A2(n388), .ZN(n387) );
  NOR2_X1 U426 ( .A1(G953), .A2(G237), .ZN(n492) );
  XNOR2_X1 U427 ( .A(G902), .B(KEYINPUT87), .ZN(n439) );
  NOR2_X1 U428 ( .A1(G237), .A2(G902), .ZN(n475) );
  XNOR2_X1 U429 ( .A(n425), .B(KEYINPUT91), .ZN(n526) );
  XNOR2_X1 U430 ( .A(G143), .B(G104), .ZN(n497) );
  INV_X1 U431 ( .A(KEYINPUT65), .ZN(n398) );
  AND2_X1 U432 ( .A1(n609), .A2(n545), .ZN(n615) );
  NAND2_X1 U433 ( .A1(n417), .A2(n646), .ZN(n415) );
  INV_X1 U434 ( .A(G902), .ZN(n503) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n605) );
  INV_X1 U436 ( .A(KEYINPUT48), .ZN(n372) );
  XNOR2_X1 U437 ( .A(G140), .B(KEYINPUT10), .ZN(n429) );
  INV_X1 U438 ( .A(G134), .ZN(n449) );
  INV_X1 U439 ( .A(n702), .ZN(n389) );
  BUF_X1 U440 ( .A(G107), .Z(n539) );
  NAND2_X1 U441 ( .A1(n371), .A2(n370), .ZN(n369) );
  AND2_X1 U442 ( .A1(n399), .A2(n394), .ZN(n371) );
  BUF_X1 U443 ( .A(n515), .Z(n458) );
  NOR2_X1 U444 ( .A1(n762), .A2(G952), .ZN(n732) );
  XNOR2_X1 U445 ( .A(n597), .B(n418), .ZN(n770) );
  INV_X1 U446 ( .A(KEYINPUT35), .ZN(n377) );
  XNOR2_X1 U447 ( .A(n612), .B(KEYINPUT32), .ZN(n657) );
  NAND2_X1 U448 ( .A1(n384), .A2(n388), .ZN(n383) );
  AND2_X1 U449 ( .A1(n657), .A2(n613), .ZN(n358) );
  AND2_X1 U450 ( .A1(n415), .A2(n680), .ZN(n359) );
  OR2_X1 U451 ( .A1(n647), .A2(n648), .ZN(n360) );
  XNOR2_X1 U452 ( .A(n381), .B(n380), .ZN(n522) );
  AND2_X1 U453 ( .A1(n355), .A2(n415), .ZN(n361) );
  AND2_X1 U454 ( .A1(n611), .A2(n623), .ZN(n362) );
  INV_X1 U455 ( .A(KEYINPUT85), .ZN(n525) );
  INV_X1 U456 ( .A(n646), .ZN(n414) );
  AND2_X1 U457 ( .A1(n646), .A2(n398), .ZN(n364) );
  XOR2_X1 U458 ( .A(G143), .B(G128), .Z(n365) );
  BUF_X1 U459 ( .A(n742), .Z(n743) );
  AND2_X1 U460 ( .A1(n355), .A2(n359), .ZN(n366) );
  NAND2_X1 U461 ( .A1(n367), .A2(n624), .ZN(n625) );
  NAND2_X1 U462 ( .A1(n367), .A2(n362), .ZN(n612) );
  AND2_X1 U463 ( .A1(n367), .A2(n664), .ZN(n557) );
  XNOR2_X2 U464 ( .A(n555), .B(n363), .ZN(n367) );
  NAND2_X1 U465 ( .A1(n368), .A2(n738), .ZN(n597) );
  NAND2_X1 U466 ( .A1(n368), .A2(n735), .ZN(n741) );
  XNOR2_X2 U467 ( .A(n596), .B(KEYINPUT39), .ZN(n368) );
  NAND2_X1 U468 ( .A1(n393), .A2(n364), .ZN(n370) );
  NAND2_X1 U469 ( .A1(n602), .A2(n374), .ZN(n373) );
  XNOR2_X1 U470 ( .A(n375), .B(KEYINPUT46), .ZN(n374) );
  XNOR2_X2 U471 ( .A(n507), .B(n429), .ZN(n756) );
  XNOR2_X2 U472 ( .A(n376), .B(G125), .ZN(n507) );
  INV_X1 U473 ( .A(n622), .ZN(n705) );
  NAND2_X1 U474 ( .A1(n379), .A2(n621), .ZN(n378) );
  XNOR2_X1 U475 ( .A(n619), .B(KEYINPUT34), .ZN(n379) );
  XNOR2_X1 U476 ( .A(n405), .B(KEYINPUT79), .ZN(n404) );
  XNOR2_X2 U477 ( .A(n755), .B(n454), .ZN(n471) );
  OR2_X2 U478 ( .A1(n628), .A2(n627), .ZN(n631) );
  NOR2_X2 U479 ( .A1(n618), .A2(n673), .ZN(n546) );
  NAND2_X1 U480 ( .A1(n639), .A2(KEYINPUT44), .ZN(n636) );
  XNOR2_X2 U481 ( .A(G116), .B(KEYINPUT3), .ZN(n382) );
  INV_X1 U482 ( .A(n392), .ZN(n384) );
  NAND2_X1 U483 ( .A1(n392), .A2(n391), .ZN(n390) );
  AND2_X1 U484 ( .A1(n702), .A2(KEYINPUT121), .ZN(n391) );
  XNOR2_X1 U485 ( .A(n510), .B(n511), .ZN(n512) );
  XNOR2_X2 U486 ( .A(G101), .B(KEYINPUT67), .ZN(n511) );
  XNOR2_X2 U487 ( .A(G143), .B(G128), .ZN(n510) );
  INV_X1 U488 ( .A(n645), .ZN(n393) );
  NAND2_X1 U489 ( .A1(n645), .A2(n400), .ZN(n399) );
  NAND2_X1 U490 ( .A1(n522), .A2(n414), .ZN(n406) );
  NOR2_X2 U491 ( .A1(n573), .A2(n572), .ZN(n599) );
  NOR2_X2 U492 ( .A1(n561), .A2(n560), .ZN(n568) );
  XNOR2_X2 U493 ( .A(n577), .B(KEYINPUT77), .ZN(n739) );
  XNOR2_X1 U494 ( .A(n507), .B(n506), .ZN(n401) );
  XNOR2_X1 U495 ( .A(n512), .B(n509), .ZN(n402) );
  NAND2_X1 U496 ( .A1(n662), .A2(n661), .ZN(n405) );
  INV_X1 U497 ( .A(n416), .ZN(n409) );
  NAND2_X1 U498 ( .A1(n412), .A2(KEYINPUT85), .ZN(n411) );
  NAND2_X1 U499 ( .A1(n361), .A2(n416), .ZN(n524) );
  NAND2_X1 U500 ( .A1(n413), .A2(n359), .ZN(n412) );
  NAND2_X1 U501 ( .A1(n357), .A2(n417), .ZN(n416) );
  INV_X1 U502 ( .A(n522), .ZN(n417) );
  XNOR2_X1 U503 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n418) );
  XOR2_X1 U504 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n419) );
  XOR2_X1 U505 ( .A(KEYINPUT89), .B(KEYINPUT14), .Z(n421) );
  XNOR2_X1 U506 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U507 ( .A(KEYINPUT73), .B(n422), .Z(n424) );
  NAND2_X1 U508 ( .A1(G952), .A2(n424), .ZN(n423) );
  XNOR2_X1 U509 ( .A(n423), .B(KEYINPUT90), .ZN(n694) );
  NOR2_X1 U510 ( .A1(n694), .A2(G953), .ZN(n530) );
  NAND2_X1 U511 ( .A1(G902), .A2(n424), .ZN(n425) );
  NAND2_X1 U512 ( .A1(G953), .A2(n526), .ZN(n426) );
  NOR2_X1 U513 ( .A1(G900), .A2(n426), .ZN(n427) );
  NOR2_X1 U514 ( .A1(n530), .A2(n427), .ZN(n428) );
  XNOR2_X1 U515 ( .A(KEYINPUT78), .B(n428), .ZN(n561) );
  XOR2_X1 U516 ( .A(G110), .B(G137), .Z(n431) );
  XNOR2_X1 U517 ( .A(G119), .B(G128), .ZN(n430) );
  XNOR2_X1 U518 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U519 ( .A(n756), .B(n432), .ZN(n437) );
  INV_X4 U520 ( .A(G953), .ZN(n762) );
  NAND2_X1 U521 ( .A1(G234), .A2(n762), .ZN(n433) );
  XOR2_X1 U522 ( .A(KEYINPUT8), .B(n433), .Z(n480) );
  NAND2_X1 U523 ( .A1(G221), .A2(n480), .ZN(n435) );
  XOR2_X1 U524 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n434) );
  XNOR2_X1 U525 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U526 ( .A(n437), .B(n436), .ZN(n707) );
  NAND2_X1 U527 ( .A1(n707), .A2(n503), .ZN(n445) );
  XOR2_X1 U528 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n441) );
  INV_X1 U529 ( .A(KEYINPUT15), .ZN(n438) );
  XNOR2_X1 U530 ( .A(n439), .B(n438), .ZN(n519) );
  NAND2_X1 U531 ( .A1(G234), .A2(n519), .ZN(n440) );
  XNOR2_X1 U532 ( .A(n441), .B(n440), .ZN(n446) );
  NAND2_X1 U533 ( .A1(n446), .A2(G217), .ZN(n443) );
  INV_X1 U534 ( .A(KEYINPUT25), .ZN(n442) );
  XNOR2_X1 U535 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X2 U536 ( .A(n445), .B(n444), .ZN(n607) );
  NAND2_X1 U537 ( .A1(G221), .A2(n446), .ZN(n448) );
  XOR2_X1 U538 ( .A(KEYINPUT21), .B(KEYINPUT94), .Z(n447) );
  XNOR2_X1 U539 ( .A(n448), .B(n447), .ZN(n666) );
  INV_X1 U540 ( .A(n663), .ZN(n545) );
  NAND2_X1 U541 ( .A1(n510), .A2(G134), .ZN(n451) );
  NAND2_X1 U542 ( .A1(n365), .A2(n449), .ZN(n450) );
  NAND2_X1 U543 ( .A1(n451), .A2(n450), .ZN(n481) );
  XNOR2_X2 U544 ( .A(n481), .B(n453), .ZN(n755) );
  XNOR2_X1 U545 ( .A(n376), .B(n511), .ZN(n454) );
  XNOR2_X2 U546 ( .A(G110), .B(G107), .ZN(n455) );
  NAND2_X1 U547 ( .A1(G227), .A2(n762), .ZN(n456) );
  XNOR2_X1 U548 ( .A(n456), .B(G140), .ZN(n457) );
  XNOR2_X1 U549 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U550 ( .A(n471), .B(n459), .ZN(n720) );
  NAND2_X1 U551 ( .A1(n720), .A2(n503), .ZN(n461) );
  XOR2_X1 U552 ( .A(KEYINPUT69), .B(G469), .Z(n460) );
  XNOR2_X2 U553 ( .A(n461), .B(n460), .ZN(n571) );
  AND2_X2 U554 ( .A1(n545), .A2(n571), .ZN(n533) );
  XNOR2_X1 U555 ( .A(n533), .B(KEYINPUT105), .ZN(n462) );
  NOR2_X1 U556 ( .A1(n561), .A2(n462), .ZN(n463) );
  XNOR2_X1 U557 ( .A(KEYINPUT76), .B(n463), .ZN(n479) );
  XNOR2_X1 U558 ( .A(n464), .B(G113), .ZN(n465) );
  XNOR2_X2 U559 ( .A(n466), .B(n465), .ZN(n516) );
  XOR2_X1 U560 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n468) );
  NAND2_X1 U561 ( .A1(n492), .A2(G210), .ZN(n467) );
  XNOR2_X1 U562 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U563 ( .A(n516), .B(n469), .ZN(n470) );
  XNOR2_X1 U564 ( .A(n471), .B(n470), .ZN(n649) );
  NAND2_X1 U565 ( .A1(n649), .A2(n503), .ZN(n474) );
  INV_X1 U566 ( .A(KEYINPUT95), .ZN(n472) );
  XNOR2_X1 U567 ( .A(n472), .B(G472), .ZN(n473) );
  XNOR2_X2 U568 ( .A(n474), .B(n473), .ZN(n670) );
  XNOR2_X1 U569 ( .A(n475), .B(KEYINPUT74), .ZN(n521) );
  INV_X1 U570 ( .A(G214), .ZN(n476) );
  OR2_X1 U571 ( .A1(n521), .A2(n476), .ZN(n680) );
  NAND2_X1 U572 ( .A1(n670), .A2(n680), .ZN(n477) );
  XOR2_X1 U573 ( .A(KEYINPUT30), .B(n477), .Z(n478) );
  AND2_X2 U574 ( .A1(n479), .A2(n478), .ZN(n595) );
  NAND2_X1 U575 ( .A1(n480), .A2(G217), .ZN(n482) );
  XNOR2_X1 U576 ( .A(n482), .B(n481), .ZN(n489) );
  XOR2_X1 U577 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n484) );
  XNOR2_X1 U578 ( .A(n539), .B(KEYINPUT100), .ZN(n483) );
  XNOR2_X1 U579 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U580 ( .A(n485), .B(KEYINPUT99), .Z(n487) );
  XNOR2_X1 U581 ( .A(G116), .B(G122), .ZN(n486) );
  XNOR2_X1 U582 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U583 ( .A(n489), .B(n488), .ZN(n710) );
  NAND2_X1 U584 ( .A1(n710), .A2(n503), .ZN(n491) );
  INV_X1 U585 ( .A(G478), .ZN(n490) );
  XNOR2_X1 U586 ( .A(n491), .B(n490), .ZN(n551) );
  INV_X1 U587 ( .A(n551), .ZN(n538) );
  XOR2_X1 U588 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n494) );
  NAND2_X1 U589 ( .A1(G214), .A2(n492), .ZN(n493) );
  XNOR2_X1 U590 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U591 ( .A(n495), .B(KEYINPUT12), .Z(n496) );
  XNOR2_X1 U592 ( .A(n756), .B(n496), .ZN(n502) );
  XOR2_X1 U593 ( .A(KEYINPUT97), .B(G122), .Z(n498) );
  XNOR2_X1 U594 ( .A(n498), .B(n497), .ZN(n500) );
  XOR2_X1 U595 ( .A(G113), .B(G131), .Z(n499) );
  XNOR2_X1 U596 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U597 ( .A(n502), .B(n501), .ZN(n713) );
  NAND2_X1 U598 ( .A1(n713), .A2(n503), .ZN(n505) );
  XNOR2_X1 U599 ( .A(KEYINPUT13), .B(G475), .ZN(n504) );
  XNOR2_X1 U600 ( .A(n505), .B(n504), .ZN(n550) );
  INV_X1 U601 ( .A(n550), .ZN(n536) );
  NAND2_X1 U602 ( .A1(n538), .A2(n536), .ZN(n620) );
  XNOR2_X1 U603 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n506) );
  NAND2_X1 U604 ( .A1(n762), .A2(G224), .ZN(n508) );
  XNOR2_X1 U605 ( .A(n508), .B(KEYINPUT4), .ZN(n509) );
  XNOR2_X1 U606 ( .A(KEYINPUT71), .B(KEYINPUT16), .ZN(n513) );
  XNOR2_X1 U607 ( .A(n513), .B(G122), .ZN(n514) );
  INV_X1 U608 ( .A(n519), .ZN(n646) );
  INV_X1 U609 ( .A(G210), .ZN(n520) );
  NOR2_X1 U610 ( .A1(n620), .A2(n524), .ZN(n523) );
  NAND2_X1 U611 ( .A1(n595), .A2(n523), .ZN(n585) );
  XNOR2_X1 U612 ( .A(n585), .B(G143), .ZN(G45) );
  NOR2_X1 U613 ( .A1(G898), .A2(n762), .ZN(n744) );
  NAND2_X1 U614 ( .A1(n526), .A2(n744), .ZN(n528) );
  INV_X1 U615 ( .A(KEYINPUT92), .ZN(n527) );
  XNOR2_X1 U616 ( .A(n528), .B(n527), .ZN(n529) );
  NOR2_X2 U617 ( .A1(n574), .A2(n531), .ZN(n532) );
  XNOR2_X2 U618 ( .A(n532), .B(KEYINPUT0), .ZN(n554) );
  INV_X1 U619 ( .A(n670), .ZN(n534) );
  AND2_X1 U620 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U621 ( .A1(n554), .A2(n535), .ZN(n627) );
  NAND2_X1 U622 ( .A1(n536), .A2(n551), .ZN(n563) );
  INV_X1 U623 ( .A(n563), .ZN(n738) );
  NAND2_X1 U624 ( .A1(n627), .A2(n738), .ZN(n537) );
  XNOR2_X1 U625 ( .A(n537), .B(G104), .ZN(G6) );
  AND2_X1 U626 ( .A1(n538), .A2(n550), .ZN(n735) );
  NAND2_X1 U627 ( .A1(n627), .A2(n735), .ZN(n544) );
  XOR2_X1 U628 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n541) );
  XNOR2_X1 U629 ( .A(n539), .B(KEYINPUT26), .ZN(n540) );
  XNOR2_X1 U630 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U631 ( .A(KEYINPUT111), .B(n542), .Z(n543) );
  XNOR2_X1 U632 ( .A(n544), .B(n543), .ZN(G9) );
  INV_X1 U633 ( .A(n554), .ZN(n618) );
  XNOR2_X2 U634 ( .A(n571), .B(KEYINPUT1), .ZN(n609) );
  NAND2_X1 U635 ( .A1(n615), .A2(n670), .ZN(n673) );
  XNOR2_X2 U636 ( .A(n546), .B(n419), .ZN(n628) );
  NAND2_X1 U637 ( .A1(n628), .A2(n735), .ZN(n548) );
  XOR2_X1 U638 ( .A(G116), .B(KEYINPUT113), .Z(n547) );
  XNOR2_X1 U639 ( .A(n548), .B(n547), .ZN(G18) );
  NAND2_X1 U640 ( .A1(n628), .A2(n738), .ZN(n549) );
  XNOR2_X1 U641 ( .A(n549), .B(G113), .ZN(G15) );
  NAND2_X1 U642 ( .A1(n551), .A2(n550), .ZN(n684) );
  INV_X1 U643 ( .A(n666), .ZN(n552) );
  NOR2_X1 U644 ( .A1(n684), .A2(n552), .ZN(n553) );
  NAND2_X1 U645 ( .A1(n553), .A2(n554), .ZN(n555) );
  NOR2_X1 U646 ( .A1(n670), .A2(n607), .ZN(n556) );
  NAND2_X1 U647 ( .A1(n557), .A2(n556), .ZN(n613) );
  XNOR2_X1 U648 ( .A(n613), .B(G110), .ZN(G12) );
  INV_X1 U649 ( .A(KEYINPUT6), .ZN(n558) );
  XNOR2_X1 U650 ( .A(n670), .B(n558), .ZN(n614) );
  INV_X1 U651 ( .A(n607), .ZN(n559) );
  NAND2_X1 U652 ( .A1(n666), .A2(n559), .ZN(n560) );
  NAND2_X1 U653 ( .A1(n614), .A2(n568), .ZN(n562) );
  NOR2_X1 U654 ( .A1(n563), .A2(n562), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n581), .A2(n680), .ZN(n564) );
  NOR2_X1 U656 ( .A1(n609), .A2(n564), .ZN(n566) );
  XNOR2_X1 U657 ( .A(KEYINPUT43), .B(KEYINPUT104), .ZN(n565) );
  XOR2_X1 U658 ( .A(n566), .B(n565), .Z(n567) );
  NAND2_X1 U659 ( .A1(n567), .A2(n524), .ZN(n603) );
  XNOR2_X1 U660 ( .A(n603), .B(G140), .ZN(G42) );
  OR2_X1 U661 ( .A1(n738), .A2(n735), .ZN(n587) );
  INV_X1 U662 ( .A(n587), .ZN(n686) );
  XOR2_X1 U663 ( .A(KEYINPUT28), .B(KEYINPUT106), .Z(n570) );
  NAND2_X1 U664 ( .A1(n670), .A2(n568), .ZN(n569) );
  XOR2_X1 U665 ( .A(n570), .B(n569), .Z(n573) );
  INV_X1 U666 ( .A(n571), .ZN(n572) );
  BUF_X1 U667 ( .A(n574), .Z(n575) );
  INV_X1 U668 ( .A(n575), .ZN(n576) );
  NAND2_X1 U669 ( .A1(n599), .A2(n576), .ZN(n577) );
  NAND2_X1 U670 ( .A1(n587), .A2(n739), .ZN(n578) );
  NAND2_X1 U671 ( .A1(n578), .A2(KEYINPUT47), .ZN(n594) );
  INV_X1 U672 ( .A(n609), .ZN(n664) );
  BUF_X1 U673 ( .A(n579), .Z(n580) );
  NAND2_X1 U674 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U675 ( .A(n582), .B(KEYINPUT36), .ZN(n583) );
  NOR2_X1 U676 ( .A1(n664), .A2(n583), .ZN(n584) );
  XNOR2_X1 U677 ( .A(KEYINPUT109), .B(n584), .ZN(n768) );
  NAND2_X1 U678 ( .A1(n768), .A2(n585), .ZN(n592) );
  INV_X1 U679 ( .A(KEYINPUT80), .ZN(n586) );
  XNOR2_X1 U680 ( .A(n587), .B(n586), .ZN(n629) );
  XNOR2_X1 U681 ( .A(KEYINPUT68), .B(KEYINPUT47), .ZN(n588) );
  NOR2_X1 U682 ( .A1(n629), .A2(n588), .ZN(n589) );
  NAND2_X1 U683 ( .A1(n739), .A2(n589), .ZN(n590) );
  XOR2_X1 U684 ( .A(KEYINPUT72), .B(n590), .Z(n591) );
  NOR2_X1 U685 ( .A1(n592), .A2(n591), .ZN(n593) );
  AND2_X1 U686 ( .A1(n594), .A2(n593), .ZN(n602) );
  XNOR2_X1 U687 ( .A(n524), .B(KEYINPUT38), .ZN(n681) );
  NAND2_X1 U688 ( .A1(n595), .A2(n681), .ZN(n596) );
  XOR2_X1 U689 ( .A(KEYINPUT42), .B(KEYINPUT108), .Z(n601) );
  NAND2_X1 U690 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U691 ( .A1(n685), .A2(n684), .ZN(n598) );
  XOR2_X1 U692 ( .A(KEYINPUT41), .B(n598), .Z(n677) );
  NAND2_X1 U693 ( .A1(n599), .A2(n677), .ZN(n600) );
  XNOR2_X1 U694 ( .A(n601), .B(n600), .ZN(n766) );
  AND2_X1 U695 ( .A1(n741), .A2(n603), .ZN(n604) );
  AND2_X2 U696 ( .A1(n605), .A2(n604), .ZN(n759) );
  INV_X1 U697 ( .A(KEYINPUT101), .ZN(n606) );
  XNOR2_X1 U698 ( .A(n607), .B(n606), .ZN(n667) );
  INV_X1 U699 ( .A(n667), .ZN(n608) );
  NAND2_X1 U700 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U701 ( .A(n610), .B(KEYINPUT103), .ZN(n611) );
  INV_X1 U702 ( .A(n614), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n615), .A2(n614), .ZN(n617) );
  INV_X1 U704 ( .A(KEYINPUT33), .ZN(n616) );
  INV_X1 U705 ( .A(n620), .ZN(n621) );
  AND2_X1 U706 ( .A1(n623), .A2(n664), .ZN(n624) );
  XNOR2_X1 U707 ( .A(n625), .B(KEYINPUT83), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n626), .A2(n667), .ZN(n655) );
  INV_X1 U709 ( .A(n629), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n655), .A2(n632), .ZN(n634) );
  INV_X1 U712 ( .A(KEYINPUT102), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n634), .B(n633), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n635), .A2(n636), .ZN(n638) );
  INV_X1 U715 ( .A(KEYINPUT84), .ZN(n637) );
  XNOR2_X1 U716 ( .A(n638), .B(n637), .ZN(n641) );
  OR2_X1 U717 ( .A1(n639), .A2(KEYINPUT44), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n759), .A2(n746), .ZN(n645) );
  INV_X1 U720 ( .A(KEYINPUT2), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n759), .A2(KEYINPUT2), .ZN(n648) );
  INV_X1 U722 ( .A(n746), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n724), .A2(G472), .ZN(n651) );
  XOR2_X1 U724 ( .A(KEYINPUT62), .B(n649), .Z(n650) );
  XNOR2_X1 U725 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U726 ( .A(KEYINPUT110), .B(KEYINPUT63), .Z(n653) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(G57) );
  BUF_X1 U728 ( .A(n655), .Z(n656) );
  XNOR2_X1 U729 ( .A(n656), .B(G101), .ZN(G3) );
  XNOR2_X1 U730 ( .A(n657), .B(G119), .ZN(G21) );
  NOR2_X2 U731 ( .A1(n658), .A2(KEYINPUT2), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(KEYINPUT81), .ZN(n662) );
  NOR2_X1 U733 ( .A1(n759), .A2(KEYINPUT2), .ZN(n660) );
  INV_X1 U734 ( .A(n660), .ZN(n661) );
  NAND2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n665), .B(KEYINPUT50), .ZN(n672) );
  NOR2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U738 ( .A(KEYINPUT49), .B(n668), .Z(n669) );
  NOR2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n676) );
  XOR2_X1 U742 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n675) );
  XNOR2_X1 U743 ( .A(n676), .B(n675), .ZN(n678) );
  INV_X1 U744 ( .A(n677), .ZN(n697) );
  NOR2_X1 U745 ( .A1(n678), .A2(n697), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n679), .B(KEYINPUT116), .ZN(n691) );
  NOR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U748 ( .A(KEYINPUT117), .B(n682), .Z(n683) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U752 ( .A1(n698), .A2(n689), .ZN(n690) );
  NOR2_X1 U753 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U754 ( .A(n692), .B(KEYINPUT118), .ZN(n693) );
  XNOR2_X1 U755 ( .A(KEYINPUT52), .B(n693), .ZN(n695) );
  NOR2_X1 U756 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U757 ( .A(KEYINPUT119), .B(n696), .Z(n701) );
  NOR2_X1 U758 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U759 ( .A(n699), .B(KEYINPUT120), .ZN(n700) );
  NOR2_X1 U760 ( .A1(n701), .A2(n700), .ZN(n702) );
  INV_X1 U761 ( .A(KEYINPUT53), .ZN(n703) );
  XNOR2_X1 U762 ( .A(n704), .B(n703), .ZN(G75) );
  XOR2_X1 U763 ( .A(n705), .B(G122), .Z(G24) );
  NAND2_X1 U764 ( .A1(n724), .A2(G217), .ZN(n706) );
  XOR2_X1 U765 ( .A(n707), .B(n706), .Z(n708) );
  NOR2_X1 U766 ( .A1(n708), .A2(n732), .ZN(G66) );
  NAND2_X1 U767 ( .A1(n724), .A2(G478), .ZN(n709) );
  XOR2_X1 U768 ( .A(n710), .B(n709), .Z(n711) );
  NOR2_X1 U769 ( .A1(n711), .A2(n732), .ZN(G63) );
  NAND2_X1 U770 ( .A1(n724), .A2(G475), .ZN(n715) );
  XOR2_X1 U771 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n712) );
  XNOR2_X1 U772 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U773 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U774 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n717) );
  XNOR2_X1 U775 ( .A(n718), .B(n717), .ZN(G60) );
  NAND2_X1 U776 ( .A1(n724), .A2(G469), .ZN(n722) );
  XNOR2_X1 U777 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n719) );
  XNOR2_X1 U778 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U779 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U780 ( .A1(n723), .A2(n732), .ZN(G54) );
  NAND2_X1 U781 ( .A1(n724), .A2(G210), .ZN(n731) );
  BUF_X1 U782 ( .A(n357), .Z(n729) );
  XOR2_X1 U783 ( .A(KEYINPUT55), .B(KEYINPUT86), .Z(n727) );
  XNOR2_X1 U784 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n726) );
  XNOR2_X1 U785 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U786 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U787 ( .A(n731), .B(n730), .ZN(n733) );
  XNOR2_X1 U788 ( .A(n734), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U789 ( .A(G128), .B(KEYINPUT29), .Z(n737) );
  NAND2_X1 U790 ( .A1(n739), .A2(n735), .ZN(n736) );
  XNOR2_X1 U791 ( .A(n737), .B(n736), .ZN(G30) );
  NAND2_X1 U792 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U793 ( .A(n740), .B(G146), .ZN(G48) );
  XNOR2_X1 U794 ( .A(G134), .B(n741), .ZN(G36) );
  XNOR2_X1 U795 ( .A(n743), .B(G101), .ZN(n745) );
  NOR2_X1 U796 ( .A1(n745), .A2(n744), .ZN(n754) );
  NAND2_X1 U797 ( .A1(n746), .A2(n762), .ZN(n752) );
  XOR2_X1 U798 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n748) );
  NAND2_X1 U799 ( .A1(G224), .A2(G953), .ZN(n747) );
  XNOR2_X1 U800 ( .A(n748), .B(n747), .ZN(n749) );
  NAND2_X1 U801 ( .A1(G898), .A2(n749), .ZN(n750) );
  XNOR2_X1 U802 ( .A(n750), .B(KEYINPUT126), .ZN(n751) );
  NAND2_X1 U803 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U804 ( .A(n754), .B(n753), .ZN(G69) );
  XNOR2_X1 U805 ( .A(n756), .B(n755), .ZN(n760) );
  XNOR2_X1 U806 ( .A(G227), .B(n760), .ZN(n757) );
  NAND2_X1 U807 ( .A1(n757), .A2(G900), .ZN(n758) );
  NAND2_X1 U808 ( .A1(n758), .A2(G953), .ZN(n765) );
  XNOR2_X1 U809 ( .A(n760), .B(n759), .ZN(n761) );
  XNOR2_X1 U810 ( .A(n761), .B(KEYINPUT127), .ZN(n763) );
  NAND2_X1 U811 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U812 ( .A1(n765), .A2(n764), .ZN(G72) );
  XOR2_X1 U813 ( .A(G137), .B(n766), .Z(G39) );
  XOR2_X1 U814 ( .A(KEYINPUT37), .B(KEYINPUT114), .Z(n767) );
  XNOR2_X1 U815 ( .A(n768), .B(n767), .ZN(n769) );
  XNOR2_X1 U816 ( .A(G125), .B(n769), .ZN(G27) );
  XOR2_X1 U817 ( .A(n770), .B(G131), .Z(G33) );
endmodule

