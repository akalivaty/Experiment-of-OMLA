//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n573, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  AND3_X1   g039(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT3), .B1(new_n464), .B2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n463), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n472), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT68), .B1(new_n473), .B2(new_n463), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(G125), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n471), .B1(new_n474), .B2(new_n481), .ZN(G160));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n483), .B1(new_n468), .B2(KEYINPUT69), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n463), .B1(new_n484), .B2(new_n485), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n463), .A2(G112), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n487), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  AND2_X1   g068(.A1(KEYINPUT4), .A2(G138), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n463), .C1(new_n475), .C2(new_n476), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n486), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n484), .B2(new_n485), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G2105), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n510), .A2(G651), .B1(G50), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n507), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT70), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n507), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n515), .B1(new_n516), .B2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(new_n527), .B1(new_n507), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n517), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n512), .A2(KEYINPUT71), .A3(new_n513), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(G543), .A3(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  OAI221_X1 g110(.A(new_n529), .B1(new_n530), .B2(new_n534), .C1(new_n522), .C2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(G168));
  AND3_X1   g112(.A1(new_n532), .A2(G543), .A3(new_n533), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G52), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G651), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n539), .B(new_n542), .C1(new_n543), .C2(new_n522), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT72), .ZN(G171));
  AOI22_X1  g120(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n541), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n522), .A2(new_n548), .B1(new_n549), .B2(new_n534), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n550), .A2(KEYINPUT73), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(KEYINPUT73), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g131(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n557));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n508), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  INV_X1    g139(.A(G91), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n522), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n532), .A2(G53), .A3(G543), .A4(new_n533), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(KEYINPUT75), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n568), .B(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(G299));
  INV_X1    g147(.A(KEYINPUT72), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n544), .B(new_n573), .ZN(G301));
  XNOR2_X1  g149(.A(new_n536), .B(KEYINPUT76), .ZN(G286));
  OAI21_X1  g150(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n576));
  INV_X1    g151(.A(G49), .ZN(new_n577));
  INV_X1    g152(.A(G87), .ZN(new_n578));
  OAI221_X1 g153(.A(new_n576), .B1(new_n577), .B2(new_n534), .C1(new_n522), .C2(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(new_n507), .A2(G61), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G48), .B2(new_n514), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n519), .A2(G86), .A3(new_n521), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT77), .ZN(G305));
  AND2_X1   g161(.A1(new_n519), .A2(new_n521), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G85), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  XOR2_X1   g164(.A(KEYINPUT78), .B(G47), .Z(new_n590));
  OAI221_X1 g165(.A(new_n588), .B1(new_n541), .B2(new_n589), .C1(new_n534), .C2(new_n590), .ZN(G290));
  NAND3_X1  g166(.A1(new_n587), .A2(KEYINPUT10), .A3(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n522), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n508), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n538), .A2(G54), .B1(new_n599), .B2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g178(.A(new_n602), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  AOI21_X1  g183(.A(KEYINPUT79), .B1(G299), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n607), .B1(new_n605), .B2(new_n609), .ZN(G297));
  AOI21_X1  g185(.A(new_n607), .B1(new_n605), .B2(new_n609), .ZN(G280));
  INV_X1    g186(.A(new_n601), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  NOR2_X1   g189(.A1(new_n601), .A2(G559), .ZN(new_n615));
  OR3_X1    g190(.A1(new_n615), .A2(KEYINPUT80), .A3(new_n608), .ZN(new_n616));
  OAI21_X1  g191(.A(KEYINPUT80), .B1(new_n615), .B2(new_n608), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n616), .B(new_n617), .C1(G868), .C2(new_n554), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g194(.A1(G123), .A2(new_n488), .B1(new_n486), .B2(G135), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n622));
  INV_X1    g197(.A(G111), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n621), .A2(new_n622), .B1(new_n623), .B2(G2105), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n622), .B2(new_n621), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(G2096), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT81), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n627), .A2(new_n628), .A3(new_n633), .ZN(G156));
  INV_X1    g209(.A(KEYINPUT14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n640), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(G401));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2096), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT20), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n663), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n663), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G229));
  NOR2_X1   g253(.A1(G16), .A2(G23), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT85), .Z(new_n680));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n681));
  XNOR2_X1  g256(.A(G288), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT33), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  MUX2_X1   g261(.A(G6), .B(G305), .S(G16), .Z(new_n687));
  XOR2_X1   g262(.A(KEYINPUT32), .B(G1981), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT84), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n683), .A2(G22), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G166), .B2(new_n683), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1971), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n690), .B2(new_n687), .ZN(new_n695));
  AND3_X1   g270(.A1(new_n686), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT34), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n488), .A2(G119), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n463), .A2(G107), .ZN(new_n701));
  OAI21_X1  g276(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n703));
  AND3_X1   g278(.A1(new_n486), .A2(new_n703), .A3(G131), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n486), .B2(G131), .ZN(new_n705));
  OAI221_X1 g280(.A(new_n700), .B1(new_n701), .B2(new_n702), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G25), .B2(G29), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT35), .B(G1991), .Z(new_n710));
  AND2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n683), .A2(G24), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G290), .B2(G16), .ZN(new_n713));
  INV_X1    g288(.A(G1986), .ZN(new_n714));
  OAI22_X1  g289(.A1(new_n713), .A2(new_n714), .B1(new_n709), .B2(new_n710), .ZN(new_n715));
  AOI211_X1 g290(.A(new_n711), .B(new_n715), .C1(new_n714), .C2(new_n713), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n698), .A2(new_n699), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT36), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT31), .B(G11), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT91), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT30), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n721), .A2(G28), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n707), .B1(new_n721), .B2(G28), .ZN(new_n723));
  OAI221_X1 g298(.A(new_n720), .B1(new_n722), .B2(new_n723), .C1(new_n626), .C2(new_n707), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT92), .Z(new_n725));
  NAND3_X1  g300(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT25), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G139), .B2(new_n486), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n463), .B2(new_n729), .ZN(new_n730));
  MUX2_X1   g305(.A(G33), .B(new_n730), .S(G29), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2072), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT24), .ZN(new_n733));
  INV_X1    g308(.A(G34), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G160), .B2(new_n707), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n725), .B(new_n732), .C1(G2084), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n683), .A2(G20), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT23), .Z(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G299), .B2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1956), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n707), .A2(G27), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G164), .B2(new_n707), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT97), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2078), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n707), .A2(G35), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n707), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT29), .Z(new_n750));
  INV_X1    g325(.A(G2090), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G4), .A2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n612), .B2(G16), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G1348), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n747), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n707), .A2(G26), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT28), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n488), .A2(G128), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT87), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n486), .A2(G140), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n463), .A2(G116), .ZN(new_n762));
  OAI21_X1  g337(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n760), .B(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n758), .B1(new_n764), .B2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2067), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n751), .B2(new_n750), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n683), .A2(G21), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G168), .B2(new_n683), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT90), .B(G1966), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G1348), .B2(new_n754), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n756), .A2(new_n767), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n488), .A2(G129), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT88), .Z(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT26), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n778), .A2(new_n779), .B1(G105), .B2(new_n469), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n486), .A2(G141), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n775), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(new_n707), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n707), .B2(G32), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT27), .B(G1996), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT89), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n683), .A2(G19), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n554), .B2(new_n683), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1341), .Z(new_n791));
  NAND4_X1  g366(.A1(new_n743), .A2(new_n773), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n737), .A2(G2084), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT95), .ZN(new_n794));
  NOR2_X1   g369(.A1(G5), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G171), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT93), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n794), .B1(new_n785), .B2(new_n786), .C1(new_n797), .C2(G1961), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n798), .A2(KEYINPUT96), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(G1961), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT94), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n798), .A2(KEYINPUT96), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n792), .A2(new_n799), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n718), .A2(new_n803), .ZN(G150));
  INV_X1    g379(.A(G150), .ZN(G311));
  NAND2_X1  g380(.A1(new_n587), .A2(G93), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n538), .A2(G55), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(new_n541), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G860), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT37), .Z(new_n812));
  INV_X1    g387(.A(KEYINPUT99), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n553), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g389(.A(KEYINPUT99), .B(new_n547), .C1(new_n551), .C2(new_n552), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n814), .A2(new_n810), .A3(new_n815), .ZN(new_n816));
  OR3_X1    g391(.A1(new_n553), .A2(new_n813), .A3(new_n810), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n612), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n822), .A2(KEYINPUT39), .ZN(new_n823));
  INV_X1    g398(.A(G860), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n822), .B2(KEYINPUT39), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n812), .B1(new_n823), .B2(new_n825), .ZN(G145));
  INV_X1    g401(.A(new_n498), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n465), .B2(new_n466), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n829));
  INV_X1    g404(.A(new_n500), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G114), .B2(new_n463), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(KEYINPUT101), .B1(new_n499), .B2(new_n502), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n497), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n764), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n488), .A2(G130), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n463), .A2(G118), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G142), .B2(new_n486), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n835), .B(new_n840), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n783), .B(new_n730), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n706), .B(new_n632), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n841), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(G162), .B(new_n626), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT100), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G160), .ZN(new_n848));
  AOI21_X1  g423(.A(G37), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n848), .B2(new_n845), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g426(.A(new_n818), .B(new_n615), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n601), .A2(G299), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n601), .A2(G299), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT42), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(KEYINPUT41), .ZN(new_n858));
  OR3_X1    g433(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT41), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n856), .A2(new_n857), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n857), .B1(new_n856), .B2(new_n861), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n682), .B(G303), .ZN(new_n865));
  XNOR2_X1  g440(.A(G305), .B(G290), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n863), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n856), .A2(new_n861), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT42), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n867), .B1(new_n871), .B2(new_n862), .ZN(new_n872));
  OAI21_X1  g447(.A(G868), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n810), .A2(new_n608), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(G295));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n874), .ZN(G331));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n878));
  NAND3_X1  g453(.A1(G171), .A2(G286), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(G301), .A2(G168), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT76), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n536), .B(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(KEYINPUT103), .B1(G301), .B2(new_n883), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n881), .A2(new_n817), .A3(new_n816), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n880), .A3(new_n879), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n818), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n885), .A2(new_n887), .A3(new_n860), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n855), .B1(new_n885), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT104), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n887), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n853), .A2(new_n854), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n885), .A2(new_n887), .A3(new_n860), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n890), .A2(new_n896), .A3(new_n868), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n888), .A2(new_n889), .ZN(new_n898));
  AOI21_X1  g473(.A(G37), .B1(new_n898), .B2(new_n867), .ZN(new_n899));
  XNOR2_X1  g474(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n893), .A2(new_n867), .A3(new_n895), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n858), .A2(new_n905), .A3(new_n859), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n855), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n906), .A2(new_n885), .A3(new_n887), .A4(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n867), .B1(new_n893), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n877), .B1(new_n901), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n900), .B1(new_n897), .B2(new_n899), .ZN(new_n912));
  INV_X1    g487(.A(new_n900), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n904), .A2(new_n913), .A3(new_n909), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n911), .B1(new_n877), .B2(new_n915), .ZN(G397));
  AND2_X1   g491(.A1(new_n467), .A2(new_n470), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n480), .B1(new_n479), .B2(G2105), .ZN(new_n918));
  AOI211_X1 g493(.A(KEYINPUT68), .B(new_n463), .C1(new_n477), .C2(new_n478), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n917), .B(G40), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G1384), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT45), .B1(new_n834), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT106), .ZN(new_n925));
  INV_X1    g500(.A(G2067), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n764), .B(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n783), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n924), .A2(G1996), .ZN(new_n931));
  XOR2_X1   g506(.A(new_n931), .B(KEYINPUT46), .Z(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n933), .B(KEYINPUT47), .Z(new_n934));
  INV_X1    g509(.A(G1996), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n783), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n925), .B1(new_n928), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n931), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n937), .B1(new_n929), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n710), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n706), .A2(new_n940), .ZN(new_n941));
  OAI22_X1  g516(.A1(new_n939), .A2(new_n941), .B1(G2067), .B2(new_n764), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n942), .A2(new_n925), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n706), .B(new_n940), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n939), .B1(new_n925), .B2(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(G290), .A2(new_n924), .A3(G1986), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT127), .Z(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT48), .ZN(new_n948));
  AOI211_X1 g523(.A(new_n934), .B(new_n943), .C1(new_n945), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n834), .A2(new_n922), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(new_n920), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(G8), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n585), .A2(G1981), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n955));
  INV_X1    g530(.A(G1981), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n583), .A2(new_n584), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n585), .A2(KEYINPUT108), .A3(G1981), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n953), .B1(new_n960), .B2(KEYINPUT49), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(new_n955), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n956), .B1(new_n583), .B2(new_n584), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n959), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT109), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n958), .A2(new_n967), .A3(new_n959), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g544(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n970));
  AOI21_X1  g545(.A(KEYINPUT111), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n972));
  INV_X1    g547(.A(new_n970), .ZN(new_n973));
  AOI211_X1 g548(.A(new_n972), .B(new_n973), .C1(new_n966), .C2(new_n968), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n961), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n463), .B(new_n494), .C1(new_n465), .C2(new_n466), .ZN(new_n976));
  INV_X1    g551(.A(new_n495), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n976), .B1(new_n977), .B2(KEYINPUT4), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n828), .A2(new_n831), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n922), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n834), .A2(KEYINPUT45), .A3(new_n922), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n921), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1971), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n950), .A2(KEYINPUT50), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n921), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n834), .B2(new_n922), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT113), .B1(new_n991), .B2(new_n920), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n990), .B(new_n922), .C1(new_n978), .C2(new_n979), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(G1384), .B1(new_n497), .B2(new_n503), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n996), .A2(KEYINPUT114), .A3(new_n990), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n989), .A2(new_n992), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n986), .B1(new_n999), .B2(G2090), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(G8), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G303), .A2(G8), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT55), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(new_n996), .B2(new_n990), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n980), .A2(KEYINPUT107), .A3(KEYINPUT50), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n834), .A2(new_n990), .A3(new_n922), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n921), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n986), .B1(new_n1010), .B2(G2090), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1003), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n951), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n682), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT52), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1018), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1017), .B(new_n1021), .C1(new_n682), .C2(new_n1018), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n975), .A2(new_n1004), .A3(new_n1015), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n984), .ZN(new_n1026));
  INV_X1    g601(.A(G2078), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT53), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1961), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n1029), .B2(new_n1010), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n921), .B1(new_n981), .B2(new_n980), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n923), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1027), .A2(KEYINPUT53), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G171), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1025), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n770), .B1(new_n1031), .B2(new_n923), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT115), .B(G2084), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1008), .A2(new_n1009), .A3(new_n921), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT124), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(new_n1040), .A3(KEYINPUT124), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(G168), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(new_n1016), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1041), .A2(G8), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT51), .B1(new_n536), .B2(G8), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n536), .A2(G8), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT62), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1045), .A2(new_n1047), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT62), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n1054), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1037), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT63), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1041), .A2(G8), .A3(new_n883), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1025), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n961), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n964), .A2(new_n965), .A3(KEYINPUT109), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n967), .B1(new_n958), .B2(new_n959), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n970), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n972), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n969), .A2(KEYINPUT111), .A3(new_n970), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1064), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(new_n1023), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1014), .B1(new_n1012), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1072), .B2(new_n1012), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1062), .A2(new_n1061), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1071), .A2(new_n1015), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1063), .A2(new_n1076), .ZN(new_n1077));
  OR2_X1    g652(.A1(G288), .A2(G1976), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n957), .B1(new_n1070), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT112), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(new_n957), .C1(new_n1070), .C2(new_n1078), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(new_n1017), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1071), .A2(new_n1014), .A3(new_n1013), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1060), .A2(new_n1077), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n567), .A2(new_n1086), .A3(new_n571), .ZN(new_n1087));
  INV_X1    g662(.A(new_n570), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n568), .B(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT57), .B1(new_n1089), .B2(new_n566), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n920), .B1(new_n950), .B2(KEYINPUT50), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1092), .A2(new_n988), .B1(new_n995), .B2(new_n997), .ZN(new_n1093));
  AOI21_X1  g668(.A(G1956), .B1(new_n1093), .B2(new_n992), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT56), .B(G2072), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(KEYINPUT117), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n921), .A2(new_n982), .A3(new_n983), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1091), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1348), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1010), .A2(new_n1100), .B1(new_n926), .B2(new_n951), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n601), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n1103));
  INV_X1    g678(.A(G1956), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n999), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1098), .A2(new_n1091), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1103), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1105), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1102), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(new_n612), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(KEYINPUT60), .B2(new_n1101), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  NAND2_X1  g688(.A1(new_n952), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT120), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1026), .A2(new_n1116), .A3(new_n935), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT119), .B1(new_n984), .B2(G1996), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n952), .A2(new_n1119), .A3(new_n1113), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n554), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1121), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1091), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1105), .B2(new_n1097), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1097), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT61), .B1(new_n1094), .B2(new_n1130), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n1126), .A2(new_n1127), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT118), .B1(new_n1094), .B2(new_n1130), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1105), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1129), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT122), .B1(new_n1135), .B2(KEYINPUT61), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1099), .B1(new_n1108), .B2(new_n1107), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1132), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1112), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AOI211_X1 g718(.A(KEYINPUT123), .B(new_n1132), .C1(new_n1136), .C2(new_n1140), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1109), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(G40), .B1(new_n473), .B2(new_n463), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n923), .A2(new_n471), .A3(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT125), .Z(new_n1148));
  NAND2_X1  g723(.A1(new_n983), .A2(new_n1033), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1030), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(G171), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(G171), .B2(new_n1035), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1030), .A2(G301), .A3(new_n1034), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT126), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1150), .A2(G171), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT54), .ZN(new_n1156));
  OAI22_X1  g731(.A1(new_n1152), .A2(KEYINPUT54), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1057), .A2(new_n1054), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1157), .A2(new_n1025), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1085), .B1(new_n1145), .B2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(G290), .B(new_n714), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n945), .B1(new_n924), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n949), .B1(new_n1160), .B2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g738(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n850), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g740(.A1(new_n915), .A2(new_n1166), .ZN(G308));
  OR2_X1    g741(.A1(new_n915), .A2(new_n1166), .ZN(G225));
endmodule


