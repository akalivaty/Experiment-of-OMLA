//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT72), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT32), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT2), .B(G113), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT70), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT69), .A2(G116), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT69), .A2(G116), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n197), .B1(new_n201), .B2(G119), .ZN(new_n202));
  OR2_X1    g016(.A1(KEYINPUT69), .A2(G116), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n198), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n204), .A2(KEYINPUT70), .A3(new_n195), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n194), .B1(new_n202), .B2(new_n205), .ZN(new_n206));
  OAI211_X1 g020(.A(KEYINPUT70), .B(new_n196), .C1(new_n204), .C2(new_n195), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT70), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n201), .A2(new_n208), .A3(G119), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n193), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G137), .ZN(new_n215));
  INV_X1    g029(.A(G137), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G134), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n215), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n214), .A2(G137), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(KEYINPUT11), .ZN(new_n223));
  OAI211_X1 g037(.A(KEYINPUT67), .B(new_n219), .C1(new_n214), .C2(G137), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n220), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n218), .B1(new_n225), .B2(new_n213), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT64), .B(G146), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT65), .B1(new_n227), .B2(G143), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT64), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(G146), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n228), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n230), .A2(new_n232), .A3(G143), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT1), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G128), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n239), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n229), .A2(G143), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n245), .A3(G128), .A4(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n240), .B1(new_n239), .B2(new_n243), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n226), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT30), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n241), .A2(KEYINPUT0), .A3(G128), .A4(new_n247), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n246), .B1(new_n227), .B2(G143), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n256), .A2(KEYINPUT66), .A3(KEYINPUT0), .A4(G128), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT0), .B(G128), .Z(new_n258));
  AOI22_X1  g072(.A1(new_n255), .A2(new_n257), .B1(new_n239), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n224), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT67), .B1(new_n217), .B2(new_n219), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(G131), .B1(new_n262), .B2(new_n220), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n225), .A2(new_n213), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n252), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n212), .B1(new_n251), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(G143), .B1(new_n230), .B2(new_n232), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n238), .B1(new_n268), .B2(new_n234), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n227), .A2(KEYINPUT65), .A3(G143), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n243), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(new_n248), .A3(new_n244), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n273), .A2(new_n226), .B1(new_n265), .B2(new_n259), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n267), .B1(KEYINPUT30), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n276));
  INV_X1    g090(.A(G237), .ZN(new_n277));
  INV_X1    g091(.A(G953), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n278), .A3(G210), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n279), .B(KEYINPUT27), .Z(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT26), .B(G101), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n282), .B1(new_n274), .B2(new_n212), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n275), .A2(new_n276), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n276), .B1(new_n275), .B2(new_n283), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT28), .ZN(new_n287));
  INV_X1    g101(.A(new_n226), .ZN(new_n288));
  INV_X1    g102(.A(new_n248), .ZN(new_n289));
  INV_X1    g103(.A(G128), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n241), .B2(KEYINPUT1), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n231), .A2(G146), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n229), .A2(KEYINPUT64), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n235), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n237), .B1(new_n294), .B2(KEYINPUT65), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n291), .B1(new_n295), .B2(new_n236), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n289), .B1(new_n296), .B2(new_n240), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n288), .B1(new_n297), .B2(new_n272), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n257), .A2(new_n255), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n239), .A2(new_n258), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n265), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n211), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n251), .A2(new_n212), .A3(new_n301), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n287), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n287), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n282), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n192), .B1(new_n286), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n301), .A2(KEYINPUT30), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n211), .B1(new_n298), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT30), .B1(new_n251), .B2(new_n301), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n282), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n304), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT31), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n275), .A2(new_n276), .A3(new_n283), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n308), .A2(new_n316), .A3(new_n192), .A4(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n191), .B1(new_n309), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G472), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT29), .B1(new_n305), .B2(new_n307), .ZN(new_n322));
  INV_X1    g136(.A(new_n304), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n212), .B1(new_n251), .B2(new_n301), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT28), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n306), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n322), .A2(new_n327), .A3(new_n314), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT73), .B(G902), .Z(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n304), .B(new_n282), .C1(new_n311), .C2(new_n312), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n330), .B1(new_n332), .B2(new_n326), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n321), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n320), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n316), .A2(new_n317), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n314), .B1(new_n325), .B2(new_n306), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT71), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n318), .ZN(new_n340));
  INV_X1    g154(.A(new_n189), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT32), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n187), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G104), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G107), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n344), .A2(G107), .ZN(new_n347));
  OAI21_X1  g161(.A(G101), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT3), .B1(new_n344), .B2(G107), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n350));
  INV_X1    g164(.A(G107), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(G104), .ZN(new_n352));
  INV_X1    g166(.A(G101), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n349), .A2(new_n352), .A3(new_n353), .A4(new_n345), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(KEYINPUT10), .B(new_n356), .C1(new_n249), .C2(new_n250), .ZN(new_n357));
  INV_X1    g171(.A(new_n265), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n349), .A2(new_n352), .A3(new_n345), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G101), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n359), .A2(KEYINPUT81), .A3(new_n360), .A4(G101), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n360), .B1(new_n359), .B2(G101), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n363), .A2(new_n364), .B1(new_n354), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n290), .B1(new_n238), .B2(KEYINPUT1), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n248), .B1(new_n256), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n356), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n259), .A2(new_n366), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n357), .A2(new_n358), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(G110), .B(G140), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n278), .A2(G227), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n358), .B1(new_n357), .B2(new_n371), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n272), .A2(new_n248), .A3(new_n244), .A4(new_n355), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n370), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT12), .B1(new_n381), .B2(new_n265), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT12), .ZN(new_n383));
  AOI211_X1 g197(.A(new_n383), .B(new_n358), .C1(new_n380), .C2(new_n370), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n372), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n379), .B1(new_n385), .B2(new_n375), .ZN(new_n386));
  OAI21_X1  g200(.A(G469), .B1(new_n386), .B2(G902), .ZN(new_n387));
  INV_X1    g201(.A(G469), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n381), .A2(new_n265), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n383), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n381), .A2(KEYINPUT12), .A3(new_n265), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n377), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n378), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n376), .B1(new_n393), .B2(new_n372), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n388), .B(new_n329), .C1(new_n392), .C2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(KEYINPUT82), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n372), .B(new_n376), .C1(new_n382), .C2(new_n384), .ZN(new_n398));
  INV_X1    g212(.A(new_n372), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n375), .B1(new_n399), .B2(new_n378), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n330), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n397), .B1(new_n401), .B2(new_n388), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n387), .B1(new_n396), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G221), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT9), .B(G234), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G902), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G214), .B1(G237), .B2(G902), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G210), .B1(G237), .B2(G902), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n366), .A2(new_n211), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(new_n207), .B2(new_n209), .ZN(new_n417));
  OAI21_X1  g231(.A(G113), .B1(new_n415), .B2(new_n196), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n206), .B(new_n356), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G110), .B(G122), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n414), .A2(new_n421), .A3(new_n419), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(G125), .B1(new_n297), .B2(new_n272), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n259), .A2(G125), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(G224), .B(new_n278), .C1(new_n426), .C2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n420), .A2(new_n430), .A3(new_n422), .ZN(new_n431));
  INV_X1    g245(.A(G125), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n273), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n278), .A2(G224), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n427), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n425), .A2(new_n429), .A3(new_n431), .A4(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(KEYINPUT7), .B(new_n434), .C1(new_n426), .C2(new_n428), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(KEYINPUT7), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n433), .A2(new_n427), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n207), .A2(new_n209), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n418), .B1(new_n441), .B2(new_n415), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n193), .B1(new_n207), .B2(new_n209), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n355), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n206), .A2(new_n356), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n418), .B1(new_n441), .B2(KEYINPUT5), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(new_n421), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n438), .A2(new_n424), .A3(new_n440), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n407), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n413), .B1(new_n437), .B2(new_n452), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n436), .A2(new_n451), .A3(new_n407), .A4(new_n412), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n411), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n403), .A2(new_n409), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n277), .A2(new_n278), .A3(G214), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(G143), .ZN(new_n458));
  AND2_X1   g272(.A1(KEYINPUT18), .A2(G131), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n461));
  INV_X1    g275(.A(G140), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n432), .A2(G140), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT77), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT77), .B1(new_n463), .B2(new_n464), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n227), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT78), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT77), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n432), .A2(G140), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n462), .A2(G125), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT77), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT78), .A3(new_n227), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(KEYINPUT76), .A2(G125), .A3(G140), .ZN(new_n478));
  AOI21_X1  g292(.A(G140), .B1(KEYINPUT76), .B2(G125), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(new_n229), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n461), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  AOI211_X1 g297(.A(KEYINPUT85), .B(new_n481), .C1(new_n469), .C2(new_n476), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n460), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G113), .B(G122), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n344), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT86), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n458), .B(new_n213), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(KEYINPUT17), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT16), .B1(new_n462), .B2(G125), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT16), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n493), .B1(new_n480), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G146), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n478), .A2(new_n479), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n492), .B1(new_n497), .B2(KEYINPUT16), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n229), .ZN(new_n499));
  INV_X1    g313(.A(new_n458), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT17), .A3(G131), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n496), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n485), .B(new_n489), .C1(new_n491), .C2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n487), .ZN(new_n504));
  INV_X1    g318(.A(new_n460), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT78), .B1(new_n475), .B2(new_n227), .ZN(new_n506));
  AOI211_X1 g320(.A(new_n468), .B(new_n233), .C1(new_n473), .C2(new_n474), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n482), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT85), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n477), .A2(new_n461), .A3(new_n482), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n491), .A2(new_n502), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n504), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(G902), .B1(new_n503), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT88), .B(G475), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n511), .A2(new_n512), .A3(new_n488), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n465), .A2(new_n466), .ZN(new_n518));
  MUX2_X1   g332(.A(new_n518), .B(new_n480), .S(KEYINPUT19), .Z(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n227), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n496), .A3(new_n490), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n487), .B1(new_n485), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT87), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n521), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n504), .B1(new_n524), .B2(new_n511), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT87), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n503), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(G475), .A2(G902), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n523), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT20), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n525), .A2(new_n503), .ZN(new_n531));
  NOR3_X1   g345(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n516), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G478), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  INV_X1    g350(.A(G217), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n405), .A2(new_n537), .A3(G953), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n235), .B2(G128), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n290), .A2(KEYINPUT89), .A3(G143), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n540), .A2(new_n541), .B1(G128), .B2(new_n235), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT13), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n214), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n203), .A2(G122), .A3(new_n198), .ZN(new_n545));
  INV_X1    g359(.A(G116), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(G122), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n351), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n351), .B1(new_n545), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n544), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n540), .A2(new_n541), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n235), .A2(G128), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n214), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n543), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT90), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n553), .A2(new_n214), .A3(new_n554), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n549), .B1(new_n560), .B2(new_n555), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n203), .A2(KEYINPUT14), .A3(G122), .A4(new_n198), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G107), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n547), .B1(new_n201), .B2(G122), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT14), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n559), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n553), .A2(new_n554), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G134), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n542), .A2(new_n214), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n545), .A2(new_n548), .ZN(new_n572));
  OAI211_X1 g386(.A(G107), .B(new_n562), .C1(new_n572), .C2(KEYINPUT14), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n571), .A2(new_n573), .A3(KEYINPUT90), .A4(new_n549), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n558), .B1(new_n567), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT91), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n538), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n567), .A2(new_n574), .ZN(new_n578));
  INV_X1    g392(.A(new_n558), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT91), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(KEYINPUT91), .A3(new_n538), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n329), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT92), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT92), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n582), .A2(new_n586), .A3(new_n329), .A4(new_n583), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n536), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n587), .A2(new_n536), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G952), .ZN(new_n591));
  AOI211_X1 g405(.A(G953), .B(new_n591), .C1(G234), .C2(G237), .ZN(new_n592));
  INV_X1    g406(.A(G234), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n330), .B(G953), .C1(new_n593), .C2(new_n277), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT93), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT21), .B(G898), .Z(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT94), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n592), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n534), .A2(new_n590), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n456), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n341), .B1(new_n309), .B2(new_n319), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n190), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n334), .B1(new_n340), .B2(new_n191), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(KEYINPUT74), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT79), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n195), .A2(G128), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n290), .A2(G119), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT24), .B(G110), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT23), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n612), .B1(new_n195), .B2(G128), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n290), .A2(KEYINPUT23), .A3(G119), .ZN(new_n614));
  INV_X1    g428(.A(G110), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .A4(new_n607), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n498), .B2(new_n229), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n469), .B2(new_n476), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n613), .A2(new_n607), .A3(new_n614), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G110), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n609), .B2(new_n610), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n496), .B2(new_n499), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n606), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n496), .B(new_n617), .C1(new_n506), .C2(new_n507), .ZN(new_n625));
  INV_X1    g439(.A(new_n622), .ZN(new_n626));
  INV_X1    g440(.A(new_n499), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n498), .A2(new_n229), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n625), .A2(new_n629), .A3(KEYINPUT79), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT22), .B(G137), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n404), .A2(new_n593), .A3(G953), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n624), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n625), .A2(new_n629), .ZN(new_n635));
  INV_X1    g449(.A(new_n633), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n606), .A3(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n634), .A2(KEYINPUT80), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT80), .B1(new_n634), .B2(new_n637), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n537), .B1(new_n329), .B2(G234), .ZN(new_n640));
  NOR4_X1   g454(.A1(new_n638), .A2(new_n639), .A3(G902), .A4(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n330), .B1(new_n634), .B2(new_n637), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT25), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n640), .B(KEYINPUT75), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n343), .A2(new_n601), .A3(new_n605), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G101), .ZN(G3));
  AOI21_X1  g461(.A(new_n330), .B1(new_n339), .B2(new_n318), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n602), .B1(new_n648), .B2(new_n321), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n403), .A2(new_n645), .A3(new_n409), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n330), .A2(new_n535), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT33), .B1(new_n582), .B2(new_n583), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT33), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT95), .ZN(new_n656));
  OR3_X1    g470(.A1(new_n575), .A2(new_n656), .A3(new_n538), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n538), .B1(new_n575), .B2(new_n656), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n653), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n584), .A2(new_n535), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n529), .A2(KEYINPUT20), .B1(new_n531), .B2(new_n532), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n662), .B1(new_n663), .B2(new_n516), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n451), .A2(new_n407), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n412), .B1(new_n665), .B2(new_n436), .ZN(new_n666));
  INV_X1    g480(.A(new_n454), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n410), .B(new_n599), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n652), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  AOI211_X1 g483(.A(new_n411), .B(new_n598), .C1(new_n453), .C2(new_n454), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n530), .A2(new_n533), .ZN(new_n671));
  INV_X1    g485(.A(new_n516), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n670), .A2(new_n673), .A3(KEYINPUT96), .A4(new_n662), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n651), .A2(new_n669), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT97), .Z(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT34), .B(G104), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  INV_X1    g492(.A(new_n590), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT20), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n523), .A2(new_n527), .A3(new_n680), .A4(new_n528), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n516), .B1(new_n530), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n670), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n649), .A2(new_n650), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT35), .B(G107), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G9));
  NOR2_X1   g500(.A1(new_n633), .A2(KEYINPUT36), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n635), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n640), .A2(G902), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n643), .B2(new_n644), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n602), .B(new_n692), .C1(new_n648), .C2(new_n321), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT98), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n329), .B1(new_n309), .B2(new_n319), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G472), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(KEYINPUT98), .A3(new_n602), .A4(new_n692), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(new_n698), .A3(new_n601), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  INV_X1    g515(.A(G900), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n592), .B1(new_n595), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n682), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n590), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n409), .A2(new_n403), .A3(new_n455), .A4(new_n692), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n343), .A2(new_n605), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  XOR2_X1   g523(.A(new_n703), .B(KEYINPUT39), .Z(new_n710));
  NAND3_X1  g524(.A1(new_n403), .A2(new_n409), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT40), .Z(new_n712));
  NAND2_X1  g526(.A1(new_n275), .A2(new_n304), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n314), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n323), .A2(new_n324), .ZN(new_n715));
  AOI21_X1  g529(.A(G902), .B1(new_n715), .B2(new_n282), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n321), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n340), .B2(new_n191), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n692), .B1(new_n603), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n666), .A2(new_n667), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT38), .ZN(new_n721));
  NOR4_X1   g535(.A1(new_n721), .A2(new_n411), .A3(new_n590), .A4(new_n534), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n712), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n235), .ZN(G45));
  AOI22_X1  g538(.A1(new_n671), .A2(new_n672), .B1(new_n661), .B2(new_n660), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n704), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n343), .A2(new_n605), .A3(new_n707), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT99), .B(G146), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G48));
  NAND2_X1  g544(.A1(new_n343), .A2(new_n605), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n395), .A2(KEYINPUT82), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n401), .A2(new_n397), .A3(new_n388), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n401), .A2(new_n388), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n734), .A2(new_n645), .A3(new_n409), .A4(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n674), .A3(new_n669), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n731), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT41), .B(G113), .Z(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT100), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n739), .B(new_n741), .ZN(G15));
  NOR2_X1   g556(.A1(new_n683), .A2(new_n736), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n343), .A2(new_n743), .A3(new_n605), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G116), .ZN(G18));
  NAND4_X1  g559(.A1(new_n734), .A2(new_n455), .A3(new_n409), .A4(new_n735), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n746), .A2(new_n600), .A3(new_n691), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n343), .A2(new_n747), .A3(new_n605), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G119), .ZN(G21));
  INV_X1    g563(.A(KEYINPUT103), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n534), .B2(new_n590), .ZN(new_n751));
  OAI221_X1 g565(.A(KEYINPUT103), .B1(new_n588), .B2(new_n589), .C1(new_n663), .C2(new_n516), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n751), .A2(new_n752), .A3(new_n455), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT101), .B1(new_n305), .B2(new_n307), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n282), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT101), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n286), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n341), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT102), .B(G472), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n645), .B(new_n758), .C1(new_n648), .C2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n734), .A2(new_n735), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n763), .A2(new_n408), .A3(new_n598), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n753), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G122), .ZN(G24));
  AOI22_X1  g580(.A1(new_n696), .A2(new_n759), .B1(new_n341), .B2(new_n757), .ZN(new_n767));
  INV_X1    g581(.A(new_n746), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n727), .A2(new_n692), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G125), .ZN(G27));
  NAND2_X1  g584(.A1(new_n385), .A2(new_n375), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT105), .ZN(new_n772));
  INV_X1    g586(.A(new_n379), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT105), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n385), .A2(new_n774), .A3(new_n375), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n772), .A2(G469), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(G469), .A2(G902), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT104), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n776), .B(new_n779), .C1(new_n396), .C2(new_n402), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n666), .A2(new_n667), .A3(new_n408), .A4(new_n411), .ZN(new_n781));
  AND4_X1   g595(.A1(new_n725), .A2(new_n780), .A3(new_n704), .A4(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(KEYINPUT42), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n603), .A2(new_n604), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n645), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT107), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT107), .B1(new_n784), .B2(new_n645), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n343), .A2(new_n782), .A3(new_n605), .A4(new_n645), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT106), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT42), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n790), .B2(KEYINPUT106), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n789), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G131), .ZN(G33));
  NAND3_X1  g609(.A1(new_n343), .A2(new_n645), .A3(new_n605), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT108), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n705), .B2(new_n590), .ZN(new_n798));
  AOI211_X1 g612(.A(new_n516), .B(new_n703), .C1(new_n530), .C2(new_n681), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n679), .A3(KEYINPUT108), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n780), .A3(new_n781), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(new_n214), .ZN(G36));
  AND3_X1   g617(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT45), .ZN(new_n805));
  OAI211_X1 g619(.A(KEYINPUT109), .B(G469), .C1(new_n386), .C2(KEYINPUT45), .ZN(new_n806));
  OAI21_X1  g620(.A(G469), .B1(new_n386), .B2(KEYINPUT45), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT109), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n805), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT110), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n804), .A2(KEYINPUT45), .B1(new_n808), .B2(new_n807), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n813), .A3(new_n806), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n778), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT112), .B1(new_n815), .B2(KEYINPUT46), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n814), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT46), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n778), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT111), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n821));
  INV_X1    g635(.A(new_n819), .ZN(new_n822));
  AOI211_X1 g636(.A(new_n821), .B(new_n822), .C1(new_n811), .C2(new_n814), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n816), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n817), .A2(new_n779), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n826), .A3(new_n818), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n734), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n409), .B(new_n710), .C1(new_n824), .C2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n534), .A2(new_n662), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT43), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n649), .A3(new_n692), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT44), .ZN(new_n836));
  OR3_X1    g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n835), .B1(new_n834), .B2(new_n836), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n666), .A2(new_n411), .A3(new_n667), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n834), .B2(new_n836), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n830), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(G137), .ZN(G39));
  OAI21_X1  g658(.A(new_n409), .B1(new_n824), .B2(new_n828), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT47), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT47), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n847), .B(new_n409), .C1(new_n824), .C2(new_n828), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n726), .A2(new_n645), .A3(new_n841), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n731), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(G140), .ZN(G42));
  NAND4_X1  g666(.A1(new_n721), .A2(new_n645), .A3(new_n409), .A4(new_n410), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n831), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n603), .A2(new_n718), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n763), .B(KEYINPUT49), .Z(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n763), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n846), .A2(new_n848), .B1(new_n408), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n833), .A2(new_n592), .A3(new_n762), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n840), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n763), .A2(new_n408), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n860), .A2(new_n411), .A3(new_n721), .A4(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT50), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n841), .A2(new_n763), .A3(new_n408), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n855), .A2(new_n645), .A3(new_n592), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n870), .A2(new_n673), .A3(new_n662), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n833), .A2(new_n592), .A3(new_n867), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n872), .A2(new_n692), .A3(new_n767), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n866), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT51), .A4(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n874), .B1(new_n859), .B2(new_n861), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT119), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n785), .B(new_n786), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n872), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT48), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n591), .B(G953), .C1(new_n860), .C2(new_n768), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n881), .B(new_n882), .C1(new_n664), .C2(new_n870), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n876), .B2(new_n877), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n875), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n691), .A2(new_n588), .A3(new_n589), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n799), .A2(new_n887), .A3(new_n840), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n403), .A2(new_n409), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n343), .A2(new_n890), .A3(new_n605), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n782), .A2(new_n692), .A3(new_n767), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n891), .B(new_n892), .C1(new_n796), .C2(new_n801), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n725), .A2(KEYINPUT115), .A3(new_n670), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT115), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n895), .B1(new_n664), .B2(new_n668), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n670), .A2(new_n679), .A3(new_n534), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n651), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n646), .A2(new_n699), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n744), .B1(new_n731), .B2(new_n738), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n748), .A2(new_n765), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT114), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n737), .A2(new_n674), .A3(new_n669), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n343), .B(new_n605), .C1(new_n905), .C2(new_n743), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT114), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n906), .A2(new_n907), .A3(new_n748), .A4(new_n765), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n901), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  AND4_X1   g723(.A1(new_n645), .A2(new_n343), .A3(new_n782), .A4(new_n605), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT106), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT42), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n790), .A2(KEYINPUT106), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n912), .A2(new_n913), .B1(new_n879), .B2(new_n783), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n708), .A2(new_n769), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n780), .A2(new_n409), .A3(new_n704), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n753), .A2(new_n719), .A3(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n916), .A2(KEYINPUT52), .A3(new_n728), .A4(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n708), .A2(new_n728), .A3(new_n918), .A4(new_n769), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT52), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n915), .B(new_n923), .C1(KEYINPUT116), .C2(KEYINPUT53), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n904), .A2(new_n908), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n925), .A2(new_n923), .A3(new_n794), .A4(new_n901), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT53), .B1(new_n923), .B2(KEYINPUT116), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n886), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT53), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n794), .A2(new_n904), .A3(new_n908), .A4(new_n901), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n920), .B(KEYINPUT52), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n902), .A2(new_n903), .A3(new_n930), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n923), .A2(new_n794), .A3(new_n901), .A4(new_n934), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n933), .A2(new_n886), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT117), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n926), .A2(new_n927), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n926), .A2(new_n927), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT54), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT117), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n933), .A2(new_n886), .A3(new_n935), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n885), .B1(new_n937), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(G952), .A2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n857), .B1(new_n944), .B2(new_n945), .ZN(G75));
  NOR2_X1   g760(.A1(new_n278), .A2(G952), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n933), .A2(new_n935), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(new_n329), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT56), .B1(new_n950), .B2(new_n413), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n425), .A2(new_n431), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n429), .A2(new_n435), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n436), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT55), .Z(new_n956));
  OAI21_X1  g770(.A(new_n948), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n951), .B2(new_n956), .ZN(G51));
  XNOR2_X1  g772(.A(new_n778), .B(KEYINPUT57), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT120), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n933), .A2(new_n960), .A3(new_n886), .A4(new_n935), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n949), .B2(new_n886), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n942), .A2(KEYINPUT120), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n959), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n392), .B2(new_n394), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n950), .A2(new_n814), .A3(new_n811), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n947), .B1(new_n966), .B2(new_n967), .ZN(G54));
  NAND2_X1  g782(.A1(new_n523), .A2(new_n527), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(KEYINPUT58), .A2(G475), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n950), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n950), .B2(new_n971), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n972), .A2(new_n973), .A3(new_n947), .ZN(G60));
  NAND2_X1  g788(.A1(new_n582), .A2(new_n583), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n659), .B1(new_n975), .B2(new_n655), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT121), .ZN(new_n977));
  NAND2_X1  g791(.A1(G478), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT59), .Z(new_n979));
  NOR2_X1   g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n886), .B1(new_n933), .B2(new_n935), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n936), .B2(new_n960), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n983), .B2(new_n963), .ZN(new_n984));
  OAI21_X1  g798(.A(KEYINPUT122), .B1(new_n984), .B2(new_n947), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n980), .B1(new_n962), .B2(new_n964), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT122), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n986), .A2(new_n987), .A3(new_n948), .ZN(new_n988));
  INV_X1    g802(.A(new_n979), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n943), .A2(new_n937), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n977), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n985), .A2(new_n988), .A3(new_n991), .ZN(G63));
  OAI21_X1  g806(.A(new_n948), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n993));
  NAND2_X1  g807(.A1(G217), .A2(G902), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT60), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n949), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n993), .B1(new_n996), .B2(new_n688), .ZN(new_n997));
  OAI22_X1  g811(.A1(new_n949), .A2(new_n995), .B1(new_n638), .B2(new_n639), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(G66));
  INV_X1    g815(.A(G224), .ZN(new_n1002));
  OAI21_X1  g816(.A(G953), .B1(new_n597), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n925), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1004), .A2(new_n900), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1003), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n952), .B1(G898), .B2(new_n278), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT124), .Z(new_n1008));
  XNOR2_X1  g822(.A(new_n1006), .B(new_n1008), .ZN(G69));
  INV_X1    g823(.A(KEYINPUT125), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n846), .A2(new_n848), .A3(new_n850), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n916), .A2(new_n728), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1012), .A2(new_n802), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n787), .A2(new_n788), .ZN(new_n1014));
  INV_X1    g828(.A(new_n753), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1016), .B1(new_n839), .B2(new_n842), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n794), .B(new_n1013), .C1(new_n1017), .C2(new_n829), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1010), .B1(new_n1011), .B2(new_n1018), .ZN(new_n1019));
  OR2_X1    g833(.A1(new_n1017), .A2(new_n829), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n1013), .A2(new_n794), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1020), .A2(new_n851), .A3(KEYINPUT125), .A4(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1019), .A2(new_n278), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n312), .B1(new_n251), .B2(new_n266), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(new_n519), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n1023), .B(new_n1025), .C1(new_n702), .C2(new_n278), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1012), .A2(new_n723), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT62), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n725), .B1(new_n679), .B2(new_n534), .ZN(new_n1029));
  OR4_X1    g843(.A1(new_n796), .A2(new_n711), .A3(new_n841), .A4(new_n1029), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1028), .A2(new_n843), .A3(new_n851), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n278), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1025), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1026), .A2(new_n1034), .ZN(new_n1035));
  OR2_X1    g849(.A1(new_n1033), .A2(KEYINPUT126), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n278), .B1(G227), .B2(G900), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1026), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(new_n1041), .ZN(G72));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT63), .Z(new_n1044));
  INV_X1    g858(.A(new_n1005), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1044), .B1(new_n1031), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1046), .A2(new_n314), .A3(new_n713), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n938), .A2(new_n939), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n714), .A2(new_n331), .A3(new_n1044), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n1019), .A2(new_n1005), .A3(new_n1022), .ZN(new_n1051));
  AND2_X1   g865(.A1(new_n1051), .A2(new_n1044), .ZN(new_n1052));
  OAI211_X1 g866(.A(KEYINPUT127), .B(new_n948), .C1(new_n1052), .C2(new_n331), .ZN(new_n1053));
  INV_X1    g867(.A(KEYINPUT127), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n331), .B1(new_n1051), .B2(new_n1044), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1054), .B1(new_n1055), .B2(new_n947), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1050), .B1(new_n1053), .B2(new_n1056), .ZN(G57));
endmodule


