

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593;

  XNOR2_X1 U322 ( .A(n411), .B(n410), .ZN(n414) );
  XOR2_X1 U323 ( .A(G169GAT), .B(G8GAT), .Z(n324) );
  XNOR2_X1 U324 ( .A(n403), .B(n402), .ZN(n404) );
  NOR2_X1 U325 ( .A1(n416), .A2(n415), .ZN(n418) );
  XNOR2_X1 U326 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n480) );
  XOR2_X1 U327 ( .A(KEYINPUT28), .B(n475), .Z(n540) );
  XOR2_X1 U328 ( .A(n323), .B(n322), .Z(n530) );
  AND2_X1 U329 ( .A1(n473), .A2(n472), .ZN(n290) );
  AND2_X1 U330 ( .A1(G229GAT), .A2(G233GAT), .ZN(n291) );
  AND2_X1 U331 ( .A1(G226GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U332 ( .A(n345), .B(KEYINPUT74), .ZN(n346) );
  XNOR2_X1 U333 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n410) );
  XNOR2_X1 U334 ( .A(n431), .B(n346), .ZN(n349) );
  INV_X1 U335 ( .A(KEYINPUT11), .ZN(n400) );
  XNOR2_X1 U336 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n417) );
  XNOR2_X1 U337 ( .A(n329), .B(n291), .ZN(n330) );
  XNOR2_X1 U338 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U339 ( .A(n324), .B(n292), .ZN(n317) );
  XNOR2_X1 U340 ( .A(n331), .B(n330), .ZN(n335) );
  XNOR2_X1 U341 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U342 ( .A(n454), .B(n317), .ZN(n319) );
  XNOR2_X1 U343 ( .A(n361), .B(n360), .ZN(n412) );
  XNOR2_X1 U344 ( .A(n481), .B(n480), .ZN(n526) );
  XOR2_X1 U345 ( .A(n343), .B(n342), .Z(n578) );
  INV_X1 U346 ( .A(G43GAT), .ZN(n484) );
  XNOR2_X1 U347 ( .A(n483), .B(KEYINPUT38), .ZN(n514) );
  XNOR2_X1 U348 ( .A(n488), .B(G190GAT), .ZN(n489) );
  XNOR2_X1 U349 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U350 ( .A(n490), .B(n489), .ZN(G1351GAT) );
  XNOR2_X1 U351 ( .A(n487), .B(n486), .ZN(G1330GAT) );
  INV_X1 U352 ( .A(KEYINPUT122), .ZN(n460) );
  XOR2_X1 U353 ( .A(KEYINPUT18), .B(KEYINPUT88), .Z(n294) );
  XNOR2_X1 U354 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n293) );
  XNOR2_X1 U355 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U356 ( .A(KEYINPUT19), .B(n295), .Z(n321) );
  XOR2_X1 U357 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n297) );
  XNOR2_X1 U358 ( .A(G120GAT), .B(KEYINPUT87), .ZN(n296) );
  XNOR2_X1 U359 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U360 ( .A(KEYINPUT89), .B(G71GAT), .Z(n299) );
  XNOR2_X1 U361 ( .A(KEYINPUT84), .B(G176GAT), .ZN(n298) );
  XNOR2_X1 U362 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U363 ( .A(n301), .B(n300), .Z(n312) );
  XOR2_X1 U364 ( .A(G127GAT), .B(KEYINPUT86), .Z(n303) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(G15GAT), .ZN(n302) );
  XNOR2_X1 U366 ( .A(n303), .B(n302), .ZN(n310) );
  XOR2_X1 U367 ( .A(G113GAT), .B(KEYINPUT0), .Z(n436) );
  XOR2_X1 U368 ( .A(G190GAT), .B(G134GAT), .Z(n305) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(G99GAT), .ZN(n304) );
  XNOR2_X1 U370 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U371 ( .A(n436), .B(n306), .Z(n308) );
  NAND2_X1 U372 ( .A1(G227GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U373 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U374 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U375 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U376 ( .A(n321), .B(n313), .Z(n539) );
  INV_X1 U377 ( .A(n539), .ZN(n533) );
  XOR2_X1 U378 ( .A(G211GAT), .B(G218GAT), .Z(n315) );
  XNOR2_X1 U379 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U380 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U381 ( .A(G197GAT), .B(n316), .Z(n454) );
  XNOR2_X1 U382 ( .A(G176GAT), .B(G92GAT), .ZN(n318) );
  XNOR2_X1 U383 ( .A(n318), .B(G64GAT), .ZN(n348) );
  XOR2_X1 U384 ( .A(n319), .B(n348), .Z(n323) );
  XNOR2_X1 U385 ( .A(G36GAT), .B(G190GAT), .ZN(n320) );
  XNOR2_X1 U386 ( .A(n320), .B(KEYINPUT81), .ZN(n399) );
  XNOR2_X1 U387 ( .A(n321), .B(n399), .ZN(n322) );
  INV_X1 U388 ( .A(n530), .ZN(n419) );
  XOR2_X1 U389 ( .A(G36GAT), .B(G29GAT), .Z(n326) );
  XOR2_X1 U390 ( .A(G15GAT), .B(G22GAT), .Z(n375) );
  XNOR2_X1 U391 ( .A(n375), .B(n324), .ZN(n325) );
  XNOR2_X1 U392 ( .A(n326), .B(n325), .ZN(n331) );
  XOR2_X1 U393 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n328) );
  XNOR2_X1 U394 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n327) );
  XNOR2_X1 U395 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U396 ( .A(G1GAT), .B(G141GAT), .Z(n333) );
  XNOR2_X1 U397 ( .A(G113GAT), .B(G197GAT), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U399 ( .A(n335), .B(n334), .Z(n343) );
  XOR2_X1 U400 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n337) );
  XNOR2_X1 U401 ( .A(G50GAT), .B(G43GAT), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U403 ( .A(KEYINPUT7), .B(n338), .Z(n396) );
  XOR2_X1 U404 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n340) );
  XNOR2_X1 U405 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n339) );
  XNOR2_X1 U406 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U407 ( .A(n396), .B(n341), .ZN(n342) );
  INV_X1 U408 ( .A(n578), .ZN(n572) );
  XNOR2_X1 U409 ( .A(G120GAT), .B(G148GAT), .ZN(n344) );
  XNOR2_X1 U410 ( .A(n344), .B(G57GAT), .ZN(n431) );
  AND2_X1 U411 ( .A1(G230GAT), .A2(G233GAT), .ZN(n345) );
  INV_X1 U412 ( .A(n349), .ZN(n347) );
  NAND2_X1 U413 ( .A1(n347), .A2(n348), .ZN(n352) );
  INV_X1 U414 ( .A(n348), .ZN(n350) );
  NAND2_X1 U415 ( .A1(n350), .A2(n349), .ZN(n351) );
  NAND2_X1 U416 ( .A1(n352), .A2(n351), .ZN(n354) );
  XOR2_X1 U417 ( .A(G106GAT), .B(G78GAT), .Z(n443) );
  XOR2_X1 U418 ( .A(G99GAT), .B(G85GAT), .Z(n392) );
  XNOR2_X1 U419 ( .A(n443), .B(n392), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U421 ( .A(n355), .B(KEYINPUT33), .Z(n361) );
  XOR2_X1 U422 ( .A(G71GAT), .B(KEYINPUT13), .Z(n365) );
  XNOR2_X1 U423 ( .A(G204GAT), .B(n365), .ZN(n359) );
  XOR2_X1 U424 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n357) );
  XNOR2_X1 U425 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n356) );
  XNOR2_X1 U426 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n412), .B(KEYINPUT41), .ZN(n561) );
  NOR2_X1 U428 ( .A1(n572), .A2(n561), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n362), .B(KEYINPUT46), .ZN(n383) );
  XOR2_X1 U430 ( .A(G78GAT), .B(G155GAT), .Z(n364) );
  XNOR2_X1 U431 ( .A(G183GAT), .B(G211GAT), .ZN(n363) );
  XNOR2_X1 U432 ( .A(n364), .B(n363), .ZN(n379) );
  XOR2_X1 U433 ( .A(G1GAT), .B(G127GAT), .Z(n429) );
  XOR2_X1 U434 ( .A(n365), .B(n429), .Z(n367) );
  NAND2_X1 U435 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U437 ( .A(KEYINPUT15), .B(G64GAT), .Z(n369) );
  XNOR2_X1 U438 ( .A(KEYINPUT82), .B(KEYINPUT14), .ZN(n368) );
  XNOR2_X1 U439 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U440 ( .A(n371), .B(n370), .Z(n377) );
  XOR2_X1 U441 ( .A(KEYINPUT83), .B(KEYINPUT12), .Z(n373) );
  XNOR2_X1 U442 ( .A(G8GAT), .B(G57GAT), .ZN(n372) );
  XNOR2_X1 U443 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U445 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U446 ( .A(n379), .B(n378), .Z(n564) );
  INV_X1 U447 ( .A(n564), .ZN(n587) );
  OR2_X1 U448 ( .A1(n383), .A2(n587), .ZN(n381) );
  INV_X1 U449 ( .A(KEYINPUT110), .ZN(n380) );
  NAND2_X1 U450 ( .A1(n381), .A2(n380), .ZN(n385) );
  NAND2_X1 U451 ( .A1(n564), .A2(KEYINPUT110), .ZN(n382) );
  OR2_X1 U452 ( .A1(n383), .A2(n382), .ZN(n384) );
  NAND2_X1 U453 ( .A1(n385), .A2(n384), .ZN(n406) );
  XOR2_X1 U454 ( .A(KEYINPUT78), .B(KEYINPUT66), .Z(n387) );
  XNOR2_X1 U455 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U457 ( .A(KEYINPUT64), .B(KEYINPUT79), .Z(n389) );
  XNOR2_X1 U458 ( .A(G92GAT), .B(KEYINPUT80), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U460 ( .A(n391), .B(n390), .ZN(n405) );
  XNOR2_X1 U461 ( .A(KEYINPUT9), .B(n392), .ZN(n394) );
  XOR2_X1 U462 ( .A(G29GAT), .B(G134GAT), .Z(n432) );
  XNOR2_X1 U463 ( .A(G218GAT), .B(n432), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U465 ( .A(n396), .B(n395), .ZN(n398) );
  NAND2_X1 U466 ( .A1(G232GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U467 ( .A(n398), .B(n397), .ZN(n403) );
  XNOR2_X1 U468 ( .A(G162GAT), .B(n399), .ZN(n401) );
  XOR2_X1 U469 ( .A(n405), .B(n404), .Z(n494) );
  INV_X1 U470 ( .A(n494), .ZN(n569) );
  NAND2_X1 U471 ( .A1(n406), .A2(n569), .ZN(n409) );
  XOR2_X1 U472 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n407) );
  XNOR2_X1 U473 ( .A(KEYINPUT47), .B(n407), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n409), .B(n408), .ZN(n416) );
  XNOR2_X1 U475 ( .A(KEYINPUT36), .B(n494), .ZN(n590) );
  NAND2_X1 U476 ( .A1(n587), .A2(n590), .ZN(n411) );
  NOR2_X1 U477 ( .A1(n412), .A2(n578), .ZN(n413) );
  AND2_X1 U478 ( .A1(n414), .A2(n413), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n541) );
  NAND2_X1 U480 ( .A1(n419), .A2(n541), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n420), .B(KEYINPUT121), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n421), .B(KEYINPUT54), .ZN(n575) );
  XOR2_X1 U483 ( .A(KEYINPUT2), .B(G162GAT), .Z(n423) );
  XNOR2_X1 U484 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U486 ( .A(G141GAT), .B(n424), .ZN(n450) );
  INV_X1 U487 ( .A(n450), .ZN(n442) );
  XOR2_X1 U488 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n426) );
  XNOR2_X1 U489 ( .A(KEYINPUT92), .B(KEYINPUT6), .ZN(n425) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n440) );
  XOR2_X1 U491 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n428) );
  XNOR2_X1 U492 ( .A(G85GAT), .B(KEYINPUT4), .ZN(n427) );
  XNOR2_X1 U493 ( .A(n428), .B(n427), .ZN(n430) );
  XOR2_X1 U494 ( .A(n430), .B(n429), .Z(n438) );
  XOR2_X1 U495 ( .A(n431), .B(n432), .Z(n434) );
  NAND2_X1 U496 ( .A1(G225GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U497 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U500 ( .A(n440), .B(n439), .Z(n441) );
  XOR2_X1 U501 ( .A(n442), .B(n441), .Z(n471) );
  XNOR2_X1 U502 ( .A(KEYINPUT93), .B(n471), .ZN(n574) );
  XOR2_X1 U503 ( .A(G148GAT), .B(n443), .Z(n445) );
  NAND2_X1 U504 ( .A1(G228GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U506 ( .A(n446), .B(KEYINPUT23), .Z(n452) );
  XOR2_X1 U507 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n448) );
  XNOR2_X1 U508 ( .A(G50GAT), .B(G22GAT), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U510 ( .A(n450), .B(n449), .Z(n451) );
  XNOR2_X1 U511 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n475) );
  INV_X1 U513 ( .A(n475), .ZN(n455) );
  AND2_X1 U514 ( .A1(n574), .A2(n455), .ZN(n456) );
  AND2_X1 U515 ( .A1(n575), .A2(n456), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n457), .B(KEYINPUT55), .ZN(n458) );
  NOR2_X1 U517 ( .A1(n533), .A2(n458), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n460), .B(n459), .ZN(n571) );
  NOR2_X1 U519 ( .A1(n571), .A2(n564), .ZN(n462) );
  INV_X1 U520 ( .A(G183GAT), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n462), .B(n461), .ZN(G1350GAT) );
  NOR2_X1 U522 ( .A1(n533), .A2(n530), .ZN(n463) );
  NOR2_X1 U523 ( .A1(n475), .A2(n463), .ZN(n464) );
  XOR2_X1 U524 ( .A(n464), .B(KEYINPUT96), .Z(n465) );
  XNOR2_X1 U525 ( .A(KEYINPUT25), .B(n465), .ZN(n469) );
  NAND2_X1 U526 ( .A1(n475), .A2(n533), .ZN(n466) );
  XNOR2_X1 U527 ( .A(KEYINPUT26), .B(n466), .ZN(n576) );
  XNOR2_X1 U528 ( .A(n530), .B(KEYINPUT27), .ZN(n474) );
  NOR2_X1 U529 ( .A1(n576), .A2(n474), .ZN(n467) );
  XOR2_X1 U530 ( .A(KEYINPUT95), .B(n467), .Z(n468) );
  NOR2_X1 U531 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n470), .B(KEYINPUT97), .ZN(n473) );
  INV_X1 U533 ( .A(n471), .ZN(n472) );
  NOR2_X1 U534 ( .A1(n474), .A2(n574), .ZN(n542) );
  NAND2_X1 U535 ( .A1(n542), .A2(n540), .ZN(n476) );
  XNOR2_X1 U536 ( .A(KEYINPUT94), .B(n476), .ZN(n477) );
  NOR2_X1 U537 ( .A1(n539), .A2(n477), .ZN(n478) );
  NOR2_X1 U538 ( .A1(n290), .A2(n478), .ZN(n497) );
  NOR2_X1 U539 ( .A1(n497), .A2(n587), .ZN(n479) );
  NAND2_X1 U540 ( .A1(n479), .A2(n590), .ZN(n481) );
  NOR2_X1 U541 ( .A1(n572), .A2(n412), .ZN(n482) );
  XOR2_X1 U542 ( .A(KEYINPUT77), .B(n482), .Z(n498) );
  NAND2_X1 U543 ( .A1(n526), .A2(n498), .ZN(n483) );
  NOR2_X1 U544 ( .A1(n514), .A2(n533), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n485) );
  NOR2_X1 U546 ( .A1(n569), .A2(n571), .ZN(n490) );
  XNOR2_X1 U547 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n488) );
  NOR2_X1 U548 ( .A1(n561), .A2(n571), .ZN(n493) );
  XNOR2_X1 U549 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n491), .B(G176GAT), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(G1349GAT) );
  NOR2_X1 U552 ( .A1(n564), .A2(n494), .ZN(n495) );
  XOR2_X1 U553 ( .A(KEYINPUT16), .B(n495), .Z(n496) );
  NOR2_X1 U554 ( .A1(n497), .A2(n496), .ZN(n517) );
  NAND2_X1 U555 ( .A1(n498), .A2(n517), .ZN(n499) );
  XNOR2_X1 U556 ( .A(KEYINPUT98), .B(n499), .ZN(n507) );
  NOR2_X1 U557 ( .A1(n507), .A2(n574), .ZN(n500) );
  XOR2_X1 U558 ( .A(KEYINPUT34), .B(n500), .Z(n501) );
  XNOR2_X1 U559 ( .A(G1GAT), .B(n501), .ZN(G1324GAT) );
  NOR2_X1 U560 ( .A1(n507), .A2(n530), .ZN(n503) );
  XNOR2_X1 U561 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U563 ( .A(G8GAT), .B(n504), .ZN(G1325GAT) );
  NOR2_X1 U564 ( .A1(n507), .A2(n533), .ZN(n506) );
  XNOR2_X1 U565 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(G1326GAT) );
  NOR2_X1 U567 ( .A1(n507), .A2(n540), .ZN(n509) );
  XNOR2_X1 U568 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n508) );
  XNOR2_X1 U569 ( .A(n509), .B(n508), .ZN(G1327GAT) );
  NOR2_X1 U570 ( .A1(n514), .A2(n574), .ZN(n511) );
  XNOR2_X1 U571 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n511), .B(n510), .ZN(G1328GAT) );
  NOR2_X1 U573 ( .A1(n514), .A2(n530), .ZN(n513) );
  XNOR2_X1 U574 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n513), .B(n512), .ZN(G1329GAT) );
  NOR2_X1 U576 ( .A1(n514), .A2(n540), .ZN(n515) );
  XOR2_X1 U577 ( .A(G50GAT), .B(n515), .Z(G1331GAT) );
  NOR2_X1 U578 ( .A1(n561), .A2(n578), .ZN(n516) );
  XOR2_X1 U579 ( .A(KEYINPUT105), .B(n516), .Z(n527) );
  NAND2_X1 U580 ( .A1(n517), .A2(n527), .ZN(n523) );
  NOR2_X1 U581 ( .A1(n574), .A2(n523), .ZN(n518) );
  XOR2_X1 U582 ( .A(G57GAT), .B(n518), .Z(n519) );
  XNOR2_X1 U583 ( .A(KEYINPUT42), .B(n519), .ZN(G1332GAT) );
  NOR2_X1 U584 ( .A1(n530), .A2(n523), .ZN(n520) );
  XOR2_X1 U585 ( .A(KEYINPUT106), .B(n520), .Z(n521) );
  XNOR2_X1 U586 ( .A(G64GAT), .B(n521), .ZN(G1333GAT) );
  NOR2_X1 U587 ( .A1(n533), .A2(n523), .ZN(n522) );
  XOR2_X1 U588 ( .A(G71GAT), .B(n522), .Z(G1334GAT) );
  NOR2_X1 U589 ( .A1(n540), .A2(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  NAND2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n535) );
  NOR2_X1 U593 ( .A1(n574), .A2(n535), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(G1336GAT) );
  NOR2_X1 U596 ( .A1(n530), .A2(n535), .ZN(n531) );
  XOR2_X1 U597 ( .A(KEYINPUT108), .B(n531), .Z(n532) );
  XNOR2_X1 U598 ( .A(G92GAT), .B(n532), .ZN(G1337GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n535), .ZN(n534) );
  XOR2_X1 U600 ( .A(G99GAT), .B(n534), .Z(G1338GAT) );
  NOR2_X1 U601 ( .A1(n540), .A2(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT109), .B(KEYINPUT44), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  AND2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U607 ( .A(KEYINPUT114), .B(n543), .Z(n555) );
  NAND2_X1 U608 ( .A1(n544), .A2(n555), .ZN(n551) );
  NOR2_X1 U609 ( .A1(n572), .A2(n551), .ZN(n545) );
  XOR2_X1 U610 ( .A(G113GAT), .B(n545), .Z(G1340GAT) );
  NOR2_X1 U611 ( .A1(n561), .A2(n551), .ZN(n547) );
  XNOR2_X1 U612 ( .A(KEYINPUT49), .B(KEYINPUT115), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U614 ( .A(G120GAT), .B(n548), .Z(G1341GAT) );
  NOR2_X1 U615 ( .A1(n564), .A2(n551), .ZN(n549) );
  XOR2_X1 U616 ( .A(KEYINPUT50), .B(n549), .Z(n550) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  NOR2_X1 U618 ( .A1(n569), .A2(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n558) );
  INV_X1 U622 ( .A(n576), .ZN(n554) );
  NAND2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(KEYINPUT116), .ZN(n568) );
  NOR2_X1 U625 ( .A1(n572), .A2(n568), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n560) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n559) );
  XNOR2_X1 U629 ( .A(n560), .B(n559), .ZN(n563) );
  NOR2_X1 U630 ( .A1(n561), .A2(n568), .ZN(n562) );
  XOR2_X1 U631 ( .A(n563), .B(n562), .Z(G1345GAT) );
  XNOR2_X1 U632 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n566) );
  NOR2_X1 U633 ( .A1(n564), .A2(n568), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(G155GAT), .B(n567), .ZN(G1346GAT) );
  NOR2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U637 ( .A(G162GAT), .B(n570), .Z(G1347GAT) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(G169GAT), .B(n573), .Z(G1348GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n577) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n591) );
  AND2_X1 U642 ( .A1(n578), .A2(n591), .ZN(n583) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n580) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(KEYINPUT124), .B(n581), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U649 ( .A1(n591), .A2(n412), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(n586), .ZN(G1353GAT) );
  XOR2_X1 U652 ( .A(G211GAT), .B(KEYINPUT127), .Z(n589) );
  NAND2_X1 U653 ( .A1(n591), .A2(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1354GAT) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(n592), .B(KEYINPUT62), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

