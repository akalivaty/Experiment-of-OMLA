//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n606, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1223, new_n1224, new_n1225;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(G2106), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G137), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n461), .A2(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n460), .A2(new_n462), .B1(new_n463), .B2(G101), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(new_n461), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G160));
  NOR2_X1   g042(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(new_n461), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  AND2_X1   g057(.A1(G126), .A2(G2105), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n461), .A2(G114), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n460), .A2(new_n483), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n489), .B(new_n490), .C1(new_n470), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n490), .B1(new_n460), .B2(new_n489), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n487), .B(KEYINPUT68), .C1(new_n493), .C2(new_n494), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  OAI21_X1  g075(.A(G543), .B1(KEYINPUT72), .B2(KEYINPUT5), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(KEYINPUT72), .B2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT70), .B(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n507), .A2(KEYINPUT70), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(KEYINPUT70), .ZN(new_n509));
  OAI211_X1 g084(.A(KEYINPUT71), .B(KEYINPUT5), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n502), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n517), .A2(new_n507), .ZN(new_n521));
  AOI21_X1  g096(.A(KEYINPUT69), .B1(new_n521), .B2(G50), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n521), .A2(KEYINPUT69), .A3(G50), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n519), .A2(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n514), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT73), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT7), .Z(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(G51), .B2(new_n521), .ZN(new_n529));
  AOI211_X1 g104(.A(new_n502), .B(new_n517), .C1(new_n506), .C2(new_n510), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n513), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n521), .A2(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n519), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(new_n511), .A2(G56), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n513), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n545), .B1(new_n544), .B2(new_n543), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n530), .A2(G81), .B1(G43), .B2(new_n521), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n553), .B(KEYINPUT75), .Z(G188));
  NAND2_X1  g129(.A1(new_n521), .A2(G53), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n530), .A2(G91), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n556), .B(new_n557), .C1(new_n558), .C2(new_n513), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G166), .ZN(G303));
  NAND2_X1  g136(.A1(new_n530), .A2(G87), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n521), .A2(G49), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  NAND2_X1  g140(.A1(new_n506), .A2(new_n510), .ZN(new_n566));
  INV_X1    g141(.A(new_n502), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n566), .A2(G86), .A3(new_n567), .A4(new_n518), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n521), .A2(G48), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G61), .ZN(new_n571));
  AOI211_X1 g146(.A(new_n571), .B(new_n502), .C1(new_n506), .C2(new_n510), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n570), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g152(.A(KEYINPUT76), .B(G651), .C1(new_n572), .C2(new_n574), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G305));
  NAND2_X1  g154(.A1(new_n521), .A2(G47), .ZN(new_n580));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n519), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n582), .A2(KEYINPUT77), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(KEYINPUT77), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n583), .A2(new_n584), .B1(new_n513), .B2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n519), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n530), .A2(KEYINPUT10), .A3(G92), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n590), .A2(new_n591), .B1(G54), .B2(new_n521), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n511), .A2(G66), .ZN(new_n593));
  AND2_X1   g168(.A1(G79), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT78), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n594), .B1(new_n511), .B2(G66), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n513), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n592), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n587), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n587), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(KEYINPUT79), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n604), .A2(KEYINPUT79), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n605), .B1(new_n606), .B2(new_n608), .ZN(G297));
  AOI21_X1  g184(.A(new_n605), .B1(new_n606), .B2(new_n608), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n601), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n601), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n548), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT80), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n475), .A2(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n477), .A2(G123), .ZN(new_n619));
  OR2_X1    g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n620), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n460), .A2(new_n463), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n628), .A2(KEYINPUT81), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n626), .B1(KEYINPUT81), .B2(new_n628), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n623), .B(new_n630), .C1(new_n631), .C2(new_n629), .ZN(G156));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G14), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT82), .ZN(new_n651));
  NOR2_X1   g226(.A1(G2072), .A2(G2078), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n442), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n649), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(KEYINPUT17), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n649), .B(new_n650), .C1(new_n442), .C2(new_n652), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n651), .A3(new_n649), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n628), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT83), .B(G2096), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n666), .A2(KEYINPUT84), .ZN(new_n667));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(KEYINPUT84), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n664), .A2(new_n665), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(new_n666), .ZN(new_n674));
  MUX2_X1   g249(.A(new_n674), .B(new_n673), .S(new_n669), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G229));
  MUX2_X1   g257(.A(G6), .B(G305), .S(G16), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT87), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT32), .B(G1981), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n686), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n689), .ZN(new_n691));
  INV_X1    g266(.A(G1971), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(G16), .A2(G23), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT88), .Z(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G288), .B2(new_n689), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT33), .ZN(new_n697));
  INV_X1    g272(.A(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND4_X1  g274(.A1(new_n687), .A2(new_n688), .A3(new_n693), .A4(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n702));
  MUX2_X1   g277(.A(G24), .B(G290), .S(G16), .Z(new_n703));
  INV_X1    g278(.A(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G25), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT85), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n477), .A2(G119), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n461), .A2(G107), .ZN(new_n710));
  OAI21_X1  g285(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n711));
  AND3_X1   g286(.A1(new_n475), .A2(KEYINPUT86), .A3(G131), .ZN(new_n712));
  AOI21_X1  g287(.A(KEYINPUT86), .B1(new_n475), .B2(G131), .ZN(new_n713));
  OAI221_X1 g288(.A(new_n709), .B1(new_n710), .B2(new_n711), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n708), .B1(new_n714), .B2(G29), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n715), .B(new_n717), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n701), .A2(new_n702), .A3(new_n705), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT36), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n706), .A2(G27), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G164), .B2(new_n706), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT97), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT96), .B(G2078), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G29), .A2(G33), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT91), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT25), .Z(new_n729));
  AOI22_X1  g304(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  INV_X1    g305(.A(new_n475), .ZN(new_n731));
  INV_X1    g306(.A(G139), .ZN(new_n732));
  OAI221_X1 g307(.A(new_n729), .B1(new_n461), .B2(new_n730), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n727), .B1(new_n733), .B2(new_n706), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2072), .ZN(new_n735));
  INV_X1    g310(.A(G2084), .ZN(new_n736));
  INV_X1    g311(.A(G34), .ZN(new_n737));
  AOI21_X1  g312(.A(G29), .B1(new_n737), .B2(KEYINPUT24), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(KEYINPUT24), .B2(new_n737), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n466), .B2(new_n706), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n735), .B1(new_n736), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n706), .A2(G32), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n460), .B(KEYINPUT67), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n743), .A2(G141), .A3(new_n461), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n743), .A2(G129), .A3(G2105), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT26), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n748), .A2(new_n749), .B1(G105), .B2(new_n463), .ZN(new_n750));
  AND3_X1   g325(.A1(new_n744), .A2(new_n745), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n742), .B1(new_n751), .B2(new_n706), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT27), .B(G1996), .Z(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n741), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n725), .B1(new_n755), .B2(KEYINPUT92), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n706), .A2(G35), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G162), .B2(new_n706), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT29), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G2090), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT98), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n689), .A2(G4), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n601), .B2(new_n689), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1348), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n689), .A2(G5), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G171), .B2(new_n689), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT94), .Z(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n765), .B1(new_n769), .B2(G1961), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n622), .A2(G29), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT30), .B(G28), .Z(new_n772));
  NOR2_X1   g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  AND2_X1   g348(.A1(KEYINPUT31), .A2(G11), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n771), .B1(G29), .B2(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT93), .ZN(new_n776));
  NAND2_X1  g351(.A1(G286), .A2(G16), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n689), .A2(G21), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n776), .B1(G1966), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n706), .A2(G26), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT28), .Z(new_n783));
  OAI211_X1 g358(.A(G140), .B(new_n461), .C1(new_n468), .C2(new_n473), .ZN(new_n784));
  OAI211_X1 g359(.A(G128), .B(G2105), .C1(new_n468), .C2(new_n473), .ZN(new_n785));
  OR2_X1    g360(.A1(G104), .A2(G2105), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n786), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n783), .B1(new_n788), .B2(G29), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT90), .B(G2067), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G1966), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n791), .B1(new_n779), .B2(new_n792), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n781), .B(new_n793), .C1(G2090), .C2(new_n759), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n689), .A2(G20), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT23), .ZN(new_n796));
  INV_X1    g371(.A(G299), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n689), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1956), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n755), .A2(KEYINPUT92), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n794), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n689), .A2(G19), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT89), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n548), .B2(new_n689), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G1341), .Z(new_n805));
  NAND4_X1  g380(.A1(new_n762), .A2(new_n770), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n752), .A2(new_n753), .B1(new_n736), .B2(new_n740), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n769), .B2(G1961), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT95), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n720), .A2(new_n810), .ZN(G311));
  NAND2_X1  g386(.A1(new_n720), .A2(new_n810), .ZN(G150));
  NAND2_X1  g387(.A1(new_n521), .A2(G55), .ZN(new_n813));
  INV_X1    g388(.A(G93), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n519), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n511), .A2(G67), .ZN(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n513), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n815), .A2(new_n818), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT99), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n546), .A2(new_n547), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n548), .A2(new_n822), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n600), .A2(new_n611), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n832), .A2(new_n833), .A3(G860), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n824), .A2(G860), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  NAND2_X1  g412(.A1(new_n475), .A2(G142), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n477), .A2(G130), .ZN(new_n839));
  OR2_X1    g414(.A1(G106), .A2(G2105), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n840), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n489), .B1(new_n491), .B2(new_n470), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT4), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n846), .A2(KEYINPUT100), .A3(new_n492), .ZN(new_n847));
  AOI21_X1  g422(.A(KEYINPUT100), .B1(new_n846), .B2(new_n492), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n487), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n487), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n493), .B2(new_n494), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n846), .A2(KEYINPUT100), .A3(new_n492), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n788), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n850), .A2(new_n751), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n751), .B1(new_n850), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT101), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n850), .A2(new_n856), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n744), .A2(new_n745), .A3(new_n750), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n864), .A3(new_n857), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n733), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n733), .A3(new_n857), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT102), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI211_X1 g444(.A(KEYINPUT102), .B(new_n733), .C1(new_n860), .C2(new_n865), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n843), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n714), .B(new_n625), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n873));
  INV_X1    g448(.A(new_n733), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT101), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n864), .B1(new_n863), .B2(new_n857), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n873), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n877), .B(new_n842), .C1(new_n866), .C2(new_n868), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n871), .A2(new_n872), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n872), .B1(new_n871), .B2(new_n878), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n622), .B(G160), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n481), .ZN(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n885));
  INV_X1    g460(.A(new_n872), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(KEYINPUT102), .A3(new_n867), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n842), .B1(new_n888), .B2(new_n877), .ZN(new_n889));
  INV_X1    g464(.A(new_n878), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n871), .A2(new_n872), .A3(new_n878), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n883), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n885), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI211_X1 g470(.A(KEYINPUT103), .B(new_n883), .C1(new_n891), .C2(new_n892), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n884), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g473(.A(new_n828), .B(new_n613), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n600), .A2(new_n797), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n600), .A2(KEYINPUT104), .A3(new_n797), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n600), .A2(new_n797), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n899), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n905), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n902), .A2(KEYINPUT41), .A3(new_n903), .A4(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT41), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n902), .A2(KEYINPUT105), .A3(new_n903), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT104), .B1(new_n600), .B2(new_n797), .ZN(new_n915));
  AOI211_X1 g490(.A(new_n901), .B(G299), .C1(new_n592), .C2(new_n599), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n917), .A3(new_n909), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n911), .B1(new_n912), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n908), .B1(new_n919), .B2(new_n899), .ZN(new_n920));
  XNOR2_X1  g495(.A(G290), .B(G303), .ZN(new_n921));
  XNOR2_X1  g496(.A(G288), .B(KEYINPUT106), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(G305), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n922), .A2(G305), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n923), .ZN(new_n926));
  XNOR2_X1  g501(.A(G290), .B(G166), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT42), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n920), .B(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(new_n607), .ZN(new_n932));
  AOI21_X1  g507(.A(G868), .B1(new_n821), .B2(new_n823), .ZN(new_n933));
  OR3_X1    g508(.A1(new_n932), .A2(KEYINPUT107), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT107), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(G295));
  OR2_X1    g511(.A1(new_n932), .A2(new_n933), .ZN(G331));
  XNOR2_X1  g512(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n918), .A2(new_n912), .ZN(new_n940));
  XNOR2_X1  g515(.A(G301), .B(G286), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n826), .A2(new_n941), .A3(new_n827), .ZN(new_n942));
  XNOR2_X1  g517(.A(G286), .B(G171), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n825), .A2(new_n819), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n821), .A2(new_n823), .B1(new_n546), .B2(new_n547), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n940), .A2(new_n910), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n929), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n942), .A2(new_n946), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n906), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n949), .B1(new_n948), .B2(new_n951), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n939), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n942), .A2(new_n946), .A3(KEYINPUT41), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n929), .B1(new_n906), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n947), .A2(KEYINPUT41), .A3(new_n918), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n948), .A2(new_n951), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n960), .B(new_n938), .C1(new_n961), .C2(new_n949), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n956), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(KEYINPUT44), .ZN(new_n964));
  INV_X1    g539(.A(new_n960), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT43), .B1(new_n965), .B2(new_n955), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n954), .A2(new_n955), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n966), .B1(new_n967), .B2(new_n939), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n964), .B1(KEYINPUT44), .B2(new_n968), .ZN(G397));
  INV_X1    g544(.A(KEYINPUT125), .ZN(new_n970));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n849), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT109), .B(G40), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n466), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n714), .B(new_n717), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT110), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n862), .B(G1996), .ZN(new_n982));
  INV_X1    g557(.A(G2067), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n844), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n788), .A2(G2067), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n981), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(G290), .B(new_n704), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n979), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(G166), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT55), .B(G8), .C1(new_n514), .C2(new_n524), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n849), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n853), .A2(new_n854), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n1000), .B2(new_n487), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(KEYINPUT111), .A3(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n497), .A2(new_n971), .A3(new_n498), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n977), .B1(new_n1004), .B2(new_n973), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1971), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n497), .A2(KEYINPUT50), .A3(new_n971), .A4(new_n498), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1008));
  INV_X1    g583(.A(G2090), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n976), .ZN(new_n1010));
  OAI211_X1 g585(.A(G8), .B(new_n996), .C1(new_n1006), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT49), .ZN(new_n1012));
  INV_X1    g587(.A(G1981), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n577), .B2(new_n578), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n574), .B1(new_n511), .B2(G61), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n576), .B1(new_n1015), .B2(new_n513), .ZN(new_n1016));
  INV_X1    g591(.A(new_n570), .ZN(new_n1017));
  AND4_X1   g592(.A1(new_n1013), .A2(new_n1016), .A3(new_n578), .A4(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1012), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1020));
  INV_X1    g595(.A(new_n578), .ZN(new_n1021));
  OAI21_X1  g596(.A(G1981), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n577), .A2(new_n1013), .A3(new_n578), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(KEYINPUT49), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n972), .A2(new_n977), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT112), .B1(new_n1025), .B2(new_n993), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1001), .A2(new_n976), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(G8), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1019), .A2(new_n1024), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G288), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G1976), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT52), .B1(G288), .B2(new_n698), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1028), .B1(new_n1027), .B2(G8), .ZN(new_n1036));
  AOI211_X1 g611(.A(KEYINPUT112), .B(new_n993), .C1(new_n1001), .C2(new_n976), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1033), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT52), .ZN(new_n1039));
  AND4_X1   g614(.A1(new_n1011), .A2(new_n1031), .A3(new_n1035), .A4(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n971), .A4(new_n498), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n976), .B(new_n1041), .C1(new_n1001), .C2(KEYINPUT45), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n977), .A2(G2084), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1042), .A2(new_n792), .B1(new_n1008), .B2(new_n1043), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1044), .A2(new_n993), .A3(G286), .ZN(new_n1045));
  OAI21_X1  g620(.A(G8), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1046));
  INV_X1    g621(.A(new_n996), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1040), .A2(KEYINPUT63), .A3(new_n1045), .A4(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1011), .A2(new_n1031), .A3(new_n1035), .A4(new_n1039), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n497), .A2(new_n1051), .A3(new_n971), .A4(new_n498), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n976), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1051), .B1(new_n849), .B2(new_n971), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1053), .A2(new_n1054), .A3(G2090), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT111), .B1(new_n1001), .B2(KEYINPUT45), .ZN(new_n1056));
  NOR4_X1   g631(.A1(new_n855), .A2(new_n998), .A3(new_n973), .A4(G1384), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1005), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1055), .B1(new_n1058), .B2(new_n692), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT113), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1006), .B2(new_n1055), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1060), .A2(new_n1062), .A3(G8), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1050), .B1(new_n1047), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT114), .B1(new_n1064), .B2(new_n1045), .ZN(new_n1065));
  OAI21_X1  g640(.A(G8), .B1(new_n1059), .B2(KEYINPUT113), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1006), .A2(new_n1061), .A3(new_n1055), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1047), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1040), .A2(new_n1068), .A3(KEYINPUT114), .A4(new_n1045), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT63), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1049), .B1(new_n1065), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n993), .B1(new_n1044), .B2(G168), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1042), .A2(new_n792), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1008), .A2(new_n1043), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G286), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1073), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1075), .A2(G168), .A3(new_n1076), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G8), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(KEYINPUT51), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT62), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1058), .B2(G2078), .ZN(new_n1085));
  OR3_X1    g660(.A1(new_n1042), .A2(new_n1084), .A3(G2078), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1008), .A2(new_n976), .ZN(new_n1087));
  INV_X1    g662(.A(G1961), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G171), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1044), .A2(G168), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT51), .B1(new_n1081), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1074), .A2(new_n1073), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1083), .A2(new_n1092), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1040), .A2(new_n1068), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT123), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1091), .B1(new_n1101), .B2(KEYINPUT62), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(new_n1064), .A3(new_n1103), .A4(new_n1097), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1031), .A2(new_n698), .A3(new_n1032), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1023), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1031), .A2(new_n1039), .A3(new_n1035), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1011), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1107), .A2(new_n1030), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1072), .A2(new_n1105), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n556), .B2(KEYINPUT117), .ZN(new_n1112));
  XNOR2_X1  g687(.A(G299), .B(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1003), .A2(new_n1005), .A3(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n976), .B(new_n1052), .C1(new_n1001), .C2(new_n1051), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT115), .B(G1956), .Z(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(KEYINPUT116), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT116), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1113), .B(new_n1115), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1025), .A2(new_n983), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1008), .A2(new_n976), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1123), .B2(G1348), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT118), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1126), .B(new_n1122), .C1(new_n1123), .C2(G1348), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT119), .B1(new_n1128), .B2(new_n600), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1117), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT116), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1118), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1115), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1113), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1129), .A2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1128), .A2(KEYINPUT119), .A3(new_n600), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1121), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1125), .A2(new_n1140), .A3(new_n1127), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n600), .B1(new_n1128), .B2(KEYINPUT60), .ZN(new_n1142));
  AOI211_X1 g717(.A(new_n1140), .B(new_n601), .C1(new_n1125), .C2(new_n1127), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1121), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1113), .B1(new_n1133), .B2(new_n1115), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT61), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1136), .A2(new_n1148), .A3(new_n1121), .ZN(new_n1149));
  INV_X1    g724(.A(G1996), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1150), .B(new_n1005), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT58), .B(G1341), .Z(new_n1152));
  NAND2_X1  g727(.A1(new_n1027), .A2(new_n1152), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1151), .A2(KEYINPUT120), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT120), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n548), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1158), .B(new_n548), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1147), .A2(new_n1149), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1144), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1163), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1139), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT54), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1168));
  INV_X1    g743(.A(G40), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1084), .A2(new_n1169), .A3(G2078), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1003), .A2(G160), .A3(new_n974), .A4(new_n1170), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1168), .A2(G301), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1167), .B1(new_n1172), .B2(new_n1092), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1173), .A2(new_n1064), .A3(new_n1101), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1090), .A2(G171), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT122), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1167), .B1(new_n1177), .B2(G171), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1174), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1166), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n991), .B1(new_n1111), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n978), .A2(new_n1150), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT46), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n978), .B1(new_n862), .B2(new_n986), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT47), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n714), .A2(new_n717), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n984), .B1(new_n988), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n978), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n979), .A2(G290), .A3(G1986), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(KEYINPUT48), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1191), .B1(new_n989), .B2(new_n979), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1190), .A2(KEYINPUT48), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1186), .B(new_n1189), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1194), .B(KEYINPUT124), .Z(new_n1195));
  OAI21_X1  g770(.A(new_n970), .B1(new_n1181), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(new_n991), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1198), .A2(new_n1173), .A3(new_n1064), .A4(new_n1101), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT121), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1201), .A2(new_n1202), .A3(new_n1144), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1199), .B1(new_n1203), .B2(new_n1139), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1072), .A2(new_n1105), .A3(new_n1110), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1197), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1194), .B(KEYINPUT124), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1206), .A2(KEYINPUT125), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1196), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g784(.A(KEYINPUT126), .ZN(new_n1211));
  OAI21_X1  g785(.A(G319), .B1(new_n646), .B2(new_n647), .ZN(new_n1212));
  NOR3_X1   g786(.A1(G229), .A2(G227), .A3(new_n1212), .ZN(new_n1213));
  AND4_X1   g787(.A1(new_n1211), .A2(new_n963), .A3(new_n897), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g788(.A(new_n1213), .ZN(new_n1215));
  OAI21_X1  g789(.A(new_n894), .B1(new_n879), .B2(new_n880), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1216), .A2(KEYINPUT103), .ZN(new_n1217));
  NAND3_X1  g791(.A1(new_n893), .A2(new_n885), .A3(new_n894), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g793(.A(new_n1215), .B1(new_n1219), .B2(new_n884), .ZN(new_n1220));
  AOI21_X1  g794(.A(new_n1211), .B1(new_n1220), .B2(new_n963), .ZN(new_n1221));
  NOR2_X1   g795(.A1(new_n1214), .A2(new_n1221), .ZN(G308));
  NAND3_X1  g796(.A1(new_n963), .A2(new_n897), .A3(new_n1213), .ZN(new_n1223));
  NAND2_X1  g797(.A1(new_n1223), .A2(KEYINPUT126), .ZN(new_n1224));
  NAND3_X1  g798(.A1(new_n1220), .A2(new_n1211), .A3(new_n963), .ZN(new_n1225));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n1225), .ZN(G225));
endmodule


