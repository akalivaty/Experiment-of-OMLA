//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1224, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND3_X1  g0012(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n224), .A2(new_n225), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n212), .B(new_n221), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT66), .Z(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G232), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G1698), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n251), .B1(G226), .B2(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G97), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(new_n214), .B2(new_n215), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT13), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G1), .A2(G13), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n266), .B1(new_n268), .B2(new_n257), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n265), .A2(G238), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n260), .A2(new_n261), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n258), .B1(new_n254), .B2(new_n255), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n272), .A2(new_n262), .A3(G274), .ZN(new_n276));
  INV_X1    g0076(.A(G238), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n276), .B1(new_n264), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT13), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G200), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G68), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n282), .A2(G50), .B1(G20), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G77), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n207), .A2(G33), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT64), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n267), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(new_n213), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT11), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G13), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n295), .A2(new_n207), .A3(G1), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n283), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT12), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n287), .A2(KEYINPUT11), .A3(new_n291), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n291), .A2(new_n296), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n206), .A2(G20), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(G68), .A3(new_n301), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n294), .A2(new_n298), .A3(new_n299), .A4(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n274), .A2(new_n279), .A3(G190), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n281), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n300), .A2(G50), .A3(new_n301), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n296), .A2(new_n202), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT8), .B(G58), .ZN(new_n310));
  INV_X1    g0110(.A(G150), .ZN(new_n311));
  INV_X1    g0111(.A(new_n282), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n310), .A2(new_n286), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(G20), .B2(new_n203), .ZN(new_n314));
  INV_X1    g0114(.A(new_n291), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n308), .B(new_n309), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT9), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G226), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n276), .B1(new_n264), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT3), .ZN(new_n321));
  INV_X1    g0121(.A(G33), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  AOI21_X1  g0124(.A(G1698), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G222), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n324), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(G223), .A3(G1698), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n326), .B(new_n328), .C1(new_n285), .C2(new_n327), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n320), .B1(new_n329), .B2(new_n259), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT67), .B(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(G190), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT10), .B1(new_n318), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n316), .B(KEYINPUT9), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT10), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n337), .A2(new_n333), .A3(new_n338), .A4(new_n334), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n331), .A2(G179), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n316), .B1(new_n330), .B2(G169), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n280), .A2(G169), .ZN(new_n346));
  NAND2_X1  g0146(.A1(KEYINPUT69), .A2(KEYINPUT14), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n274), .A2(new_n279), .A3(G179), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n261), .B1(new_n260), .B2(new_n273), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n275), .A2(new_n278), .A3(KEYINPUT13), .ZN(new_n352));
  OAI211_X1 g0152(.A(G169), .B(new_n347), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n349), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  AOI211_X1 g0154(.A(new_n307), .B(new_n345), .C1(new_n303), .C2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT17), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n327), .B2(G20), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n252), .A2(new_n253), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n283), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G58), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(new_n283), .ZN(new_n364));
  OAI21_X1  g0164(.A(G20), .B1(new_n364), .B2(new_n201), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n282), .A2(G159), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n357), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT7), .B1(new_n360), .B2(new_n207), .ZN(new_n369));
  NOR4_X1   g0169(.A1(new_n252), .A2(new_n253), .A3(new_n358), .A4(G20), .ZN(new_n370));
  OAI21_X1  g0170(.A(G68), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n367), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(KEYINPUT16), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n368), .A2(new_n373), .A3(new_n291), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n310), .B1(new_n206), .B2(G20), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n300), .A2(new_n375), .B1(new_n296), .B2(new_n310), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n319), .A2(G1698), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n377), .B1(G223), .B2(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G87), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n259), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n276), .B1(new_n264), .B2(new_n250), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G190), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G200), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n258), .B1(new_n378), .B2(new_n379), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n382), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n374), .A2(new_n376), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT70), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT70), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n374), .A2(new_n389), .A3(new_n392), .A4(new_n376), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n356), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n376), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n371), .A2(new_n372), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n315), .B1(new_n396), .B2(new_n357), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n395), .B1(new_n397), .B2(new_n373), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n387), .A2(new_n382), .ZN(new_n399));
  INV_X1    g0199(.A(G179), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G169), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n387), .B2(new_n382), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT18), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n374), .A2(new_n376), .ZN(new_n406));
  INV_X1    g0206(.A(new_n404), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT17), .B1(new_n398), .B2(new_n389), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n394), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G20), .A2(G77), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT15), .B(G87), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n413), .B1(new_n310), .B2(new_n312), .C1(new_n286), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n291), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n300), .A2(G77), .A3(new_n301), .ZN(new_n417));
  INV_X1    g0217(.A(new_n296), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(G77), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n416), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G1698), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n327), .A2(G232), .A3(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(G238), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n360), .A2(G107), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n259), .ZN(new_n427));
  INV_X1    g0227(.A(G244), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n276), .B1(new_n264), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n332), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n421), .A2(new_n432), .A3(KEYINPUT68), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n419), .B1(new_n415), .B2(new_n291), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n429), .B1(new_n426), .B2(new_n259), .ZN(new_n435));
  INV_X1    g0235(.A(new_n332), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n434), .B(new_n417), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT68), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n435), .A2(G190), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n433), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n431), .A2(new_n402), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n434), .A2(new_n417), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n435), .A2(new_n400), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n355), .A2(new_n412), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT5), .ZN(new_n448));
  OR3_X1    g0248(.A1(new_n448), .A2(KEYINPUT74), .A3(G41), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT74), .B1(new_n448), .B2(G41), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n269), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n206), .B(G45), .C1(new_n270), .C2(KEYINPUT5), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT72), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n448), .A2(G41), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT72), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(new_n206), .A4(G45), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n454), .A2(KEYINPUT73), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT73), .B1(new_n454), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n452), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n327), .A2(G264), .A3(G1698), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n327), .A2(G257), .A3(new_n422), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n360), .A2(G303), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n259), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n454), .A2(new_n457), .A3(new_n449), .A4(new_n450), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(G270), .A3(new_n262), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n460), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n206), .A2(G33), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n300), .A2(G116), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n296), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(G20), .B1(G33), .B2(G283), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n322), .A2(G97), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n473), .A2(new_n474), .B1(G20), .B2(new_n471), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n475), .A2(new_n291), .A3(KEYINPUT20), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT20), .B1(new_n475), .B2(new_n291), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n470), .B(new_n472), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G169), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT21), .B1(new_n468), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n460), .A2(new_n465), .A3(new_n467), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT21), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n481), .A2(new_n482), .A3(G169), .A4(new_n478), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT78), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n468), .A2(new_n485), .A3(G179), .A4(new_n478), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n460), .A2(new_n465), .A3(G179), .A4(new_n467), .ZN(new_n487));
  INV_X1    g0287(.A(new_n478), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT78), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n478), .B1(new_n481), .B2(G200), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n384), .B2(new_n481), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n484), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT23), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(G20), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT79), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n494), .A2(new_n497), .A3(new_n498), .A4(KEYINPUT79), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n207), .B(G87), .C1(new_n252), .C2(new_n253), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT22), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n327), .A2(new_n506), .A3(new_n207), .A4(G87), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT80), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT24), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n501), .A2(new_n502), .B1(new_n505), .B2(new_n507), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT24), .B1(new_n512), .B2(KEYINPUT80), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n503), .A2(new_n508), .A3(KEYINPUT80), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n511), .B(new_n291), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n300), .A2(new_n469), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n496), .B1(KEYINPUT81), .B2(KEYINPUT25), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n418), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n296), .A2(KEYINPUT81), .A3(KEYINPUT25), .A4(new_n496), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n517), .A2(G107), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n466), .A2(G264), .A3(new_n262), .ZN(new_n523));
  OAI211_X1 g0323(.A(G257), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n524));
  OAI211_X1 g0324(.A(G250), .B(new_n422), .C1(new_n252), .C2(new_n253), .ZN(new_n525));
  INV_X1    g0325(.A(G294), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n524), .B(new_n525), .C1(new_n322), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n259), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n460), .A2(G190), .A3(new_n523), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n460), .A2(new_n523), .A3(new_n528), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G200), .ZN(new_n531));
  AND4_X1   g0331(.A1(new_n515), .A2(new_n522), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n523), .A2(new_n528), .ZN(new_n533));
  INV_X1    g0333(.A(new_n459), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n454), .A2(KEYINPUT73), .A3(new_n457), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n451), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n402), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n460), .A2(new_n400), .A3(new_n523), .A4(new_n528), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n515), .B2(new_n522), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n532), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G283), .ZN(new_n542));
  OAI211_X1 g0342(.A(G250), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n543));
  OAI211_X1 g0343(.A(G244), .B(new_n422), .C1(new_n252), .C2(new_n253), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT4), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n542), .B(new_n543), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT4), .B1(new_n325), .B2(G244), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n259), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n466), .A2(G257), .A3(new_n262), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n460), .A2(new_n548), .A3(new_n384), .A4(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n460), .A2(new_n548), .A3(new_n549), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(G200), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n418), .A2(G97), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G97), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n516), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n496), .B1(new_n359), .B2(new_n361), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT71), .ZN(new_n558));
  OAI21_X1  g0358(.A(G107), .B1(new_n369), .B2(new_n370), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT71), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n282), .A2(G77), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT6), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n563), .A2(new_n555), .A3(G107), .ZN(new_n564));
  XNOR2_X1  g0364(.A(G97), .B(G107), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G20), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n558), .A2(new_n561), .A3(new_n562), .A4(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n556), .B1(new_n569), .B2(new_n291), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n552), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT19), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n207), .B1(new_n255), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G87), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(new_n555), .A3(new_n496), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n207), .B(G68), .C1(new_n252), .C2(new_n253), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n572), .B1(new_n286), .B2(new_n555), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n291), .ZN(new_n580));
  INV_X1    g0380(.A(new_n414), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n300), .A2(new_n581), .A3(new_n469), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n414), .A2(new_n296), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT76), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n579), .A2(new_n291), .B1(new_n296), .B2(new_n414), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT76), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n582), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(G250), .ZN(new_n590));
  OAI22_X1  g0390(.A1(KEYINPUT75), .A2(new_n590), .B1(new_n271), .B2(G1), .ZN(new_n591));
  NAND2_X1  g0391(.A1(KEYINPUT75), .A2(G250), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n592), .A2(new_n206), .A3(G45), .A4(new_n266), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n591), .A2(new_n593), .A3(new_n262), .ZN(new_n594));
  OAI211_X1 g0394(.A(G238), .B(new_n422), .C1(new_n252), .C2(new_n253), .ZN(new_n595));
  OAI211_X1 g0395(.A(G244), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n595), .B(new_n596), .C1(new_n322), .C2(new_n471), .ZN(new_n597));
  AOI211_X1 g0397(.A(G179), .B(new_n594), .C1(new_n597), .C2(new_n259), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n259), .ZN(new_n599));
  INV_X1    g0399(.A(new_n594), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n598), .B1(new_n402), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n594), .B1(new_n597), .B2(new_n259), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(new_n436), .ZN(new_n604));
  AOI211_X1 g0404(.A(new_n384), .B(new_n594), .C1(new_n597), .C2(new_n259), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n580), .A2(new_n583), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT77), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n516), .B2(new_n574), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n300), .A2(KEYINPUT77), .A3(G87), .A4(new_n469), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n589), .A2(new_n602), .B1(new_n606), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n460), .A2(new_n548), .A3(new_n400), .A4(new_n549), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n460), .A2(new_n548), .A3(new_n549), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n402), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n562), .B1(new_n566), .B2(new_n207), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(KEYINPUT71), .B2(new_n557), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n315), .B1(new_n617), .B2(new_n561), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n613), .B(new_n615), .C1(new_n618), .C2(new_n556), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n571), .A2(new_n612), .A3(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n447), .A2(new_n493), .A3(new_n541), .A4(new_n620), .ZN(G372));
  NAND2_X1  g0421(.A1(new_n391), .A2(new_n393), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n411), .B1(new_n622), .B2(KEYINPUT17), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n353), .A2(new_n350), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n347), .B1(new_n280), .B2(G169), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n303), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n445), .B2(new_n307), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n410), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n343), .B1(new_n630), .B2(new_n340), .ZN(new_n631));
  INV_X1    g0431(.A(new_n447), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n601), .A2(new_n332), .ZN(new_n634));
  INV_X1    g0434(.A(new_n605), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n611), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n588), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n587), .B1(new_n586), .B2(new_n582), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n603), .A2(new_n400), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(G169), .B2(new_n603), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n636), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n633), .B1(new_n642), .B2(new_n619), .ZN(new_n643));
  INV_X1    g0443(.A(new_n570), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n615), .A2(new_n613), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n612), .A2(KEYINPUT26), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n589), .A2(new_n602), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n515), .A2(new_n522), .A3(new_n529), .A4(new_n531), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n650), .A2(new_n571), .A3(new_n612), .A4(new_n619), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n480), .A2(new_n483), .B1(new_n486), .B2(new_n489), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n515), .A2(new_n522), .ZN(new_n653));
  INV_X1    g0453(.A(new_n539), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n651), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n631), .B1(new_n632), .B2(new_n657), .ZN(G369));
  NAND2_X1  g0458(.A1(new_n484), .A2(new_n490), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n488), .A2(new_n666), .ZN(new_n667));
  MUX2_X1   g0467(.A(new_n493), .B(new_n659), .S(new_n667), .Z(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(G330), .ZN(new_n669));
  INV_X1    g0469(.A(new_n541), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n666), .B1(new_n515), .B2(new_n522), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n670), .A2(new_n671), .B1(new_n655), .B2(new_n666), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n673), .B(KEYINPUT82), .Z(new_n674));
  NAND2_X1  g0474(.A1(new_n659), .A2(new_n666), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n676), .A2(new_n541), .B1(new_n540), .B2(new_n666), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n674), .A2(new_n677), .ZN(G399));
  INV_X1    g0478(.A(new_n210), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G41), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n575), .A2(G116), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n219), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n657), .A2(KEYINPUT29), .A3(new_n665), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT31), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n666), .A2(new_n688), .ZN(new_n689));
  AND4_X1   g0489(.A1(G179), .A2(new_n460), .A3(new_n465), .A4(new_n467), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n603), .A2(new_n523), .A3(new_n528), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(new_n551), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n603), .A2(G179), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n481), .A2(new_n614), .A3(new_n530), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n698), .A2(KEYINPUT83), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n690), .A2(KEYINPUT30), .A3(new_n551), .A4(new_n692), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n698), .B2(KEYINPUT83), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n689), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(KEYINPUT84), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n487), .A2(new_n614), .A3(new_n691), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(KEYINPUT30), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n700), .B1(KEYINPUT84), .B2(new_n697), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n665), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n688), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n541), .A2(new_n493), .A3(new_n620), .A4(new_n666), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n702), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT85), .B1(new_n659), .B2(new_n540), .ZN(new_n713));
  AND4_X1   g0513(.A1(new_n650), .A2(new_n571), .A3(new_n612), .A4(new_n619), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT85), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n655), .A2(new_n715), .A3(new_n490), .A4(new_n484), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n649), .B1(new_n717), .B2(KEYINPUT86), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT86), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n713), .A2(new_n719), .A3(new_n714), .A4(new_n716), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n665), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n687), .B(new_n711), .C1(new_n712), .C2(new_n721), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT87), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n685), .B1(new_n724), .B2(G1), .ZN(G364));
  NOR2_X1   g0525(.A1(new_n295), .A2(G20), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n206), .B1(new_n726), .B2(G45), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n680), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n669), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(G330), .B2(new_n668), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n679), .A2(new_n360), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G355), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G116), .B2(new_n210), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n679), .A2(new_n327), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n271), .B2(new_n220), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n245), .A2(new_n271), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n216), .B1(G20), .B2(new_n402), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n729), .B1(new_n739), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(G20), .A2(G179), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n747), .A2(new_n384), .A3(G200), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n327), .B1(G322), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G311), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n747), .A2(G190), .A3(G200), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n749), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n384), .A2(G179), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n207), .ZN(new_n755));
  XOR2_X1   g0555(.A(KEYINPUT33), .B(G317), .Z(new_n756));
  INV_X1    g0556(.A(new_n747), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n384), .A3(G200), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n755), .A2(new_n526), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G303), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n207), .A2(new_n384), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n332), .A2(new_n400), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n760), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n207), .A2(G190), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n332), .A2(new_n400), .A3(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n207), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n767), .A2(G283), .B1(G329), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT90), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT88), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(KEYINPUT88), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT89), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n764), .B(new_n770), .C1(G326), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT91), .ZN(new_n778));
  INV_X1    g0578(.A(new_n748), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n327), .B1(new_n752), .B2(new_n285), .C1(new_n363), .C2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(G107), .B2(new_n767), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n768), .A2(G159), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT32), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n755), .A2(new_n555), .B1(new_n758), .B2(new_n283), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n763), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G87), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n774), .A2(G50), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n781), .A2(new_n785), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n777), .A2(KEYINPUT91), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n778), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n746), .B1(new_n791), .B2(new_n740), .ZN(new_n792));
  INV_X1    g0592(.A(new_n743), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n668), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n731), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(G396));
  NAND2_X1  g0596(.A1(new_n443), .A2(new_n665), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n440), .B1(new_n437), .B2(new_n438), .ZN(new_n798));
  AOI21_X1  g0598(.A(KEYINPUT68), .B1(new_n421), .B2(new_n432), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n445), .B(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT93), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n445), .A2(new_n666), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n441), .A2(KEYINPUT93), .A3(new_n445), .A4(new_n797), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n657), .B2(new_n665), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n802), .A2(new_n804), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n666), .B(new_n808), .C1(new_n649), .C2(new_n656), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n711), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n729), .B1(new_n810), .B2(new_n711), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n806), .A2(new_n741), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n740), .A2(new_n741), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n729), .B1(new_n816), .B2(G77), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G143), .A2(new_n748), .B1(new_n751), .B2(G159), .ZN(new_n818));
  INV_X1    g0618(.A(new_n774), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n818), .B1(new_n311), .B2(new_n758), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT34), .Z(new_n822));
  NOR2_X1   g0622(.A1(new_n766), .A2(new_n283), .ZN(new_n823));
  INV_X1    g0623(.A(new_n768), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n327), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n755), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n823), .B(new_n826), .C1(G58), .C2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n202), .B2(new_n763), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n766), .A2(new_n574), .B1(new_n824), .B2(new_n750), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT92), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n360), .B1(new_n779), .B2(new_n526), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G116), .B2(new_n751), .ZN(new_n833));
  INV_X1    g0633(.A(new_n758), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n827), .A2(G97), .B1(new_n834), .B2(G283), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n836), .B1(new_n496), .B2(new_n763), .C1(new_n761), .C2(new_n819), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n822), .A2(new_n829), .B1(new_n831), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n817), .B1(new_n838), .B2(new_n740), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n812), .A2(new_n813), .B1(new_n814), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G384));
  NOR2_X1   g0641(.A1(new_n726), .A2(new_n206), .ZN(new_n842));
  INV_X1    g0642(.A(G330), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  INV_X1    g0644(.A(new_n663), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n406), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n623), .B2(new_n629), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n406), .B1(new_n407), .B2(new_n845), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n390), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT37), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT37), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n848), .A2(new_n391), .A3(new_n851), .A4(new_n393), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n844), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n848), .A2(new_n391), .A3(new_n393), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n852), .ZN(new_n857));
  OAI211_X1 g0657(.A(KEYINPUT38), .B(new_n857), .C1(new_n412), .C2(new_n846), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n303), .B(new_n665), .C1(new_n354), .C2(new_n307), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n303), .A2(new_n665), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n626), .A2(new_n306), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n805), .A2(new_n863), .ZN(new_n864));
  AND4_X1   g0664(.A1(new_n481), .A2(new_n614), .A3(new_n530), .A4(new_n696), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT84), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n865), .A2(new_n866), .B1(new_n704), .B2(KEYINPUT30), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n693), .A2(new_n694), .B1(new_n697), .B2(KEYINPUT84), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n688), .B(new_n666), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n481), .A2(new_n696), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n870), .A2(new_n866), .A3(new_n530), .A4(new_n614), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n695), .A2(new_n871), .A3(new_n700), .A4(new_n703), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT31), .B1(new_n872), .B2(new_n665), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n864), .B1(new_n874), .B2(new_n709), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n859), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n872), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n709), .A2(new_n708), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n805), .A2(new_n863), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n857), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n844), .B1(new_n882), .B2(new_n847), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n858), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n876), .A2(KEYINPUT40), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n447), .A2(new_n878), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n843), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n887), .B2(new_n886), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT94), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n859), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n354), .A2(new_n303), .A3(new_n666), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n892), .B(new_n894), .C1(new_n891), .C2(new_n884), .ZN(new_n895));
  INV_X1    g0695(.A(new_n863), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n445), .A2(new_n665), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n809), .B2(new_n898), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n899), .A2(new_n884), .B1(new_n410), .B2(new_n663), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n631), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n687), .B1(new_n721), .B2(new_n712), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n904), .B2(new_n447), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n902), .B(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n842), .B1(new_n890), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n890), .B2(new_n906), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n567), .A2(KEYINPUT35), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n567), .A2(KEYINPUT35), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n909), .A2(G116), .A3(new_n217), .A4(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT36), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n219), .A2(new_n285), .A3(new_n364), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n283), .A2(G50), .ZN(new_n914));
  OAI211_X1 g0714(.A(G1), .B(new_n295), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n908), .A2(new_n912), .A3(new_n915), .ZN(G367));
  NAND2_X1  g0716(.A1(new_n676), .A2(new_n541), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n571), .B(new_n619), .C1(new_n570), .C2(new_n666), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n644), .A2(new_n645), .A3(new_n665), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT42), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n619), .B1(new_n918), .B2(new_n655), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n666), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT96), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT43), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT95), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n611), .A2(new_n666), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(new_n589), .A3(new_n602), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n929), .B(new_n931), .C1(new_n642), .C2(new_n930), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n931), .A2(new_n929), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n926), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n928), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n934), .B2(new_n928), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n674), .A2(new_n921), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n938), .B(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n727), .B(KEYINPUT98), .Z(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n677), .A2(new_n920), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT97), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT45), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n677), .A2(new_n920), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT44), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(new_n674), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n917), .B1(new_n672), .B2(new_n676), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n669), .B(new_n952), .Z(new_n953));
  NOR2_X1   g0753(.A1(new_n723), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n724), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n680), .B(KEYINPUT41), .Z(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n942), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n935), .A2(new_n793), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n744), .B1(new_n210), .B2(new_n414), .C1(new_n736), .C2(new_n236), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT99), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n729), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n775), .A2(G143), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n779), .A2(new_n311), .B1(new_n752), .B2(new_n202), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n327), .B1(new_n824), .B2(new_n820), .ZN(new_n968));
  INV_X1    g0768(.A(G159), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n755), .A2(new_n283), .B1(new_n758), .B2(new_n969), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G58), .A2(new_n786), .B1(new_n767), .B2(G77), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n966), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n775), .A2(G311), .B1(G303), .B2(new_n748), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT100), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n827), .A2(G107), .B1(new_n751), .B2(G283), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT46), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n763), .B2(new_n471), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n977), .B(new_n979), .C1(new_n526), .C2(new_n758), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT102), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n327), .B1(new_n768), .B2(G317), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n555), .B2(new_n766), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n980), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n763), .A2(new_n978), .A3(new_n471), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n983), .A2(new_n981), .B1(new_n985), .B2(KEYINPUT101), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(KEYINPUT101), .B2(new_n985), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n976), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n974), .A2(new_n975), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n973), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT47), .Z(new_n991));
  INV_X1    g0791(.A(new_n740), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n965), .B1(new_n962), .B2(new_n961), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n940), .A2(new_n959), .B1(new_n960), .B2(new_n993), .ZN(G387));
  XOR2_X1   g0794(.A(new_n680), .B(KEYINPUT105), .Z(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n954), .A2(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n997), .A2(KEYINPUT106), .B1(new_n723), .B2(new_n953), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(KEYINPUT106), .B2(new_n997), .ZN(new_n999));
  INV_X1    g0799(.A(new_n682), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n732), .A2(new_n1000), .B1(new_n496), .B2(new_n679), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n241), .A2(new_n271), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n310), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n202), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT50), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n682), .B(new_n271), .C1(new_n283), .C2(new_n285), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n735), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1001), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n744), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n729), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n672), .A2(new_n793), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n768), .A2(G150), .B1(new_n751), .B2(G68), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1012), .B(new_n327), .C1(new_n202), .C2(new_n779), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n755), .A2(new_n414), .B1(new_n758), .B2(new_n310), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n285), .A2(new_n763), .B1(new_n766), .B2(new_n555), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n969), .B2(new_n819), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT103), .Z(new_n1018));
  XNOR2_X1  g0818(.A(KEYINPUT104), .B(G322), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n775), .A2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G303), .A2(new_n751), .B1(new_n748), .B2(G317), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(new_n750), .C2(new_n758), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(G283), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n763), .A2(new_n526), .B1(new_n755), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(KEYINPUT49), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n327), .B1(new_n768), .B2(G326), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(new_n471), .C2(new_n766), .ZN(new_n1030));
  AOI21_X1  g0830(.A(KEYINPUT49), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1018), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1010), .B(new_n1011), .C1(new_n1032), .C2(new_n740), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n953), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1033), .B1(new_n1034), .B2(new_n942), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n999), .A2(new_n1035), .ZN(G393));
  AOI21_X1  g0836(.A(new_n996), .B1(new_n951), .B2(new_n954), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n954), .B2(new_n951), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n951), .A2(new_n942), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n736), .A2(new_n248), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n744), .B1(new_n555), .B2(new_n210), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n729), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n827), .A2(G116), .B1(new_n751), .B2(G294), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n761), .B2(new_n758), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT107), .Z(new_n1045));
  NAND2_X1  g0845(.A1(new_n767), .A2(G107), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n786), .A2(G283), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n327), .B1(new_n768), .B2(new_n1019), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n774), .A2(G317), .B1(G311), .B2(new_n748), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT52), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n774), .A2(G150), .B1(G159), .B2(new_n748), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n768), .A2(G143), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1054), .B(new_n327), .C1(new_n310), .C2(new_n752), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n755), .A2(new_n285), .B1(new_n758), .B2(new_n202), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n283), .B2(new_n763), .C1(new_n574), .C2(new_n766), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1049), .A2(new_n1051), .B1(new_n1053), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1042), .B1(new_n1059), .B2(new_n740), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n920), .B2(new_n793), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1038), .A2(new_n1039), .A3(new_n1061), .ZN(G390));
  AND3_X1   g0862(.A1(new_n883), .A2(KEYINPUT39), .A3(new_n858), .ZN(new_n1063));
  AOI21_X1  g0863(.A(KEYINPUT39), .B1(new_n854), .B2(new_n858), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n741), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n729), .B1(new_n816), .B2(new_n1003), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n824), .A2(new_n526), .B1(new_n752), .B2(new_n555), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n327), .B(new_n1067), .C1(G116), .C2(new_n748), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n774), .A2(G283), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n827), .A2(G77), .B1(new_n834), .B2(G107), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n823), .B1(G87), .B2(new_n786), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n774), .A2(G128), .B1(G132), .B2(new_n748), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT109), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n763), .A2(new_n311), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT53), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n360), .B1(new_n768), .B2(G125), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(KEYINPUT54), .B(G143), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n752), .B2(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n755), .A2(new_n969), .B1(new_n758), .B2(new_n820), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1076), .B(new_n1081), .C1(new_n202), .C2(new_n766), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1072), .B1(new_n1074), .B2(new_n1082), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1083), .A2(KEYINPUT110), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n992), .B1(new_n1083), .B2(KEYINPUT110), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1066), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1065), .A2(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1063), .A2(new_n1064), .B1(new_n899), .B2(new_n894), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n714), .A2(new_n716), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n715), .B1(new_n652), .B2(new_n655), .ZN(new_n1090));
  OAI21_X1  g0890(.A(KEYINPUT86), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n649), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n1092), .A3(new_n720), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1093), .A2(new_n666), .A3(new_n808), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n896), .B1(new_n1094), .B2(new_n898), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n859), .A2(new_n893), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1088), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n843), .B1(new_n874), .B2(new_n709), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n879), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n710), .A2(G330), .A3(new_n805), .A4(new_n863), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1088), .B(new_n1102), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1087), .B1(new_n1104), .B2(new_n941), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n897), .B1(new_n721), .B2(new_n808), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n859), .B(new_n893), .C1(new_n1106), .C2(new_n896), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1099), .B1(new_n1107), .B2(new_n1088), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1103), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n447), .A2(new_n1098), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n905), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n896), .B1(new_n711), .B2(new_n806), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1099), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n809), .A2(new_n898), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n878), .A2(G330), .A3(new_n805), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n896), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1117), .A2(new_n1102), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1114), .A2(new_n1115), .B1(new_n1118), .B2(new_n1106), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT108), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n996), .B1(new_n1110), .B2(new_n1120), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n905), .A2(new_n1111), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1118), .A2(new_n1106), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1126), .A2(KEYINPUT108), .A3(new_n1104), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1105), .B1(new_n1121), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(G378));
  NAND2_X1  g0929(.A1(new_n360), .A2(new_n270), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1130), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT111), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n767), .A2(G58), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1130), .B1(G283), .B2(new_n768), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(new_n285), .C2(new_n763), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT112), .Z(new_n1136));
  NOR2_X1   g0936(.A1(new_n819), .A2(new_n471), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n581), .A2(new_n751), .B1(new_n748), .B2(G107), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n283), .B2(new_n755), .C1(new_n555), .C2(new_n758), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1132), .B1(new_n1140), .B2(KEYINPUT58), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT113), .Z(new_n1142));
  NOR2_X1   g0942(.A1(new_n763), .A2(new_n1078), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G128), .A2(new_n748), .B1(new_n751), .B2(G137), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n825), .B2(new_n758), .C1(new_n311), .C2(new_n755), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(G125), .C2(new_n774), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT114), .Z(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  AOI211_X1 g0948(.A(G33), .B(G41), .C1(new_n768), .C2(G124), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n969), .B2(new_n766), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n1147), .B2(KEYINPUT59), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1148), .A2(new_n1151), .B1(KEYINPUT58), .B2(new_n1140), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1142), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n992), .B1(new_n1153), .B2(KEYINPUT115), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(KEYINPUT115), .B2(new_n1153), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n729), .C1(G50), .C2(new_n816), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT116), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n316), .A2(new_n845), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n340), .B2(new_n344), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n340), .A2(new_n344), .A3(new_n1159), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1158), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1159), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1164), .B(new_n343), .C1(new_n336), .C2(new_n339), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1158), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1160), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1157), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1161), .A2(new_n1162), .A3(new_n1158), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1166), .B1(new_n1160), .B2(new_n1165), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n1170), .A3(KEYINPUT116), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1172), .A2(new_n742), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1156), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n885), .B2(new_n843), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n881), .A2(new_n884), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n880), .B1(new_n859), .B2(new_n875), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1172), .B(G330), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1176), .A2(new_n901), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n901), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1174), .B1(new_n1182), .B2(new_n942), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1180), .A2(new_n1181), .A3(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1101), .A2(new_n1125), .A3(new_n1103), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n1122), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1186), .A2(KEYINPUT117), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT117), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1188), .A2(new_n1182), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n996), .B1(new_n1192), .B2(new_n1185), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1184), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(G375));
  NAND2_X1  g0995(.A1(new_n896), .A2(new_n741), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n729), .B1(new_n816), .B2(G68), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT118), .Z(new_n1198));
  NAND2_X1  g0998(.A1(new_n774), .A2(G132), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT119), .Z(new_n1200));
  OAI22_X1  g1000(.A1(new_n779), .A2(new_n820), .B1(new_n752), .B2(new_n311), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n360), .B(new_n1201), .C1(G128), .C2(new_n768), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1078), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n827), .A2(G50), .B1(new_n834), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n786), .A2(G159), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1202), .A2(new_n1133), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n819), .A2(new_n526), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G77), .A2(new_n767), .B1(new_n786), .B2(G97), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n327), .B1(G283), .B2(new_n748), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n768), .A2(G303), .B1(new_n751), .B2(G107), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n827), .A2(new_n581), .B1(new_n834), .B2(G116), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1200), .A2(new_n1206), .B1(new_n1207), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1198), .B1(new_n1213), .B2(new_n740), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1125), .A2(new_n942), .B1(new_n1196), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1126), .A2(new_n958), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(G381));
  INV_X1    g1018(.A(G387), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n999), .A2(new_n795), .A3(new_n1035), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(G390), .A2(G378), .A3(G384), .A4(G381), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(new_n1221), .A3(new_n1194), .A4(new_n1222), .ZN(G407));
  NAND2_X1  g1023(.A1(new_n664), .A2(G213), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1194), .A2(new_n1128), .A3(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(G407), .A2(G213), .A3(new_n1226), .ZN(G409));
  INV_X1    g1027(.A(G390), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G387), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT122), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G393), .A2(G396), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1220), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(G387), .B(new_n1228), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1233), .B(new_n1234), .Z(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(KEYINPUT61), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT63), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1188), .A2(new_n1182), .A3(new_n958), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1183), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1128), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT120), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n1128), .A3(KEYINPUT120), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1194), .A2(G378), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(KEYINPUT121), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1190), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1186), .A2(KEYINPUT117), .A3(new_n1188), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1193), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(G378), .A3(new_n1183), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1246), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT121), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1245), .A2(new_n1253), .A3(new_n1224), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1217), .A2(KEYINPUT60), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1217), .A2(KEYINPUT60), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1256), .A2(new_n995), .A3(new_n1126), .A4(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1215), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n840), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(G384), .A3(new_n1215), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1237), .B1(new_n1255), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT123), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1244), .B2(new_n1225), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1251), .A2(KEYINPUT123), .A3(new_n1224), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1262), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1225), .A2(G2897), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1262), .A2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1260), .A2(G2897), .A3(new_n1225), .A4(new_n1261), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1255), .A2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1236), .A2(new_n1263), .A3(new_n1268), .A4(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1225), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1262), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .A4(new_n1245), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n1267), .B2(new_n1276), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1265), .A2(new_n1266), .A3(new_n1272), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT125), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT125), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1280), .A2(new_n1284), .A3(new_n1281), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1279), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1235), .B1(new_n1286), .B2(KEYINPUT126), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1288), .B(new_n1279), .C1(new_n1283), .C2(new_n1285), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1274), .B1(new_n1287), .B2(new_n1289), .ZN(G405));
  NAND2_X1  g1090(.A1(G375), .A2(new_n1128), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1250), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(new_n1262), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT127), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1293), .B1(new_n1235), .B2(new_n1294), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1233), .B(new_n1234), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT127), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1295), .B(new_n1297), .ZN(G402));
endmodule


