//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G128), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT64), .A3(G146), .ZN(new_n196));
  AOI22_X1  g010(.A1(new_n194), .A2(new_n196), .B1(G143), .B2(new_n193), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(G143), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT67), .B1(new_n197), .B2(new_n200), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n195), .A2(KEYINPUT64), .A3(G146), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT64), .B1(new_n195), .B2(G146), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n199), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT1), .B1(new_n195), .B2(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n191), .B1(new_n201), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G134), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G137), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n212), .B2(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n213), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n215), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n209), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT0), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(new_n198), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n204), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n195), .A2(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n199), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT11), .B1(new_n210), .B2(G134), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n210), .A2(G134), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n238), .A2(new_n239), .A3(new_n219), .A4(new_n218), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n217), .A2(new_n218), .A3(new_n213), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n219), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n238), .A2(KEYINPUT66), .A3(new_n218), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n235), .B1(new_n242), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n187), .B1(new_n224), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT2), .B(G113), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G116), .B(G119), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(KEYINPUT68), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n254));
  INV_X1    g068(.A(G119), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G116), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G119), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n254), .B1(new_n259), .B2(new_n250), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n250), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n197), .A2(KEYINPUT67), .A3(new_n200), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n205), .B1(new_n204), .B2(new_n207), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n190), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n240), .A2(new_n241), .B1(G131), .B2(new_n214), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n247), .A2(new_n242), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n230), .A2(new_n234), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n271), .A3(KEYINPUT30), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n249), .A2(new_n263), .A3(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(KEYINPUT26), .B(G101), .Z(new_n274));
  NOR2_X1   g088(.A1(G237), .A2(G953), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G210), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n274), .B(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n263), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n268), .A2(new_n271), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n273), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT31), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n263), .B1(new_n224), .B2(new_n248), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n268), .A2(new_n271), .A3(KEYINPUT28), .A4(new_n281), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n279), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n273), .A2(new_n291), .A3(new_n280), .A4(new_n282), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n284), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n284), .A2(new_n295), .A3(new_n290), .A4(new_n292), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT32), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n297), .A2(KEYINPUT32), .A3(new_n298), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n287), .A2(KEYINPUT71), .A3(new_n282), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n304), .B(new_n263), .C1(new_n224), .C2(new_n248), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(KEYINPUT28), .A3(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n306), .A2(KEYINPUT29), .A3(new_n280), .A4(new_n286), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT72), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n307), .A2(new_n311), .A3(new_n308), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n273), .A2(new_n282), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n279), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n289), .A2(new_n280), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT29), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G472), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n301), .A2(new_n302), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G217), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(G234), .B2(new_n308), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n255), .A2(G128), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT23), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT74), .B(G110), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n198), .A2(G119), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n324), .B(new_n325), .C1(new_n328), .C2(new_n323), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n330), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n323), .A2(new_n326), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT24), .B(G110), .Z(new_n334));
  OAI211_X1 g148(.A(new_n331), .B(new_n332), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(G125), .ZN(new_n339));
  INV_X1    g153(.A(G125), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G140), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(G146), .B(new_n338), .C1(new_n342), .C2(new_n336), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n344));
  AND4_X1   g158(.A1(new_n344), .A2(new_n339), .A3(new_n341), .A4(new_n193), .ZN(new_n345));
  XNOR2_X1  g159(.A(G125), .B(G140), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n346), .B2(new_n193), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n335), .B(new_n343), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G110), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n324), .B1(new_n328), .B2(new_n323), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(new_n350), .B2(KEYINPUT73), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(KEYINPUT73), .B2(new_n350), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n338), .B1(new_n342), .B2(new_n336), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n193), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n343), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n333), .A2(new_n334), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n348), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT22), .B(G137), .ZN(new_n359));
  INV_X1    g173(.A(G221), .ZN(new_n360));
  INV_X1    g174(.A(G234), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n360), .A2(new_n361), .A3(G953), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n359), .B(new_n362), .Z(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n363), .B1(new_n348), .B2(new_n357), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT25), .B1(new_n367), .B2(new_n308), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT25), .ZN(new_n369));
  NOR4_X1   g183(.A1(new_n365), .A2(new_n366), .A3(new_n369), .A4(G902), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n322), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n367), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n322), .A2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n371), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G469), .ZN(new_n377));
  XNOR2_X1  g191(.A(G110), .B(G140), .ZN(new_n378));
  INV_X1    g192(.A(G953), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G227), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n378), .B(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(new_n382), .B2(G107), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G104), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(G107), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT77), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n383), .A2(new_n386), .A3(KEYINPUT77), .A4(new_n387), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(G101), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G101), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n383), .A2(new_n386), .A3(new_n393), .A4(new_n387), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n390), .A2(new_n397), .A3(G101), .A4(new_n391), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n270), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n382), .A2(G107), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n385), .A2(G104), .ZN(new_n401));
  OAI21_X1  g215(.A(G101), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n266), .A2(KEYINPUT10), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT78), .B1(new_n200), .B2(new_n188), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT78), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n207), .A2(new_n407), .A3(new_n232), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n190), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT10), .B1(new_n409), .B2(new_n404), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT79), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI211_X1 g226(.A(KEYINPUT79), .B(KEYINPUT10), .C1(new_n409), .C2(new_n404), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n399), .B(new_n405), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n381), .B1(new_n414), .B2(new_n269), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n409), .A2(new_n404), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n266), .B2(new_n404), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n417), .A2(KEYINPUT12), .A3(new_n269), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT12), .B1(new_n417), .B2(new_n269), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n410), .B(new_n411), .ZN(new_n422));
  INV_X1    g236(.A(new_n269), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n399), .A4(new_n405), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n414), .A2(new_n269), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n381), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n377), .B(new_n308), .C1(new_n421), .C2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n377), .A2(new_n308), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n381), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n414), .A2(new_n269), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n430), .B1(new_n420), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n424), .A2(new_n425), .A3(new_n381), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n427), .B(new_n429), .C1(new_n434), .C2(new_n377), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT9), .B(G234), .Z(new_n436));
  AOI21_X1  g250(.A(new_n360), .B1(new_n436), .B2(new_n308), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G128), .B(G143), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n212), .B1(new_n440), .B2(KEYINPUT13), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n195), .A2(G128), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n441), .B1(KEYINPUT13), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n212), .ZN(new_n444));
  INV_X1    g258(.A(G122), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G116), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n257), .A2(G122), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT94), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT94), .B1(new_n446), .B2(new_n447), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n448), .A2(new_n449), .A3(G107), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT94), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n257), .A2(G122), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n445), .A2(G116), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT94), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n385), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n443), .B(new_n444), .C1(new_n450), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT95), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n440), .B(new_n212), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n454), .A2(new_n385), .A3(new_n455), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n385), .B1(new_n453), .B2(KEYINPUT14), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n446), .A2(new_n447), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n461), .B1(KEYINPUT14), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G107), .B1(new_n448), .B2(new_n449), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n460), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT95), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n466), .A2(new_n467), .A3(new_n444), .A4(new_n443), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n458), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n436), .A2(G217), .A3(new_n379), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT96), .ZN(new_n472));
  INV_X1    g286(.A(new_n470), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n458), .A2(new_n464), .A3(new_n468), .A4(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n469), .A2(KEYINPUT96), .A3(new_n470), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n308), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT15), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(G478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(G478), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n475), .A2(new_n308), .A3(new_n480), .A4(new_n476), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT92), .ZN(new_n484));
  INV_X1    g298(.A(G237), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n379), .A3(G214), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n195), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n275), .A2(G143), .A3(G214), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT18), .A4(G131), .ZN(new_n491));
  OAI22_X1  g305(.A1(new_n347), .A2(new_n345), .B1(new_n193), .B2(new_n346), .ZN(new_n492));
  NAND2_X1  g306(.A1(KEYINPUT18), .A2(G131), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n486), .A2(new_n195), .ZN(new_n494));
  AOI21_X1  g308(.A(G143), .B1(new_n275), .B2(G214), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n493), .B1(new_n496), .B2(KEYINPUT87), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(KEYINPUT87), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n491), .B(new_n492), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT90), .B(G104), .Z(new_n500));
  XNOR2_X1  g314(.A(G113), .B(G122), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G131), .B1(new_n494), .B2(new_n495), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n487), .A2(new_n219), .A3(new_n488), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n489), .A2(KEYINPUT17), .A3(G131), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n506), .A2(new_n343), .A3(new_n354), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n499), .A2(new_n502), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT91), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n499), .A2(new_n508), .A3(new_n511), .A4(new_n502), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n503), .A2(new_n505), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT88), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT88), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n503), .A2(new_n516), .A3(new_n505), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n343), .A3(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n346), .A2(KEYINPUT89), .A3(KEYINPUT19), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT19), .B1(new_n346), .B2(KEYINPUT89), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(G146), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n499), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n502), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n484), .B1(new_n513), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n510), .A2(new_n512), .B1(new_n523), .B2(new_n524), .ZN(new_n527));
  NOR2_X1   g341(.A1(G475), .A2(G902), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OAI22_X1  g343(.A1(new_n526), .A2(KEYINPUT20), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n513), .A2(new_n525), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT20), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n531), .A2(new_n484), .A3(new_n532), .A4(new_n528), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n510), .A2(new_n512), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n502), .B1(new_n499), .B2(new_n508), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n308), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT93), .B(G475), .Z(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n530), .A2(new_n533), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(G902), .B(G953), .C1(new_n361), .C2(new_n485), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n540), .B(KEYINPUT97), .Z(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT21), .B(G898), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n379), .A2(G952), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n361), .B2(new_n485), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n483), .A2(new_n539), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(G210), .B1(G237), .B2(G902), .ZN(new_n548));
  XOR2_X1   g362(.A(new_n548), .B(KEYINPUT86), .Z(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT5), .ZN(new_n551));
  OR3_X1    g365(.A1(new_n257), .A2(KEYINPUT5), .A3(G119), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(G113), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT80), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT80), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n551), .A2(new_n552), .A3(new_n555), .A4(G113), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n554), .A2(new_n556), .B1(new_n260), .B2(new_n253), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT85), .B1(new_n557), .B2(new_n404), .ZN(new_n558));
  INV_X1    g372(.A(G113), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(new_n252), .B2(KEYINPUT5), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n555), .B1(new_n560), .B2(new_n552), .ZN(new_n561));
  INV_X1    g375(.A(new_n556), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n261), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT85), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n403), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n261), .A2(new_n404), .A3(new_n553), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n558), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(G110), .B(G122), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT81), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g384(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n396), .A2(new_n263), .A3(new_n398), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n261), .B(new_n404), .C1(new_n561), .C2(new_n562), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT83), .B1(new_n270), .B2(new_n340), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n209), .A2(new_n340), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT83), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n235), .A2(new_n579), .A3(G125), .ZN(new_n580));
  INV_X1    g394(.A(G224), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(G953), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT7), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n577), .A2(new_n578), .A3(new_n580), .A4(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n578), .B1(new_n340), .B2(new_n270), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n584), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n573), .A2(new_n576), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n308), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n574), .A2(new_n570), .A3(new_n575), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT82), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n570), .B(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n574), .B2(new_n575), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT6), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n574), .A2(new_n575), .ZN(new_n596));
  INV_X1    g410(.A(new_n593), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT6), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n582), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n577), .A2(new_n578), .A3(new_n583), .A4(new_n580), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n595), .A2(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n550), .B1(new_n590), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(G214), .B1(G237), .B2(G902), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n603), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n599), .B1(new_n598), .B2(new_n576), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n594), .A2(KEYINPUT6), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n610), .A2(new_n308), .A3(new_n549), .A4(new_n589), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n605), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n439), .A2(new_n547), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n320), .A2(new_n376), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  AOI21_X1  g429(.A(G902), .B1(new_n294), .B2(new_n296), .ZN(new_n616));
  INV_X1    g430(.A(G472), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n299), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n439), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n376), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT98), .B1(new_n469), .B2(new_n470), .ZN(new_n623));
  INV_X1    g437(.A(new_n474), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT33), .B1(new_n474), .B2(KEYINPUT98), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT99), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n626), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n628), .B(new_n629), .C1(new_n624), .C2(new_n623), .ZN(new_n630));
  INV_X1    g444(.A(G478), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(G902), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n475), .A2(new_n633), .A3(new_n476), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n627), .A2(new_n630), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n477), .A2(new_n631), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n530), .A2(new_n533), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n536), .A2(new_n538), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n605), .A2(new_n611), .A3(new_n606), .A4(new_n546), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n622), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n636), .A2(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n644));
  INV_X1    g458(.A(new_n612), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n644), .A2(KEYINPUT100), .A3(new_n645), .A4(new_n546), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n621), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT34), .B(G104), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  NAND3_X1  g463(.A1(new_n531), .A2(new_n532), .A3(new_n528), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT20), .B1(new_n527), .B2(new_n529), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n650), .A2(new_n651), .B1(new_n536), .B2(new_n538), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n546), .B(KEYINPUT101), .Z(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n482), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n482), .A2(new_n652), .A3(KEYINPUT102), .A4(new_n654), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n657), .A2(new_n645), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n621), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT35), .B(G107), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  NOR2_X1   g477(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n358), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n373), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n371), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n619), .A2(new_n613), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT37), .B(G110), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G12));
  AOI21_X1  g484(.A(new_n612), .B1(new_n371), .B2(new_n666), .ZN(new_n671));
  INV_X1    g485(.A(new_n545), .ZN(new_n672));
  INV_X1    g486(.A(G900), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n672), .B1(new_n541), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n482), .A2(new_n652), .A3(new_n675), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n320), .A2(new_n620), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  NAND2_X1  g493(.A1(new_n640), .A2(new_n482), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n674), .B(KEYINPUT39), .Z(new_n682));
  NAND2_X1  g496(.A1(new_n620), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n681), .B1(new_n683), .B2(KEYINPUT40), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(KEYINPUT40), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n314), .A2(new_n280), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n303), .A2(new_n305), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n686), .B1(new_n687), .B2(new_n280), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT103), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n686), .B(new_n690), .C1(new_n280), .C2(new_n687), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n308), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G472), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n301), .A2(new_n302), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n605), .A2(new_n611), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT38), .ZN(new_n696));
  INV_X1    g510(.A(new_n606), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n696), .A2(new_n697), .A3(new_n667), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n685), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G143), .ZN(G45));
  NAND2_X1  g514(.A1(new_n644), .A2(new_n675), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n320), .A2(new_n620), .A3(new_n671), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  NAND2_X1  g518(.A1(new_n643), .A2(new_n646), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n308), .B1(new_n421), .B2(new_n426), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n438), .A3(new_n427), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n707), .A2(KEYINPUT104), .A3(new_n438), .A4(new_n427), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n705), .A2(new_n320), .A3(new_n712), .A4(new_n376), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n320), .A2(new_n712), .A3(new_n376), .A4(new_n659), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT105), .B(G116), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G18));
  AND3_X1   g532(.A1(new_n710), .A2(new_n671), .A3(new_n711), .ZN(new_n719));
  INV_X1    g533(.A(new_n547), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n320), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  NAND2_X1  g536(.A1(new_n297), .A2(new_n308), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT107), .B(G472), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n280), .B1(new_n306), .B2(new_n286), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n284), .ZN(new_n728));
  INV_X1    g542(.A(new_n284), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT106), .B1(new_n729), .B2(new_n725), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n728), .A2(new_n730), .A3(new_n292), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n723), .A2(new_n724), .B1(new_n731), .B2(new_n298), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n680), .A2(new_n612), .A3(new_n653), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n712), .A2(new_n376), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT108), .B(G122), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G24));
  NAND3_X1  g550(.A1(new_n719), .A2(new_n702), .A3(new_n732), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  AOI21_X1  g552(.A(KEYINPUT32), .B1(new_n297), .B2(new_n298), .ZN(new_n739));
  INV_X1    g553(.A(new_n298), .ZN(new_n740));
  AOI211_X1 g554(.A(new_n300), .B(new_n740), .C1(new_n294), .C2(new_n296), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n375), .B1(new_n742), .B2(new_n319), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT109), .B1(new_n695), .B2(new_n606), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n745));
  AOI211_X1 g559(.A(new_n745), .B(new_n697), .C1(new_n605), .C2(new_n611), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n439), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n743), .A2(KEYINPUT42), .A3(new_n702), .A4(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n320), .A2(new_n376), .A3(new_n702), .A4(new_n747), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  AND4_X1   g567(.A1(new_n320), .A2(new_n676), .A3(new_n376), .A4(new_n747), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n212), .ZN(G36));
  INV_X1    g569(.A(new_n427), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n434), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n432), .A2(KEYINPUT45), .A3(new_n433), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(G469), .A3(new_n759), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n428), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n756), .B1(new_n763), .B2(KEYINPUT46), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(KEYINPUT46), .B2(new_n763), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n438), .A3(new_n682), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n744), .A2(new_n746), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n637), .A2(new_n539), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT43), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n618), .A3(new_n667), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n767), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n766), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n210), .ZN(G39));
  NAND2_X1  g590(.A1(new_n765), .A2(new_n438), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT47), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT47), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n765), .A2(new_n779), .A3(new_n438), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n701), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n320), .A2(new_n376), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n767), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  XNOR2_X1  g599(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n781), .A2(KEYINPUT112), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n778), .A2(new_n788), .A3(new_n780), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n707), .A2(new_n437), .A3(new_n427), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n770), .A2(new_n672), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n732), .A2(new_n376), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n767), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n794), .A2(new_n697), .A3(new_n696), .A4(new_n712), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n732), .A2(new_n667), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n712), .A2(new_n767), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n545), .B1(new_n805), .B2(KEYINPUT113), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n712), .A2(new_n767), .A3(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n810), .A3(new_n770), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n806), .A2(new_n770), .A3(new_n808), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT114), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n804), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n637), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n694), .A2(new_n375), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n539), .A2(new_n809), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n803), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n786), .B1(new_n797), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n814), .ZN(new_n820));
  INV_X1    g634(.A(new_n817), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(KEYINPUT51), .A3(new_n802), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n795), .B1(new_n781), .B2(new_n790), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n544), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n809), .A2(new_n816), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n644), .ZN(new_n827));
  INV_X1    g641(.A(new_n712), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n792), .A2(new_n828), .A3(new_n793), .A4(new_n612), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT115), .Z(new_n830));
  NOR2_X1   g644(.A1(new_n439), .A2(new_n612), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n667), .A2(new_n674), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n694), .A2(new_n831), .A3(new_n681), .A4(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n703), .A2(new_n833), .A3(new_n737), .A4(new_n678), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n834), .B(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n667), .ZN(new_n837));
  INV_X1    g651(.A(new_n747), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n652), .A2(new_n675), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n320), .A2(new_n483), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n732), .A2(new_n702), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n837), .B(new_n838), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n713), .A2(new_n716), .A3(new_n721), .A4(new_n734), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n539), .A2(new_n482), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n612), .B(new_n653), .C1(new_n641), .C2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n619), .A3(new_n376), .A4(new_n620), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n614), .A3(new_n668), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n843), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n754), .B1(new_n748), .B2(new_n751), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n836), .A2(KEYINPUT53), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n841), .A2(new_n842), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n667), .A3(new_n747), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n713), .A2(new_n716), .A3(new_n721), .A4(new_n734), .ZN(new_n855));
  INV_X1    g669(.A(new_n848), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n850), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n439), .B1(new_n742), .B2(new_n319), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n731), .A2(new_n298), .ZN(new_n860));
  INV_X1    g674(.A(new_n724), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n616), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n860), .A2(new_n862), .A3(new_n701), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n859), .A2(new_n677), .B1(new_n863), .B2(new_n719), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n835), .A3(new_n703), .A4(new_n833), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n858), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n852), .B1(new_n857), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n851), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT54), .Z(new_n869));
  NAND4_X1  g683(.A1(new_n825), .A2(new_n827), .A3(new_n830), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n743), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n811), .B2(new_n813), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT48), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n870), .A2(new_n873), .B1(G952), .B2(G953), .ZN(new_n874));
  INV_X1    g688(.A(new_n696), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n707), .A2(new_n427), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n376), .B1(new_n876), .B2(KEYINPUT49), .ZN(new_n877));
  AOI211_X1 g691(.A(new_n875), .B(new_n877), .C1(KEYINPUT49), .C2(new_n876), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n768), .A2(new_n697), .A3(new_n437), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n742), .A3(new_n693), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n874), .A2(new_n880), .ZN(G75));
  NAND2_X1  g695(.A1(new_n595), .A2(new_n600), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT116), .Z(new_n883));
  AOI21_X1  g697(.A(new_n308), .B1(new_n851), .B2(new_n867), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n549), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n886), .A3(new_n883), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n607), .B(KEYINPUT55), .Z(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n888), .B2(new_n889), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n379), .A2(G952), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(G51));
  XNOR2_X1  g709(.A(new_n868), .B(KEYINPUT54), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT57), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n428), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n429), .A2(KEYINPUT57), .ZN(new_n899));
  OAI22_X1  g713(.A1(new_n898), .A2(new_n899), .B1(new_n426), .B2(new_n421), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n884), .A2(new_n761), .A3(new_n762), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n894), .B1(new_n900), .B2(new_n901), .ZN(G54));
  NAND2_X1  g716(.A1(KEYINPUT58), .A2(G475), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT117), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n903), .A2(KEYINPUT117), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n884), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n527), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n894), .ZN(G60));
  AND3_X1   g722(.A1(new_n627), .A2(new_n630), .A3(new_n634), .ZN(new_n909));
  NAND2_X1  g723(.A1(G478), .A2(G902), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT59), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n896), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n894), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n912), .A2(KEYINPUT118), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT118), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n909), .B1(new_n896), .B2(new_n911), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(G63));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n321), .A2(new_n308), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n868), .A2(new_n665), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT61), .ZN(new_n923));
  INV_X1    g737(.A(new_n921), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n851), .B2(new_n867), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n913), .B1(new_n925), .B2(new_n367), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n918), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT61), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n925), .B2(new_n665), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n844), .A2(new_n848), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n930), .A2(new_n854), .A3(new_n850), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT53), .B1(new_n931), .B2(new_n836), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n857), .A2(new_n866), .A3(new_n852), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n921), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n372), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n929), .A2(new_n935), .A3(KEYINPUT121), .A4(new_n913), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n927), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n868), .A2(KEYINPUT120), .A3(new_n665), .A4(new_n921), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n938), .B(new_n913), .C1(new_n367), .C2(new_n925), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT120), .B1(new_n925), .B2(new_n665), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n928), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n937), .A2(new_n941), .A3(KEYINPUT122), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(G66));
  OAI21_X1  g760(.A(G953), .B1(new_n542), .B2(new_n581), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n930), .B2(G953), .ZN(new_n948));
  INV_X1    g762(.A(new_n883), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(G898), .B2(new_n379), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  NOR2_X1   g765(.A1(new_n871), .A2(new_n838), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n641), .A2(new_n845), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n953), .A2(new_n682), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n775), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n699), .A2(new_n703), .A3(new_n864), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(KEYINPUT124), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n957), .A2(KEYINPUT124), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n956), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n784), .A2(new_n955), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n962), .A2(new_n379), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n249), .A2(new_n272), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(new_n521), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT123), .ZN(new_n966));
  NOR4_X1   g780(.A1(new_n766), .A2(new_n871), .A3(new_n612), .A4(new_n680), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n864), .A2(new_n703), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n967), .A2(new_n775), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n784), .A2(new_n850), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n965), .B1(new_n970), .B2(G953), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n673), .A2(new_n379), .ZN(new_n972));
  OAI22_X1  g786(.A1(new_n963), .A2(new_n966), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n379), .B1(G227), .B2(G900), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(G72));
  XNOR2_X1  g789(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n617), .A2(new_n308), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n976), .B(new_n977), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n930), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n979), .B1(new_n962), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n686), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n981), .A2(KEYINPUT126), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(KEYINPUT126), .B1(new_n981), .B2(new_n982), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n979), .B1(new_n970), .B2(new_n980), .ZN(new_n986));
  INV_X1    g800(.A(new_n316), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n894), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n982), .B1(new_n851), .B2(new_n867), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n987), .A2(new_n978), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n989), .A2(KEYINPUT127), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(KEYINPUT127), .B1(new_n989), .B2(new_n990), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n985), .A2(new_n993), .ZN(G57));
endmodule


