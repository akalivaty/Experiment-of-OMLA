//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT76), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G137), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT66), .A2(G134), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT66), .A2(G134), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(G137), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n197), .A2(G131), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n199), .A2(new_n200), .ZN(new_n204));
  INV_X1    g018(.A(new_n196), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n198), .A2(KEYINPUT11), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT66), .A2(G134), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n203), .B1(new_n204), .B2(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n202), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G104), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n212), .A2(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G101), .ZN(new_n219));
  INV_X1    g033(.A(G101), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n213), .A2(new_n216), .A3(new_n220), .A4(new_n217), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G143), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G146), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n223), .A2(KEYINPUT65), .A3(G143), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n225), .B2(G146), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n225), .A2(G146), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT0), .ZN(new_n234));
  INV_X1    g048(.A(G128), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT64), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(KEYINPUT0), .B2(G128), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n227), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n228), .B1(new_n233), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n218), .A2(new_n241), .A3(G101), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n222), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n212), .A2(G107), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n215), .A2(G104), .ZN(new_n245));
  OAI21_X1  g059(.A(G101), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n221), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT65), .B1(new_n223), .B2(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n224), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT1), .B1(new_n225), .B2(G146), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n249), .A2(new_n229), .B1(G128), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT1), .ZN(new_n252));
  AND4_X1   g066(.A1(new_n252), .A2(new_n224), .A3(new_n226), .A4(G128), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n247), .B(KEYINPUT10), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n243), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n250), .A2(G128), .B1(new_n224), .B2(new_n226), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT78), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n235), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n259));
  XNOR2_X1  g073(.A(G143), .B(G146), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT78), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n252), .A3(G128), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT10), .B1(new_n263), .B2(new_n247), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n211), .B1(new_n255), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n262), .B1(new_n256), .B2(new_n257), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT78), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n247), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT10), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n270), .A2(new_n210), .A3(new_n243), .A4(new_n254), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G110), .B(G140), .ZN(new_n273));
  INV_X1    g087(.A(G953), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G227), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n273), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT12), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n221), .A2(new_n246), .ZN(new_n280));
  INV_X1    g094(.A(new_n229), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(new_n224), .B2(new_n248), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n280), .B(new_n262), .C1(new_n282), .C2(new_n259), .ZN(new_n283));
  AOI211_X1 g097(.A(new_n279), .B(new_n210), .C1(new_n268), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n268), .A2(new_n283), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT12), .B1(new_n285), .B2(new_n211), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n271), .B(new_n276), .C1(new_n284), .C2(new_n286), .ZN(new_n287));
  AOI211_X1 g101(.A(G469), .B(G902), .C1(new_n278), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n271), .B1(new_n284), .B2(new_n286), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n276), .B(KEYINPUT77), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n271), .A2(new_n276), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n265), .ZN(new_n292));
  OAI21_X1  g106(.A(G469), .B1(new_n292), .B2(G902), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT79), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n289), .A2(new_n290), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n291), .A2(new_n265), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n296), .B1(new_n299), .B2(new_n190), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT79), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n192), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G214), .B1(G237), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(G224), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT7), .B1(new_n305), .B2(G953), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n251), .A2(G125), .A3(new_n253), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT81), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n311), .B(new_n262), .C1(new_n282), .C2(new_n259), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n312), .B(KEYINPUT81), .C1(new_n311), .C2(new_n240), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n310), .A2(new_n313), .A3(KEYINPUT82), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT82), .B1(new_n310), .B2(new_n313), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT2), .B(G113), .ZN(new_n317));
  AND2_X1   g131(.A1(KEYINPUT67), .A2(G119), .ZN(new_n318));
  NOR2_X1   g132(.A1(KEYINPUT67), .A2(G119), .ZN(new_n319));
  INV_X1    g133(.A(G116), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G119), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(G116), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n317), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n317), .ZN(new_n325));
  OR2_X1    g139(.A1(KEYINPUT67), .A2(G119), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT67), .A2(G119), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(G116), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n323), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n222), .A3(new_n242), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(KEYINPUT5), .A3(new_n329), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G113), .B1(new_n328), .B2(KEYINPUT5), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n247), .B(new_n330), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G122), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n332), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n312), .B(new_n307), .C1(new_n311), .C2(new_n240), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n328), .A2(KEYINPUT5), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n328), .A2(KEYINPUT80), .A3(KEYINPUT5), .A4(new_n329), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n341), .A2(G113), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n330), .A2(new_n221), .A3(new_n246), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n330), .B1(new_n334), .B2(new_n335), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n344), .A2(new_n345), .B1(new_n346), .B2(new_n280), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n337), .B(KEYINPUT8), .Z(new_n348));
  OAI211_X1 g162(.A(new_n338), .B(new_n339), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n190), .B1(new_n316), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n332), .A2(new_n336), .ZN(new_n351));
  INV_X1    g165(.A(new_n337), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(KEYINPUT6), .A3(new_n338), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n355), .A3(new_n352), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n312), .B1(new_n311), .B2(new_n240), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n305), .A2(G953), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n357), .B(new_n358), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n354), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(G210), .B1(G237), .B2(G902), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n350), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n310), .A2(new_n313), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n310), .A2(new_n313), .A3(KEYINPUT82), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n338), .A2(new_n339), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n344), .A2(new_n345), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n346), .A2(new_n280), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n348), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(G902), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n354), .A2(new_n356), .A3(new_n359), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n361), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n304), .B1(new_n363), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n303), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n240), .B1(new_n202), .B2(new_n209), .ZN(new_n379));
  INV_X1    g193(.A(new_n331), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n204), .A2(new_n208), .A3(new_n203), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n203), .B1(G134), .B2(G137), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n205), .A2(new_n207), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n382), .B1(new_n383), .B2(G137), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n381), .B(new_n384), .C1(new_n251), .C2(new_n253), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n379), .A2(new_n380), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n380), .B1(new_n379), .B2(new_n385), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT28), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT70), .B1(new_n386), .B2(KEYINPUT28), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n379), .A2(new_n380), .A3(new_n385), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT70), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT28), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G237), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT68), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT68), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G237), .ZN(new_n398));
  AOI21_X1  g212(.A(G953), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G210), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT26), .B(G101), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n394), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n379), .A2(new_n407), .A3(new_n385), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n379), .B2(new_n385), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n331), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n404), .A3(new_n390), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT31), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT31), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n410), .A2(new_n413), .A3(new_n404), .A4(new_n390), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n406), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G472), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(new_n190), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT71), .B(KEYINPUT32), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n415), .A2(KEYINPUT32), .A3(new_n416), .A4(new_n190), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n410), .A2(new_n390), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n405), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT29), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n388), .A2(new_n389), .A3(new_n404), .A4(new_n393), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n190), .B1(new_n425), .B2(new_n424), .ZN(new_n427));
  OAI21_X1  g241(.A(G472), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n420), .A2(new_n421), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G217), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(G234), .B2(new_n190), .ZN(new_n431));
  INV_X1    g245(.A(G140), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G125), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n311), .A2(G140), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT16), .ZN(new_n435));
  OR3_X1    g249(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n223), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n436), .A3(G146), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n326), .A2(G128), .A3(new_n327), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT24), .B(G110), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT72), .B1(new_n322), .B2(G128), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT72), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n235), .A3(G119), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OR3_X1    g261(.A1(new_n442), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n235), .B1(new_n318), .B2(new_n319), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT23), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n235), .A2(KEYINPUT23), .A3(G119), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n451), .A2(new_n441), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G110), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n440), .B(new_n448), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n433), .A2(new_n434), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(G146), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n451), .A2(new_n454), .A3(new_n441), .A4(new_n452), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n443), .B1(new_n442), .B2(new_n447), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT73), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n439), .B(new_n461), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n460), .A2(new_n462), .A3(KEYINPUT74), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT74), .B1(new_n460), .B2(new_n462), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n455), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT75), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT75), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n467), .B(new_n455), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT22), .B(G137), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n274), .A2(G221), .A3(G234), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n469), .B(new_n470), .Z(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n466), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n465), .A2(KEYINPUT75), .A3(new_n471), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT25), .B1(new_n475), .B2(new_n190), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT25), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n477), .B(G902), .C1(new_n473), .C2(new_n474), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n431), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n431), .A2(G902), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n429), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G475), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT85), .ZN(new_n484));
  NAND2_X1  g298(.A1(KEYINPUT18), .A2(G131), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n396), .A2(new_n398), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n225), .A2(KEYINPUT83), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n487), .A2(G214), .A3(new_n274), .A4(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT83), .B(G143), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n399), .B2(G214), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n486), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT84), .ZN(new_n494));
  INV_X1    g308(.A(G214), .ZN(new_n495));
  AOI211_X1 g309(.A(new_n495), .B(G953), .C1(new_n396), .C2(new_n398), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n489), .B1(new_n496), .B2(new_n491), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT84), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n486), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n456), .B(new_n223), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n490), .A2(new_n492), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n501), .B1(new_n502), .B2(new_n485), .ZN(new_n503));
  OAI21_X1  g317(.A(G131), .B1(new_n490), .B2(new_n492), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n397), .A2(G237), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n395), .A2(KEYINPUT68), .ZN(new_n507));
  OAI211_X1 g321(.A(G214), .B(new_n274), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n491), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n203), .A3(new_n489), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n203), .B1(new_n510), .B2(new_n489), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n440), .B1(new_n513), .B2(KEYINPUT17), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n500), .A2(new_n503), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(G113), .B(G122), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(new_n212), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n484), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  AOI211_X1 g332(.A(KEYINPUT84), .B(new_n485), .C1(new_n510), .C2(new_n489), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n498), .B1(new_n497), .B2(new_n486), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n503), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n514), .A2(new_n512), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n484), .A4(new_n517), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  OAI22_X1  g338(.A1(new_n518), .A2(new_n524), .B1(new_n517), .B2(new_n515), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n483), .B1(new_n525), .B2(new_n190), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT19), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT19), .B1(new_n433), .B2(new_n434), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n223), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n511), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n462), .B(new_n529), .C1(new_n530), .C2(new_n513), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n517), .B1(new_n521), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n518), .B2(new_n524), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT86), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(G475), .A2(G902), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n521), .A2(new_n522), .A3(new_n517), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT85), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n532), .B1(new_n539), .B2(new_n523), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT86), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n536), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT20), .ZN(new_n543));
  INV_X1    g357(.A(new_n537), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(KEYINPUT20), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n534), .A2(KEYINPUT87), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT87), .ZN(new_n547));
  INV_X1    g361(.A(new_n545), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n547), .B1(new_n540), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n526), .B1(new_n543), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n225), .A2(G128), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n235), .A2(G143), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n383), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(G116), .B(G122), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n215), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n320), .A2(KEYINPUT14), .A3(G122), .ZN(new_n559));
  INV_X1    g373(.A(new_n557), .ZN(new_n560));
  OAI211_X1 g374(.A(G107), .B(new_n559), .C1(new_n560), .C2(KEYINPUT14), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n556), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n557), .B(new_n215), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT13), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n553), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n554), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n553), .A2(new_n564), .ZN(new_n567));
  OAI21_X1  g381(.A(G134), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n383), .A2(new_n555), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n563), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n188), .A2(new_n430), .A3(G953), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n562), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n562), .B2(new_n570), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT15), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G478), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n190), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n190), .B1(new_n572), .B2(new_n573), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n575), .A3(G478), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n274), .A2(G952), .ZN(new_n581));
  NAND2_X1  g395(.A1(G234), .A2(G237), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT88), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(G902), .A3(G953), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT21), .B(G898), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n580), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n378), .A2(new_n482), .A3(new_n552), .A4(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  XOR2_X1   g406(.A(new_n574), .B(KEYINPUT33), .Z(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G478), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n578), .A2(G478), .ZN(new_n595));
  NAND2_X1  g409(.A1(G478), .A2(G902), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n552), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n377), .A2(new_n589), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n599), .A2(new_n479), .A3(new_n481), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n405), .A2(new_n394), .B1(new_n411), .B2(KEYINPUT31), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n601), .B2(new_n414), .ZN(new_n602));
  OR3_X1    g416(.A1(new_n602), .A2(KEYINPUT89), .A3(new_n416), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n415), .A2(new_n190), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(G472), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(KEYINPUT89), .A3(new_n417), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n598), .A2(new_n600), .A3(new_n302), .A4(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT34), .B(G104), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  INV_X1    g426(.A(KEYINPUT93), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n526), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n515), .A2(new_n517), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n523), .B2(new_n539), .ZN(new_n616));
  OAI21_X1  g430(.A(G475), .B1(new_n616), .B2(G902), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT93), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n614), .A2(new_n618), .A3(new_n580), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n540), .A2(KEYINPUT86), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n535), .B(new_n532), .C1(new_n539), .C2(new_n523), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n620), .A2(new_n621), .A3(new_n548), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT92), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n622), .B1(new_n543), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n542), .A2(KEYINPUT92), .A3(KEYINPUT20), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n619), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND4_X1   g440(.A1(new_n302), .A2(new_n626), .A3(new_n600), .A4(new_n607), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT35), .B(G107), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NOR2_X1   g443(.A1(new_n472), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n465), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n480), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n603), .A2(new_n606), .B1(new_n479), .B2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n378), .A2(new_n633), .A3(new_n552), .A4(new_n590), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT37), .B(G110), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT94), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n634), .B(new_n636), .ZN(G12));
  NOR3_X1   g451(.A1(new_n620), .A2(new_n621), .A3(new_n544), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT20), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n623), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n622), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n625), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n304), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n362), .B1(new_n350), .B2(new_n360), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n374), .A2(new_n361), .A3(new_n375), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n619), .ZN(new_n647));
  INV_X1    g461(.A(new_n584), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n649), .B2(new_n586), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n650), .A2(KEYINPUT95), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(KEYINPUT95), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n642), .A2(new_n646), .A3(new_n647), .A4(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT96), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n626), .A2(KEYINPUT96), .A3(new_n646), .A4(new_n653), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n479), .A2(new_n632), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n429), .A3(new_n302), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n656), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  XOR2_X1   g476(.A(new_n653), .B(KEYINPUT39), .Z(new_n663));
  NOR2_X1   g477(.A1(new_n303), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n665), .A2(KEYINPUT40), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(KEYINPUT40), .ZN(new_n667));
  INV_X1    g481(.A(new_n658), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n405), .B1(new_n390), .B2(new_n410), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n386), .A2(new_n387), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n190), .B1(new_n670), .B2(new_n404), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n420), .A2(new_n421), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n644), .A2(new_n645), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n304), .A3(new_n580), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n674), .A2(new_n552), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n666), .A2(new_n667), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT98), .B(G143), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G45));
  NAND4_X1  g496(.A1(new_n658), .A2(new_n302), .A3(new_n429), .A4(new_n646), .ZN(new_n683));
  INV_X1    g497(.A(new_n597), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n550), .B1(KEYINPUT20), .B2(new_n542), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n684), .B(new_n653), .C1(new_n685), .C2(new_n526), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n223), .ZN(G48));
  AOI21_X1  g502(.A(new_n210), .B1(new_n268), .B2(new_n283), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT12), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n690), .A2(new_n291), .B1(new_n272), .B2(new_n277), .ZN(new_n691));
  OAI21_X1  g505(.A(G469), .B1(new_n691), .B2(G902), .ZN(new_n692));
  INV_X1    g506(.A(new_n191), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n278), .A2(new_n287), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n296), .A3(new_n190), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n429), .A2(new_n479), .A3(new_n481), .A4(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n598), .A3(new_n599), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NAND3_X1  g515(.A1(new_n626), .A2(new_n698), .A3(new_n599), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  AND2_X1   g517(.A1(new_n428), .A2(new_n421), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n704), .A2(new_n420), .B1(new_n479), .B2(new_n632), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT99), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n706), .B1(new_n377), .B2(new_n696), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n296), .B1(new_n694), .B2(new_n190), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n288), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n646), .A2(new_n709), .A3(KEYINPUT99), .A4(new_n693), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n705), .A2(new_n552), .A3(new_n590), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  NAND2_X1  g527(.A1(new_n646), .A2(new_n580), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n696), .A2(new_n589), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n552), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT100), .ZN(new_n717));
  OAI21_X1  g531(.A(G472), .B1(new_n602), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n604), .A2(KEYINPUT100), .A3(new_n416), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND4_X1   g534(.A1(KEYINPUT101), .A2(new_n720), .A3(new_n479), .A4(new_n481), .ZN(new_n721));
  INV_X1    g535(.A(new_n481), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n468), .A2(new_n472), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n458), .A2(new_n459), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n439), .A2(KEYINPUT73), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n439), .A2(KEYINPUT73), .ZN(new_n726));
  INV_X1    g540(.A(new_n457), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n724), .A2(new_n725), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT74), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n460), .A2(new_n462), .A3(KEYINPUT74), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n467), .B1(new_n732), .B2(new_n455), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n723), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n474), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n190), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n477), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n475), .A2(KEYINPUT25), .A3(new_n190), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n722), .B1(new_n739), .B2(new_n431), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT101), .B1(new_n740), .B2(new_n720), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n716), .B1(new_n721), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT102), .B(G122), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G24));
  AOI22_X1  g558(.A1(new_n479), .A2(new_n632), .B1(new_n718), .B2(new_n719), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n711), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n686), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n311), .ZN(G27));
  OAI21_X1  g562(.A(new_n693), .B1(new_n300), .B2(new_n288), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n644), .A2(new_n304), .A3(new_n645), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n429), .A3(new_n479), .A4(new_n481), .ZN(new_n752));
  OR3_X1    g566(.A1(new_n686), .A2(new_n752), .A3(KEYINPUT103), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT103), .B1(new_n686), .B2(new_n752), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n740), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT32), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n417), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n757), .B1(new_n704), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n686), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(KEYINPUT42), .A3(new_n761), .A4(new_n751), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n756), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  NAND4_X1  g578(.A1(new_n626), .A2(new_n482), .A3(new_n653), .A4(new_n751), .ZN(new_n765));
  XOR2_X1   g579(.A(KEYINPUT104), .B(G134), .Z(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G36));
  AND2_X1   g581(.A1(new_n552), .A2(KEYINPUT106), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n684), .B1(new_n552), .B2(KEYINPUT106), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT43), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n552), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n771), .A2(KEYINPUT43), .A3(new_n597), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n773), .A2(new_n603), .A3(new_n606), .A4(new_n658), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(G469), .A2(G902), .ZN(new_n777));
  OAI21_X1  g591(.A(G469), .B1(new_n292), .B2(KEYINPUT45), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT105), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n292), .A2(KEYINPUT45), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n778), .B2(new_n779), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n777), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT46), .B(new_n777), .C1(new_n780), .C2(new_n782), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n695), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n693), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n663), .ZN(new_n789));
  INV_X1    g603(.A(new_n750), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n774), .B2(new_n775), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n776), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(KEYINPUT107), .B(G137), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(G39));
  NOR4_X1   g609(.A1(new_n686), .A2(new_n429), .A3(new_n740), .A4(new_n750), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n787), .A2(KEYINPUT47), .A3(new_n693), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT47), .B1(new_n787), .B2(new_n693), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(KEYINPUT108), .B(G140), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(G42));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n742), .A2(new_n591), .A3(new_n608), .A4(new_n702), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n580), .B(KEYINPUT111), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n685), .A2(new_n526), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(new_n600), .A3(new_n302), .A4(new_n607), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n634), .A2(new_n699), .A3(new_n806), .A4(new_n712), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n614), .A2(new_n618), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n804), .A2(new_n653), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n810), .A2(new_n811), .A3(new_n750), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n642), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n658), .A2(new_n720), .A3(new_n751), .ZN(new_n814));
  OAI22_X1  g628(.A1(new_n813), .A2(new_n659), .B1(new_n814), .B2(new_n686), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n642), .A2(new_n647), .A3(new_n653), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n752), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n809), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n686), .A2(new_n814), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n705), .A2(new_n642), .A3(new_n812), .A4(new_n302), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n765), .A3(KEYINPUT112), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n808), .A2(new_n822), .A3(new_n763), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n686), .B1(new_n746), .B2(new_n683), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n653), .B(KEYINPUT113), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n749), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n673), .A3(new_n479), .A4(new_n632), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n827), .A2(new_n552), .A3(new_n714), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT52), .B1(new_n661), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n661), .A2(new_n829), .A3(KEYINPUT52), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n823), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND4_X1   g650(.A1(KEYINPUT53), .A2(new_n808), .A3(new_n763), .A4(new_n822), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n833), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n802), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n721), .A2(new_n741), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n584), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n773), .A2(new_n711), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n757), .A2(new_n673), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n696), .A2(new_n750), .A3(new_n584), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n598), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n773), .A2(new_n760), .A3(new_n846), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n849), .A2(KEYINPUT48), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(KEYINPUT48), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n677), .A2(new_n304), .A3(new_n696), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n843), .A2(new_n770), .A3(new_n772), .A4(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT50), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n773), .A2(new_n745), .A3(new_n846), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n845), .A2(new_n552), .A3(new_n597), .A4(new_n846), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n773), .A2(new_n790), .A3(new_n843), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n692), .A2(new_n695), .ZN(new_n859));
  INV_X1    g673(.A(new_n192), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n797), .A2(new_n798), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n856), .B(new_n857), .C1(new_n858), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n852), .B1(new_n864), .B2(KEYINPUT51), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(KEYINPUT116), .A3(KEYINPUT51), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT50), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n854), .B(new_n867), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n858), .A2(new_n862), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n856), .A2(new_n857), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n868), .A2(KEYINPUT51), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n865), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n837), .A2(new_n875), .A3(new_n833), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n808), .A2(new_n822), .A3(new_n763), .A4(KEYINPUT53), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n661), .A2(KEYINPUT52), .A3(new_n829), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n830), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT115), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n876), .A2(new_n880), .B1(new_n834), .B2(new_n835), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n840), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n836), .A2(new_n838), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(KEYINPUT114), .A3(KEYINPUT54), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n841), .A2(new_n874), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(G953), .B1(new_n885), .B2(KEYINPUT117), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n581), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n740), .A2(new_n304), .A3(new_n860), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT109), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n890), .A2(new_n768), .A3(new_n769), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n891), .A2(KEYINPUT110), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(KEYINPUT110), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n859), .B(KEYINPUT49), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n894), .A2(new_n677), .A3(new_n673), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n886), .A2(new_n888), .A3(new_n896), .ZN(G75));
  NOR2_X1   g711(.A1(new_n881), .A2(new_n190), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT56), .B1(new_n898), .B2(G210), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n354), .A2(new_n356), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT118), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n359), .B(KEYINPUT55), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n901), .B(new_n902), .Z(new_n903));
  AND2_X1   g717(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n899), .A2(new_n903), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n274), .A2(G952), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G51));
  AOI21_X1  g721(.A(new_n875), .B1(new_n837), .B2(new_n833), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT115), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n836), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT54), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n882), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n777), .B(KEYINPUT57), .Z(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n694), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n780), .A2(new_n782), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n898), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n906), .B1(new_n915), .B2(new_n917), .ZN(G54));
  NAND3_X1  g732(.A1(new_n898), .A2(KEYINPUT58), .A3(G475), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n620), .A2(new_n621), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n919), .A2(KEYINPUT119), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n906), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n919), .B2(new_n921), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT119), .B1(new_n919), .B2(new_n921), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(G60));
  INV_X1    g740(.A(new_n593), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n841), .A2(new_n882), .A3(new_n884), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n596), .B(KEYINPUT59), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n912), .A2(new_n927), .A3(new_n929), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n906), .A3(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT60), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n910), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n475), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n906), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n910), .A2(new_n631), .A3(new_n935), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n938), .A2(KEYINPUT121), .A3(KEYINPUT61), .A4(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n937), .B1(new_n881), .B2(new_n934), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n941), .A2(new_n939), .A3(KEYINPUT61), .A4(new_n923), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT121), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n941), .A2(new_n939), .A3(new_n923), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT120), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n947), .B1(new_n946), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(G66));
  OAI21_X1  g765(.A(G953), .B1(new_n587), .B2(new_n305), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n808), .B2(G953), .ZN(new_n953));
  INV_X1    g767(.A(new_n901), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(G898), .B2(new_n274), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT122), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n953), .B(new_n956), .ZN(G69));
  NOR2_X1   g771(.A1(new_n408), .A2(new_n409), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n527), .A2(new_n528), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n958), .B(new_n959), .Z(new_n960));
  NAND3_X1  g774(.A1(new_n664), .A2(new_n482), .A3(new_n790), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n598), .A2(new_n805), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n799), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n824), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n661), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT123), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT123), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n661), .A2(new_n968), .A3(new_n965), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n680), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n793), .B(new_n964), .C1(new_n971), .C2(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n971), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n960), .B1(new_n977), .B2(G953), .ZN(new_n978));
  INV_X1    g792(.A(new_n960), .ZN(new_n979));
  AND4_X1   g793(.A1(new_n646), .A2(new_n760), .A3(new_n771), .A4(new_n580), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n817), .B1(new_n980), .B2(new_n789), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n981), .A2(new_n763), .A3(new_n799), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n793), .A2(new_n970), .A3(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n983), .A2(new_n274), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n649), .A2(G953), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT125), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n979), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n978), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n274), .B1(G227), .B2(G900), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(G72));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n991));
  INV_X1    g805(.A(new_n669), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n977), .A2(new_n808), .ZN(new_n993));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  AOI21_X1  g809(.A(new_n992), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n793), .A2(new_n808), .A3(new_n970), .A4(new_n982), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n995), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n998), .A2(new_n405), .A3(new_n390), .A4(new_n410), .ZN(new_n999));
  INV_X1    g813(.A(new_n995), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n423), .B2(new_n411), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT126), .Z(new_n1002));
  OAI211_X1 g816(.A(new_n999), .B(new_n923), .C1(new_n839), .C2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n991), .B1(new_n996), .B2(new_n1003), .ZN(new_n1004));
  AOI211_X1 g818(.A(new_n404), .B(new_n422), .C1(new_n997), .C2(new_n995), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n839), .A2(new_n1002), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n1005), .A2(new_n1006), .A3(new_n906), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1000), .B1(new_n977), .B2(new_n808), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n1007), .B(KEYINPUT127), .C1(new_n1008), .C2(new_n992), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1004), .A2(new_n1009), .ZN(G57));
endmodule


