

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593;

  NAND2_X1 U323 ( .A1(n418), .A2(n417), .ZN(n420) );
  XNOR2_X1 U324 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U325 ( .A(G36GAT), .B(G190GAT), .Z(n376) );
  XNOR2_X1 U326 ( .A(n373), .B(n432), .ZN(n374) );
  INV_X1 U327 ( .A(KEYINPUT25), .ZN(n385) );
  NOR2_X1 U328 ( .A1(n591), .A2(n421), .ZN(n423) );
  XNOR2_X1 U329 ( .A(n376), .B(n291), .ZN(n377) );
  AND2_X1 U330 ( .A1(G226GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U331 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n467) );
  XNOR2_X1 U332 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U333 ( .A(n386), .B(n385), .ZN(n387) );
  NAND2_X1 U334 ( .A1(n388), .A2(n387), .ZN(n413) );
  XNOR2_X1 U335 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n482) );
  INV_X1 U336 ( .A(G197GAT), .ZN(n364) );
  XNOR2_X1 U337 ( .A(n365), .B(n364), .ZN(n373) );
  INV_X1 U338 ( .A(KEYINPUT101), .ZN(n419) );
  XNOR2_X1 U339 ( .A(n326), .B(n456), .ZN(n327) );
  XNOR2_X1 U340 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n479) );
  XNOR2_X1 U341 ( .A(n420), .B(n419), .ZN(n502) );
  XNOR2_X1 U342 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U343 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U344 ( .A(n461), .B(n460), .ZN(n466) );
  OR2_X1 U345 ( .A1(n536), .A2(n505), .ZN(n462) );
  INV_X1 U346 ( .A(G43GAT), .ZN(n463) );
  XNOR2_X1 U347 ( .A(n462), .B(KEYINPUT38), .ZN(n518) );
  XNOR2_X1 U348 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n490) );
  XNOR2_X1 U349 ( .A(n463), .B(KEYINPUT40), .ZN(n464) );
  XNOR2_X1 U350 ( .A(n491), .B(n490), .ZN(G1351GAT) );
  XNOR2_X1 U351 ( .A(n465), .B(n464), .ZN(G1330GAT) );
  XOR2_X1 U352 ( .A(KEYINPUT20), .B(G71GAT), .Z(n293) );
  XNOR2_X1 U353 ( .A(G169GAT), .B(G113GAT), .ZN(n292) );
  XNOR2_X1 U354 ( .A(n293), .B(n292), .ZN(n309) );
  XOR2_X1 U355 ( .A(G15GAT), .B(G127GAT), .Z(n332) );
  XOR2_X1 U356 ( .A(G134GAT), .B(G190GAT), .Z(n295) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(G99GAT), .ZN(n294) );
  XNOR2_X1 U358 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U359 ( .A(n332), .B(n296), .Z(n298) );
  NAND2_X1 U360 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U361 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U362 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n300) );
  XNOR2_X1 U363 ( .A(KEYINPUT85), .B(G176GAT), .ZN(n299) );
  XNOR2_X1 U364 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U365 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U366 ( .A(G183GAT), .B(KEYINPUT18), .Z(n304) );
  XNOR2_X1 U367 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n303) );
  XNOR2_X1 U368 ( .A(n304), .B(n303), .ZN(n372) );
  XNOR2_X1 U369 ( .A(G120GAT), .B(KEYINPUT0), .ZN(n305) );
  XNOR2_X1 U370 ( .A(n305), .B(KEYINPUT84), .ZN(n400) );
  XNOR2_X1 U371 ( .A(n372), .B(n400), .ZN(n306) );
  XNOR2_X1 U372 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U373 ( .A(n309), .B(n308), .ZN(n549) );
  INV_X1 U374 ( .A(n549), .ZN(n541) );
  XNOR2_X1 U375 ( .A(KEYINPUT36), .B(KEYINPUT105), .ZN(n331) );
  XOR2_X1 U376 ( .A(KEYINPUT9), .B(KEYINPUT75), .Z(n311) );
  NAND2_X1 U377 ( .A1(G232GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U378 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U379 ( .A(KEYINPUT78), .B(n312), .ZN(n330) );
  XOR2_X1 U380 ( .A(KEYINPUT10), .B(n376), .Z(n314) );
  XOR2_X1 U381 ( .A(G134GAT), .B(KEYINPUT79), .Z(n399) );
  XNOR2_X1 U382 ( .A(G106GAT), .B(n399), .ZN(n313) );
  XNOR2_X1 U383 ( .A(n314), .B(n313), .ZN(n316) );
  INV_X1 U384 ( .A(KEYINPUT77), .ZN(n315) );
  XNOR2_X1 U385 ( .A(n316), .B(n315), .ZN(n321) );
  XOR2_X1 U386 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n318) );
  XNOR2_X1 U387 ( .A(G92GAT), .B(KEYINPUT76), .ZN(n317) );
  XNOR2_X1 U388 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U389 ( .A(G218GAT), .B(n319), .ZN(n320) );
  NAND2_X1 U390 ( .A1(n321), .A2(n320), .ZN(n323) );
  OR2_X1 U391 ( .A1(n321), .A2(n320), .ZN(n322) );
  NAND2_X1 U392 ( .A1(n323), .A2(n322), .ZN(n328) );
  XOR2_X1 U393 ( .A(G29GAT), .B(G43GAT), .Z(n325) );
  XNOR2_X1 U394 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n324) );
  XNOR2_X1 U395 ( .A(n325), .B(n324), .ZN(n434) );
  XOR2_X1 U396 ( .A(G50GAT), .B(G162GAT), .Z(n353) );
  XNOR2_X1 U397 ( .A(n434), .B(n353), .ZN(n326) );
  XNOR2_X1 U398 ( .A(G99GAT), .B(G85GAT), .ZN(n456) );
  XNOR2_X1 U399 ( .A(n330), .B(n329), .ZN(n471) );
  XOR2_X1 U400 ( .A(n331), .B(n471), .Z(n591) );
  XOR2_X1 U401 ( .A(G22GAT), .B(G155GAT), .Z(n352) );
  XOR2_X1 U402 ( .A(n352), .B(G78GAT), .Z(n334) );
  XNOR2_X1 U403 ( .A(n332), .B(G211GAT), .ZN(n333) );
  XNOR2_X1 U404 ( .A(n334), .B(n333), .ZN(n339) );
  XNOR2_X1 U405 ( .A(G71GAT), .B(G57GAT), .ZN(n335) );
  XNOR2_X1 U406 ( .A(n335), .B(KEYINPUT13), .ZN(n455) );
  XOR2_X1 U407 ( .A(n455), .B(KEYINPUT81), .Z(n337) );
  NAND2_X1 U408 ( .A1(G231GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U409 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U410 ( .A(n339), .B(n338), .Z(n341) );
  XNOR2_X1 U411 ( .A(G1GAT), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U412 ( .A(n341), .B(n340), .ZN(n349) );
  XOR2_X1 U413 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n343) );
  XNOR2_X1 U414 ( .A(G8GAT), .B(G64GAT), .ZN(n342) );
  XNOR2_X1 U415 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U416 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n345) );
  XNOR2_X1 U417 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n344) );
  XNOR2_X1 U418 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U419 ( .A(n347), .B(n346), .Z(n348) );
  XNOR2_X1 U420 ( .A(n349), .B(n348), .ZN(n559) );
  XOR2_X1 U421 ( .A(G204GAT), .B(KEYINPUT23), .Z(n351) );
  XNOR2_X1 U422 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n350) );
  XNOR2_X1 U423 ( .A(n351), .B(n350), .ZN(n357) );
  XOR2_X1 U424 ( .A(KEYINPUT88), .B(KEYINPUT90), .Z(n355) );
  XNOR2_X1 U425 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U426 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U427 ( .A(n357), .B(n356), .Z(n359) );
  NAND2_X1 U428 ( .A1(G228GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U429 ( .A(n359), .B(n358), .ZN(n361) );
  XNOR2_X1 U430 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n360) );
  XNOR2_X1 U431 ( .A(n360), .B(KEYINPUT2), .ZN(n395) );
  XOR2_X1 U432 ( .A(n361), .B(n395), .Z(n368) );
  XOR2_X1 U433 ( .A(KEYINPUT21), .B(G218GAT), .Z(n363) );
  XNOR2_X1 U434 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n362) );
  XNOR2_X1 U435 ( .A(n363), .B(n362), .ZN(n365) );
  XNOR2_X1 U436 ( .A(G106GAT), .B(G78GAT), .ZN(n366) );
  XNOR2_X1 U437 ( .A(n366), .B(G148GAT), .ZN(n443) );
  XNOR2_X1 U438 ( .A(n373), .B(n443), .ZN(n367) );
  XNOR2_X1 U439 ( .A(n368), .B(n367), .ZN(n486) );
  NOR2_X1 U440 ( .A1(n549), .A2(n486), .ZN(n369) );
  XNOR2_X1 U441 ( .A(n369), .B(KEYINPUT26), .ZN(n567) );
  INV_X1 U442 ( .A(n567), .ZN(n381) );
  XOR2_X1 U443 ( .A(G64GAT), .B(G92GAT), .Z(n371) );
  XNOR2_X1 U444 ( .A(G176GAT), .B(G204GAT), .ZN(n370) );
  XNOR2_X1 U445 ( .A(n371), .B(n370), .ZN(n454) );
  XNOR2_X1 U446 ( .A(n372), .B(n454), .ZN(n380) );
  XOR2_X1 U447 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n375) );
  XOR2_X1 U448 ( .A(G169GAT), .B(G8GAT), .Z(n432) );
  XNOR2_X1 U449 ( .A(n375), .B(n374), .ZN(n378) );
  XOR2_X1 U450 ( .A(n380), .B(n379), .Z(n383) );
  XNOR2_X1 U451 ( .A(n383), .B(KEYINPUT27), .ZN(n414) );
  NOR2_X1 U452 ( .A1(n381), .A2(n414), .ZN(n382) );
  XOR2_X1 U453 ( .A(KEYINPUT100), .B(n382), .Z(n388) );
  OR2_X1 U454 ( .A1(n383), .A2(n541), .ZN(n384) );
  NAND2_X1 U455 ( .A1(n486), .A2(n384), .ZN(n386) );
  XOR2_X1 U456 ( .A(KEYINPUT94), .B(G57GAT), .Z(n390) );
  XNOR2_X1 U457 ( .A(G127GAT), .B(G155GAT), .ZN(n389) );
  XNOR2_X1 U458 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U459 ( .A(G85GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U460 ( .A(G29GAT), .B(G148GAT), .ZN(n391) );
  XNOR2_X1 U461 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U462 ( .A(n394), .B(n393), .ZN(n412) );
  XOR2_X1 U463 ( .A(n395), .B(KEYINPUT1), .Z(n397) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U466 ( .A(n399), .B(n398), .Z(n402) );
  XOR2_X1 U467 ( .A(G113GAT), .B(G1GAT), .Z(n437) );
  XNOR2_X1 U468 ( .A(n437), .B(n400), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n402), .B(n401), .ZN(n410) );
  XOR2_X1 U470 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n404) );
  XNOR2_X1 U471 ( .A(KEYINPUT91), .B(KEYINPUT4), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U473 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n406) );
  XNOR2_X1 U474 ( .A(KEYINPUT93), .B(KEYINPUT95), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U476 ( .A(n408), .B(n407), .Z(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U478 ( .A(n412), .B(n411), .ZN(n537) );
  NAND2_X1 U479 ( .A1(n413), .A2(n537), .ZN(n418) );
  XOR2_X1 U480 ( .A(n486), .B(KEYINPUT28), .Z(n552) );
  NOR2_X1 U481 ( .A1(n537), .A2(n414), .ZN(n415) );
  XNOR2_X1 U482 ( .A(n415), .B(KEYINPUT99), .ZN(n547) );
  NOR2_X1 U483 ( .A1(n552), .A2(n547), .ZN(n416) );
  NAND2_X1 U484 ( .A1(n541), .A2(n416), .ZN(n417) );
  NAND2_X1 U485 ( .A1(n559), .A2(n502), .ZN(n421) );
  XNOR2_X1 U486 ( .A(KEYINPUT106), .B(KEYINPUT37), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n536) );
  XOR2_X1 U488 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n425) );
  XNOR2_X1 U489 ( .A(G22GAT), .B(G15GAT), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U491 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n427) );
  XNOR2_X1 U492 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n442) );
  XOR2_X1 U495 ( .A(G141GAT), .B(G197GAT), .Z(n431) );
  XNOR2_X1 U496 ( .A(G50GAT), .B(G36GAT), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n433) );
  XOR2_X1 U498 ( .A(n433), .B(n432), .Z(n440) );
  XOR2_X1 U499 ( .A(n434), .B(KEYINPUT68), .Z(n436) );
  NAND2_X1 U500 ( .A1(G229GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U504 ( .A(n442), .B(n441), .ZN(n521) );
  XNOR2_X1 U505 ( .A(n443), .B(KEYINPUT74), .ZN(n447) );
  INV_X1 U506 ( .A(n447), .ZN(n445) );
  AND2_X1 U507 ( .A1(G230GAT), .A2(G233GAT), .ZN(n446) );
  INV_X1 U508 ( .A(n446), .ZN(n444) );
  NAND2_X1 U509 ( .A1(n445), .A2(n444), .ZN(n449) );
  NAND2_X1 U510 ( .A1(n447), .A2(n446), .ZN(n448) );
  NAND2_X1 U511 ( .A1(n449), .A2(n448), .ZN(n453) );
  XOR2_X1 U512 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n451) );
  XNOR2_X1 U513 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n450) );
  XNOR2_X1 U514 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U515 ( .A(n453), .B(n452), .ZN(n461) );
  XOR2_X1 U516 ( .A(n455), .B(n454), .Z(n459) );
  XNOR2_X1 U517 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n457), .B(n456), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n521), .A2(n466), .ZN(n505) );
  NOR2_X1 U520 ( .A1(n541), .A2(n518), .ZN(n465) );
  INV_X1 U521 ( .A(n471), .ZN(n576) );
  XNOR2_X1 U522 ( .A(n466), .B(KEYINPUT41), .ZN(n570) );
  NAND2_X1 U523 ( .A1(n570), .A2(n521), .ZN(n468) );
  NAND2_X1 U524 ( .A1(n469), .A2(n559), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(KEYINPUT115), .ZN(n472) );
  NAND2_X1 U526 ( .A1(n472), .A2(n471), .ZN(n473) );
  XNOR2_X1 U527 ( .A(n473), .B(KEYINPUT47), .ZN(n478) );
  NOR2_X1 U528 ( .A1(n591), .A2(n559), .ZN(n474) );
  XNOR2_X1 U529 ( .A(n474), .B(KEYINPUT45), .ZN(n475) );
  NAND2_X1 U530 ( .A1(n475), .A2(n466), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n476), .A2(n521), .ZN(n477) );
  NOR2_X1 U532 ( .A1(n478), .A2(n477), .ZN(n480) );
  XNOR2_X1 U533 ( .A(n480), .B(n479), .ZN(n548) );
  XOR2_X1 U534 ( .A(n383), .B(KEYINPUT121), .Z(n481) );
  NOR2_X1 U535 ( .A1(n548), .A2(n481), .ZN(n483) );
  XNOR2_X1 U536 ( .A(n483), .B(n482), .ZN(n484) );
  NAND2_X1 U537 ( .A1(n484), .A2(n537), .ZN(n485) );
  XNOR2_X1 U538 ( .A(n485), .B(KEYINPUT65), .ZN(n495) );
  NAND2_X1 U539 ( .A1(n486), .A2(n495), .ZN(n487) );
  XNOR2_X1 U540 ( .A(n487), .B(KEYINPUT55), .ZN(n488) );
  NAND2_X1 U541 ( .A1(n488), .A2(n549), .ZN(n489) );
  XNOR2_X1 U542 ( .A(n489), .B(KEYINPUT123), .ZN(n580) );
  NAND2_X1 U543 ( .A1(n576), .A2(n580), .ZN(n491) );
  NAND2_X1 U544 ( .A1(n580), .A2(n570), .ZN(n494) );
  XOR2_X1 U545 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n492) );
  XNOR2_X1 U546 ( .A(n492), .B(G176GAT), .ZN(n493) );
  XNOR2_X1 U547 ( .A(n494), .B(n493), .ZN(G1349GAT) );
  INV_X1 U548 ( .A(G204GAT), .ZN(n500) );
  XOR2_X1 U549 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n498) );
  NAND2_X1 U550 ( .A1(n495), .A2(n567), .ZN(n496) );
  XNOR2_X1 U551 ( .A(n496), .B(KEYINPUT125), .ZN(n588) );
  INV_X1 U552 ( .A(n588), .ZN(n590) );
  OR2_X1 U553 ( .A1(n590), .A2(n466), .ZN(n497) );
  XNOR2_X1 U554 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U555 ( .A(n500), .B(n499), .ZN(G1353GAT) );
  NOR2_X1 U556 ( .A1(n576), .A2(n559), .ZN(n501) );
  XNOR2_X1 U557 ( .A(KEYINPUT16), .B(n501), .ZN(n503) );
  NAND2_X1 U558 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U559 ( .A(n504), .B(KEYINPUT102), .ZN(n523) );
  OR2_X1 U560 ( .A1(n523), .A2(n505), .ZN(n512) );
  NOR2_X1 U561 ( .A1(n537), .A2(n512), .ZN(n506) );
  XOR2_X1 U562 ( .A(n506), .B(KEYINPUT34), .Z(n507) );
  XNOR2_X1 U563 ( .A(G1GAT), .B(n507), .ZN(G1324GAT) );
  NOR2_X1 U564 ( .A1(n383), .A2(n512), .ZN(n509) );
  XNOR2_X1 U565 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n508) );
  XNOR2_X1 U566 ( .A(n509), .B(n508), .ZN(G1325GAT) );
  NOR2_X1 U567 ( .A1(n541), .A2(n512), .ZN(n511) );
  XNOR2_X1 U568 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n510) );
  XNOR2_X1 U569 ( .A(n511), .B(n510), .ZN(G1326GAT) );
  INV_X1 U570 ( .A(n552), .ZN(n544) );
  NOR2_X1 U571 ( .A1(n544), .A2(n512), .ZN(n513) );
  XOR2_X1 U572 ( .A(KEYINPUT104), .B(n513), .Z(n514) );
  XNOR2_X1 U573 ( .A(G22GAT), .B(n514), .ZN(G1327GAT) );
  NOR2_X1 U574 ( .A1(n518), .A2(n537), .ZN(n516) );
  XNOR2_X1 U575 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n515) );
  XNOR2_X1 U576 ( .A(n516), .B(n515), .ZN(G1328GAT) );
  NOR2_X1 U577 ( .A1(n518), .A2(n383), .ZN(n517) );
  XOR2_X1 U578 ( .A(G36GAT), .B(n517), .Z(G1329GAT) );
  NOR2_X1 U579 ( .A1(n518), .A2(n544), .ZN(n520) );
  XNOR2_X1 U580 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n519) );
  XNOR2_X1 U581 ( .A(n520), .B(n519), .ZN(G1331GAT) );
  INV_X1 U582 ( .A(n521), .ZN(n553) );
  NAND2_X1 U583 ( .A1(n570), .A2(n553), .ZN(n522) );
  XNOR2_X1 U584 ( .A(n522), .B(KEYINPUT108), .ZN(n535) );
  OR2_X1 U585 ( .A1(n523), .A2(n535), .ZN(n531) );
  NOR2_X1 U586 ( .A1(n537), .A2(n531), .ZN(n525) );
  XNOR2_X1 U587 ( .A(KEYINPUT42), .B(KEYINPUT109), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G57GAT), .B(n526), .ZN(G1332GAT) );
  NOR2_X1 U590 ( .A1(n383), .A2(n531), .ZN(n527) );
  XOR2_X1 U591 ( .A(KEYINPUT110), .B(n527), .Z(n528) );
  XNOR2_X1 U592 ( .A(G64GAT), .B(n528), .ZN(G1333GAT) );
  NOR2_X1 U593 ( .A1(n541), .A2(n531), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(G1334GAT) );
  NOR2_X1 U596 ( .A1(n544), .A2(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(KEYINPUT43), .B(KEYINPUT112), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G78GAT), .B(n534), .ZN(G1335GAT) );
  OR2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n543) );
  NOR2_X1 U601 ( .A1(n537), .A2(n543), .ZN(n539) );
  XNOR2_X1 U602 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1336GAT) );
  NOR2_X1 U604 ( .A1(n383), .A2(n543), .ZN(n540) );
  XOR2_X1 U605 ( .A(G92GAT), .B(n540), .Z(G1337GAT) );
  NOR2_X1 U606 ( .A1(n541), .A2(n543), .ZN(n542) );
  XOR2_X1 U607 ( .A(G99GAT), .B(n542), .Z(G1338GAT) );
  NOR2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U609 ( .A(KEYINPUT44), .B(n545), .Z(n546) );
  XNOR2_X1 U610 ( .A(G106GAT), .B(n546), .ZN(G1339GAT) );
  NOR2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n568) );
  NAND2_X1 U612 ( .A1(n568), .A2(n549), .ZN(n550) );
  XNOR2_X1 U613 ( .A(KEYINPUT116), .B(n550), .ZN(n551) );
  NOR2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n563) );
  NAND2_X1 U615 ( .A1(n563), .A2(n521), .ZN(n554) );
  XNOR2_X1 U616 ( .A(n554), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n556) );
  NAND2_X1 U618 ( .A1(n563), .A2(n570), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n556), .B(n555), .ZN(n558) );
  XOR2_X1 U620 ( .A(G120GAT), .B(KEYINPUT117), .Z(n557) );
  XNOR2_X1 U621 ( .A(n558), .B(n557), .ZN(G1341GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n561) );
  INV_X1 U623 ( .A(n559), .ZN(n587) );
  NAND2_X1 U624 ( .A1(n563), .A2(n587), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U626 ( .A(G127GAT), .B(n562), .ZN(G1342GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n565) );
  NAND2_X1 U628 ( .A1(n563), .A2(n576), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(G134GAT), .B(n566), .ZN(G1343GAT) );
  AND2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n521), .A2(n575), .ZN(n569) );
  XNOR2_X1 U633 ( .A(G141GAT), .B(n569), .ZN(G1344GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n572) );
  NAND2_X1 U635 ( .A1(n575), .A2(n570), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G148GAT), .B(n573), .ZN(G1345GAT) );
  NAND2_X1 U638 ( .A1(n575), .A2(n587), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U642 ( .A1(n580), .A2(n521), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT124), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n587), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U647 ( .A1(n521), .A2(n588), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT60), .ZN(n584) );
  INV_X1 U649 ( .A(KEYINPUT59), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

