//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n187));
  INV_X1    g001(.A(G217), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(G234), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(G125), .ZN(new_n195));
  INV_X1    g009(.A(G125), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n194), .B1(new_n198), .B2(new_n192), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  OAI211_X1 g015(.A(G146), .B(new_n194), .C1(new_n198), .C2(new_n192), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G119), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT24), .B(G110), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n206), .B2(G128), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(new_n207), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n210), .B1(G110), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n203), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G137), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n217), .B(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n198), .A2(G146), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n196), .A2(KEYINPUT16), .A3(G140), .ZN(new_n222));
  XNOR2_X1  g036(.A(G125), .B(G140), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(KEYINPUT16), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n221), .B1(new_n224), .B2(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n208), .A2(new_n209), .ZN(new_n226));
  INV_X1    g040(.A(G110), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n212), .A2(new_n213), .A3(new_n227), .A4(new_n207), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT69), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(new_n200), .ZN(new_n231));
  AND4_X1   g045(.A1(KEYINPUT69), .A2(new_n229), .A3(new_n202), .A4(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n216), .B(new_n220), .C1(new_n230), .C2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT71), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n229), .A2(new_n202), .A3(new_n231), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n225), .A2(KEYINPUT69), .A3(new_n229), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n240), .A2(KEYINPUT71), .A3(new_n216), .A4(new_n220), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n189), .A2(KEYINPUT25), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n216), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n220), .A2(KEYINPUT70), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n220), .A2(KEYINPUT70), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n243), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n242), .A2(KEYINPUT72), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT72), .B1(new_n242), .B2(new_n248), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n235), .A2(new_n241), .B1(new_n244), .B2(new_n247), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT25), .B1(new_n252), .B2(new_n189), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n191), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n190), .A2(G902), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n187), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n242), .A2(new_n248), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n242), .A2(KEYINPUT72), .A3(new_n248), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n190), .B1(new_n264), .B2(new_n253), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT73), .A3(new_n257), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(G472), .A2(G902), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT11), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(G137), .ZN(new_n271));
  INV_X1    g085(.A(G137), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT11), .A3(G134), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(G137), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G131), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n271), .A2(new_n273), .A3(new_n277), .A4(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G143), .B(G146), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT0), .B(G128), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n200), .A2(G143), .ZN(new_n283));
  INV_X1    g097(.A(G143), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G146), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(KEYINPUT0), .A2(G128), .ZN(new_n287));
  OR2_X1    g101(.A1(KEYINPUT0), .A2(G128), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n286), .A2(KEYINPUT64), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n279), .A2(new_n282), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT1), .B1(new_n284), .B2(G146), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n284), .A2(G146), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n200), .A2(G143), .ZN(new_n293));
  OAI211_X1 g107(.A(G128), .B(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n270), .A2(G137), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n272), .A2(G134), .ZN(new_n296));
  OAI21_X1  g110(.A(G131), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n283), .B(new_n285), .C1(KEYINPUT1), .C2(new_n204), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n294), .A2(new_n278), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n206), .A2(G116), .ZN(new_n300));
  INV_X1    g114(.A(G116), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G119), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(G113), .ZN(new_n304));
  INV_X1    g118(.A(G113), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n300), .B(new_n302), .C1(new_n304), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n300), .A2(new_n302), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT2), .B(G113), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n290), .A2(new_n299), .A3(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G237), .A2(G953), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G210), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT27), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT26), .B(G101), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n271), .A2(new_n273), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n296), .A2(G131), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n320), .A2(new_n321), .B1(new_n275), .B2(G131), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n282), .A2(new_n289), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n299), .A2(KEYINPUT30), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n311), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT30), .B1(new_n290), .B2(new_n299), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT65), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n299), .A2(KEYINPUT30), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n312), .B1(new_n329), .B2(new_n290), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT65), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n299), .B1(new_n322), .B2(new_n323), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n319), .B1(new_n328), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT67), .B(KEYINPUT31), .Z(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(new_n311), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n313), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT28), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n313), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n318), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n336), .A2(new_n337), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n319), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT65), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n331), .B1(new_n330), .B2(new_n334), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT66), .B1(new_n349), .B2(KEYINPUT31), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT66), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT31), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n336), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(KEYINPUT68), .B(new_n345), .C1(new_n350), .C2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n349), .A2(KEYINPUT66), .A3(KEYINPUT31), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n351), .B1(new_n336), .B2(new_n352), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT68), .B1(new_n358), .B2(new_n345), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n268), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT32), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G472), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n343), .A2(new_n344), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(KEYINPUT29), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n313), .B1(new_n347), .B2(new_n348), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n365), .B1(new_n318), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(G902), .B1(new_n364), .B2(KEYINPUT29), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n345), .B1(new_n350), .B2(new_n353), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT68), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n354), .ZN(new_n374));
  INV_X1    g188(.A(new_n268), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(new_n361), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n370), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n267), .B1(new_n362), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n218), .A2(G227), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(KEYINPUT74), .ZN(new_n381));
  XNOR2_X1  g195(.A(G110), .B(G140), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n381), .B(new_n382), .Z(new_n383));
  NAND2_X1  g197(.A1(new_n294), .A2(new_n298), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(new_n385), .B2(G107), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  INV_X1    g201(.A(G107), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G104), .ZN(new_n389));
  INV_X1    g203(.A(G101), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(G107), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n386), .A2(new_n389), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n385), .A2(G107), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n388), .A2(G104), .ZN(new_n394));
  OAI21_X1  g208(.A(G101), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n384), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n294), .A2(new_n298), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n392), .A2(new_n395), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT77), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT77), .B1(new_n384), .B2(new_n396), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n384), .A2(new_n396), .A3(KEYINPUT79), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n399), .A2(new_n403), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n322), .A2(KEYINPUT78), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(KEYINPUT12), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n406), .B(new_n407), .C1(KEYINPUT12), .C2(new_n409), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n386), .A2(new_n389), .A3(new_n391), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G101), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT75), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n392), .A2(KEYINPUT4), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT75), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n418), .A3(G101), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  XOR2_X1   g234(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n421));
  NAND3_X1  g235(.A1(new_n414), .A2(G101), .A3(new_n421), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n422), .A2(new_n282), .A3(new_n289), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n384), .A2(new_n396), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n420), .A2(new_n423), .B1(new_n424), .B2(KEYINPUT10), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT10), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n403), .A2(new_n426), .A3(new_n404), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n322), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n383), .B1(new_n413), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n383), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n322), .B1(new_n425), .B2(new_n427), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n379), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n430), .ZN(new_n434));
  INV_X1    g248(.A(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n428), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n412), .B2(new_n411), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n436), .B(KEYINPUT80), .C1(new_n438), .C2(new_n383), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n433), .A2(G469), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G469), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(new_n189), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n413), .A2(new_n434), .ZN(new_n443));
  INV_X1    g257(.A(new_n383), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n437), .B2(new_n431), .ZN(new_n445));
  AOI21_X1  g259(.A(G902), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n442), .B1(new_n446), .B2(new_n441), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT9), .B(G234), .ZN(new_n449));
  OAI21_X1  g263(.A(G221), .B1(new_n449), .B2(G902), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n311), .A2(new_n422), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n420), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT5), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n206), .A3(G116), .ZN(new_n456));
  OAI211_X1 g270(.A(G113), .B(new_n456), .C1(new_n308), .C2(new_n455), .ZN(new_n457));
  AND4_X1   g271(.A1(new_n307), .A2(new_n457), .A3(new_n392), .A4(new_n395), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n458), .B1(new_n420), .B2(new_n453), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n461), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(KEYINPUT6), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n282), .A2(new_n289), .A3(G125), .ZN(new_n467));
  INV_X1    g281(.A(G224), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G953), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n294), .A2(new_n196), .A3(new_n298), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n467), .B2(new_n471), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT81), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n461), .B1(new_n454), .B2(new_n459), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR4_X1   g292(.A1(new_n464), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n461), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n466), .B(new_n474), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n461), .B(KEYINPUT8), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n401), .B1(new_n307), .B2(new_n457), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(new_n458), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n467), .A2(new_n484), .A3(new_n470), .A4(new_n471), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n469), .A2(KEYINPUT7), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n472), .A2(new_n473), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(G902), .B1(new_n489), .B2(new_n465), .ZN(new_n490));
  OAI21_X1  g304(.A(G210), .B1(G237), .B2(G902), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n480), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n480), .A2(new_n490), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n491), .B(KEYINPUT82), .Z(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(G234), .A2(G237), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n497), .A2(G952), .A3(new_n218), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n497), .A2(G902), .A3(G953), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT21), .B(G898), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G214), .B1(G237), .B2(G902), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n496), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n314), .A2(G143), .A3(G214), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(G143), .B1(new_n314), .B2(G214), .ZN(new_n507));
  OAI211_X1 g321(.A(KEYINPUT18), .B(G131), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n314), .A2(G214), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n284), .ZN(new_n510));
  NAND2_X1  g324(.A1(KEYINPUT18), .A2(G131), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n223), .A2(new_n200), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n508), .B(new_n512), .C1(new_n221), .C2(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n506), .A2(new_n507), .A3(G131), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n277), .B1(new_n510), .B2(new_n505), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT17), .ZN(new_n517));
  OAI211_X1 g331(.A(KEYINPUT17), .B(G131), .C1(new_n506), .C2(new_n507), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n201), .A2(new_n518), .A3(new_n202), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n514), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(G113), .B(G122), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n521), .A2(G104), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(G104), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n520), .A2(KEYINPUT85), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT85), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n514), .B(new_n525), .C1(new_n517), .C2(new_n519), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT84), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n522), .A2(new_n528), .A3(new_n523), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n522), .B2(new_n523), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n531), .B(new_n514), .C1(new_n517), .C2(new_n519), .ZN(new_n532));
  AOI21_X1  g346(.A(G902), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G475), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT20), .ZN(new_n535));
  AND2_X1   g349(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n536));
  NOR2_X1   g350(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n223), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n538), .B(new_n200), .C1(new_n223), .C2(new_n537), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n539), .B(new_n202), .C1(new_n516), .C2(new_n515), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n514), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n522), .A2(new_n523), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n532), .ZN(new_n544));
  NOR2_X1   g358(.A1(G475), .A2(G902), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n535), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n545), .ZN(new_n547));
  AOI211_X1 g361(.A(KEYINPUT20), .B(new_n547), .C1(new_n543), .C2(new_n532), .ZN(new_n548));
  OAI22_X1  g362(.A1(new_n533), .A2(new_n534), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(G128), .B(G143), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT13), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n284), .A2(G128), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n551), .B(G134), .C1(KEYINPUT13), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n270), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n554), .A2(KEYINPUT88), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n554), .A2(KEYINPUT88), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT86), .B1(new_n301), .B2(G122), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n559));
  INV_X1    g373(.A(G122), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(G116), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT87), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n301), .A2(G122), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n563), .B1(new_n562), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n388), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n567), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(G107), .A3(new_n565), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n557), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n550), .A2(new_n270), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n554), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT89), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OR3_X1    g390(.A1(new_n564), .A2(KEYINPUT90), .A3(KEYINPUT14), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n564), .A2(KEYINPUT14), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT90), .B1(new_n564), .B2(KEYINPUT14), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n577), .A2(new_n562), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G107), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n573), .A2(KEYINPUT89), .A3(new_n554), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n568), .A2(new_n576), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n449), .A2(new_n188), .A3(G953), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n572), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n584), .ZN(new_n586));
  INV_X1    g400(.A(new_n583), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(new_n571), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G478), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT15), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR4_X1   g409(.A1(new_n451), .A2(new_n504), .A3(new_n549), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n378), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  AOI21_X1  g412(.A(G902), .B1(new_n373), .B2(new_n354), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n360), .B1(new_n599), .B2(new_n363), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n600), .A2(new_n267), .A3(new_n451), .ZN(new_n601));
  INV_X1    g415(.A(new_n549), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n585), .A2(new_n588), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT33), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n585), .A2(new_n588), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(G478), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n590), .A2(new_n189), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n589), .B2(new_n590), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n602), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n502), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n480), .A2(new_n490), .A3(new_n491), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n491), .B1(new_n480), .B2(new_n490), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n503), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n601), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G104), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  NOR2_X1   g434(.A1(new_n546), .A2(new_n548), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT92), .B1(new_n533), .B2(new_n534), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT92), .ZN(new_n623));
  INV_X1    g437(.A(new_n532), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n524), .B2(new_n526), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n623), .B(G475), .C1(new_n625), .C2(G902), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n621), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n502), .A3(new_n595), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT93), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n630), .A2(new_n631), .A3(new_n615), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n601), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  INV_X1    g449(.A(new_n600), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT36), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n638), .B1(new_n245), .B2(new_n246), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT94), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT94), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n641), .B(new_n638), .C1(new_n245), .C2(new_n246), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n244), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n640), .A2(new_n240), .A3(new_n216), .A4(new_n642), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n256), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n637), .B1(new_n255), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n646), .B(KEYINPUT95), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n265), .A2(KEYINPUT96), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n596), .A2(new_n636), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT37), .B(G110), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT97), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n653), .B(new_n655), .ZN(G12));
  OAI21_X1  g470(.A(new_n376), .B1(new_n355), .B2(new_n359), .ZN(new_n657));
  INV_X1    g471(.A(new_n370), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n375), .B1(new_n373), .B2(new_n354), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n657), .B(new_n658), .C1(new_n659), .C2(KEYINPUT32), .ZN(new_n660));
  INV_X1    g474(.A(new_n450), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n440), .B2(new_n447), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n662), .A2(new_n649), .A3(new_n651), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n498), .B1(new_n499), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n627), .A2(new_n595), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n615), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n660), .A2(new_n663), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  XNOR2_X1  g484(.A(new_n496), .B(KEYINPUT38), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n265), .A2(new_n650), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n595), .A2(new_n549), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  AND4_X1   g489(.A1(new_n503), .A2(new_n671), .A3(new_n673), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n366), .A2(new_n318), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n344), .A2(new_n338), .A3(new_n313), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n677), .A2(KEYINPUT98), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n189), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT98), .B1(new_n677), .B2(new_n678), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n362), .A2(new_n657), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n665), .B(KEYINPUT39), .Z(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n451), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n689), .A2(KEYINPUT40), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(KEYINPUT40), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n676), .A2(KEYINPUT99), .A3(new_n683), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n686), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  NAND4_X1  g509(.A1(new_n549), .A2(new_n607), .A3(new_n609), .A4(new_n666), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT100), .B1(new_n615), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n503), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n480), .A2(new_n490), .ZN(new_n699));
  INV_X1    g513(.A(new_n491), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n698), .B1(new_n701), .B2(new_n492), .ZN(new_n702));
  AND4_X1   g516(.A1(new_n549), .A2(new_n607), .A3(new_n609), .A4(new_n666), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT100), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n660), .A2(new_n663), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  AND2_X1   g522(.A1(new_n259), .A2(new_n266), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n430), .B1(new_n412), .B2(new_n411), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n383), .B1(new_n435), .B2(new_n428), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n189), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G469), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n441), .B(new_n189), .C1(new_n710), .C2(new_n711), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n450), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n660), .A2(new_n616), .A3(new_n709), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT101), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND3_X1  g534(.A1(new_n632), .A2(new_n378), .A3(new_n716), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  NOR2_X1   g536(.A1(new_n715), .A2(new_n615), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n595), .A2(new_n501), .A3(new_n549), .ZN(new_n724));
  AND4_X1   g538(.A1(new_n649), .A2(new_n723), .A3(new_n651), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n660), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  OAI21_X1  g541(.A(KEYINPUT103), .B1(new_n599), .B2(new_n363), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n189), .B1(new_n355), .B2(new_n359), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n730), .A3(G472), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n255), .A2(new_n258), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n268), .B(KEYINPUT102), .Z(new_n734));
  INV_X1    g548(.A(new_n345), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n336), .A2(new_n352), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR4_X1   g551(.A1(new_n715), .A2(new_n615), .A3(new_n674), .A4(new_n501), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n732), .A2(new_n733), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  INV_X1    g554(.A(new_n723), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n696), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n732), .A2(new_n672), .A3(new_n742), .A4(new_n737), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT104), .B(G125), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G27));
  NAND2_X1  g559(.A1(new_n660), .A2(new_n733), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n496), .A2(new_n698), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n703), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n436), .B(G469), .C1(new_n438), .C2(new_n383), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n442), .B(KEYINPUT105), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n714), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n753), .A2(KEYINPUT106), .A3(new_n450), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT106), .B1(new_n753), .B2(new_n450), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n750), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n495), .B1(new_n480), .B2(new_n490), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n613), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n503), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n754), .A2(new_n755), .A3(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n660), .A2(new_n760), .A3(new_n709), .A4(new_n703), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n748), .A2(new_n756), .B1(new_n747), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n277), .ZN(G33));
  INV_X1    g577(.A(new_n667), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n378), .A2(new_n764), .A3(new_n760), .ZN(new_n765));
  XOR2_X1   g579(.A(KEYINPUT107), .B(G134), .Z(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G36));
  AOI21_X1  g581(.A(KEYINPUT45), .B1(new_n433), .B2(new_n439), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n436), .B1(new_n438), .B2(new_n383), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  OAI21_X1  g584(.A(G469), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(KEYINPUT46), .B(new_n752), .C1(new_n768), .C2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT108), .A3(new_n714), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n768), .A2(new_n771), .ZN(new_n774));
  INV_X1    g588(.A(new_n752), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n773), .B1(new_n776), .B2(KEYINPUT46), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT108), .B1(new_n772), .B2(new_n714), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n450), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n779), .A2(new_n688), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n610), .A2(KEYINPUT43), .A3(new_n549), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT43), .B1(new_n610), .B2(new_n549), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n673), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(KEYINPUT44), .A3(new_n600), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n749), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT109), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n785), .A2(new_n600), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n781), .B(new_n788), .C1(KEYINPUT44), .C2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  XNOR2_X1  g605(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n779), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n779), .A2(new_n793), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n660), .A2(new_n709), .A3(new_n750), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  NAND3_X1  g613(.A1(new_n733), .A2(new_n450), .A3(new_n503), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT111), .Z(new_n801));
  AND2_X1   g615(.A1(new_n713), .A2(new_n714), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n804), .A2(new_n549), .A3(new_n610), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(new_n803), .B2(new_n802), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n801), .A2(new_n806), .A3(new_n683), .A4(new_n671), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT112), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n660), .B(new_n663), .C1(new_n668), .C2(new_n706), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n675), .A2(new_n702), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n753), .A2(new_n450), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n672), .A2(new_n813), .A3(new_n665), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n659), .A2(KEYINPUT32), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n657), .A2(new_n682), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n812), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(new_n818), .B2(new_n743), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n743), .A2(KEYINPUT52), .A3(new_n810), .A4(new_n817), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n809), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  INV_X1    g637(.A(new_n743), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n810), .A2(new_n817), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(KEYINPUT116), .A3(new_n820), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n765), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n732), .A2(new_n756), .A3(new_n672), .A4(new_n737), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n595), .A2(new_n665), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n749), .A2(new_n627), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n660), .A2(new_n663), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n762), .A2(new_n829), .A3(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n378), .A2(new_n596), .B1(new_n725), .B2(new_n660), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n612), .A2(new_n698), .A3(new_n758), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n601), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n836), .A2(new_n838), .A3(new_n721), .A4(new_n739), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT101), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n717), .B(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n267), .A2(new_n451), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n595), .A2(new_n602), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n504), .A2(KEYINPUT113), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT113), .B1(new_n504), .B2(new_n844), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n636), .A2(new_n843), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT114), .B1(new_n847), .B2(new_n653), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n847), .A2(new_n653), .A3(KEYINPUT114), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n835), .A2(new_n842), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n828), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n835), .A2(new_n842), .A3(new_n851), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n820), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n826), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n856), .B(new_n823), .C1(new_n824), .C2(new_n825), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT53), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT54), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n853), .B1(new_n828), .B2(new_n852), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n842), .A2(new_n851), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n860), .A3(KEYINPUT53), .A4(new_n835), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n862), .B1(KEYINPUT54), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n749), .A2(new_n716), .A3(new_n498), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n709), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n683), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n602), .A3(new_n610), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n732), .A2(new_n737), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n672), .ZN(new_n873));
  INV_X1    g687(.A(new_n784), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n871), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n872), .A2(new_n733), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n874), .A2(new_n498), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n759), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n802), .A2(new_n661), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n794), .A2(new_n795), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n876), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n671), .A2(new_n503), .A3(new_n715), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n872), .A2(new_n733), .A3(new_n878), .A4(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT50), .B1(new_n885), .B2(KEYINPUT117), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n885), .A2(KEYINPUT117), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n877), .A2(KEYINPUT50), .A3(new_n878), .A4(new_n884), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n886), .A2(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n887), .A2(new_n889), .A3(new_n886), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n883), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(KEYINPUT51), .B(new_n883), .C1(new_n890), .C2(new_n891), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n879), .A2(new_n741), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n746), .A2(new_n875), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n897), .A2(KEYINPUT119), .A3(KEYINPUT48), .ZN(new_n898));
  XOR2_X1   g712(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n870), .A2(new_n611), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n901), .A3(G952), .A4(new_n218), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n896), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n894), .A2(new_n895), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n867), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n808), .B1(new_n905), .B2(new_n906), .ZN(G75));
  NOR2_X1   g721(.A1(new_n218), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n189), .B1(new_n863), .B2(new_n865), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT56), .B1(new_n910), .B2(G210), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n466), .B1(new_n478), .B2(new_n479), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n474), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n909), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT56), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n910), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(new_n495), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(KEYINPUT120), .B(new_n917), .C1(new_n918), .C2(new_n495), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n915), .B1(new_n921), .B2(new_n922), .ZN(G51));
  XOR2_X1   g737(.A(new_n752), .B(KEYINPUT57), .Z(new_n924));
  NOR2_X1   g738(.A1(new_n866), .A2(KEYINPUT54), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n863), .B2(new_n865), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n924), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n443), .A2(new_n445), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n910), .A2(new_n774), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n908), .B1(new_n930), .B2(new_n931), .ZN(G54));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n933));
  AND2_X1   g747(.A1(KEYINPUT58), .A2(G475), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n910), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n544), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n908), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n910), .A2(KEYINPUT121), .A3(new_n544), .A4(new_n934), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(G60));
  NAND2_X1  g754(.A1(new_n604), .A2(new_n606), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT122), .Z(new_n942));
  XOR2_X1   g756(.A(new_n608), .B(KEYINPUT59), .Z(new_n943));
  OAI211_X1 g757(.A(new_n942), .B(new_n943), .C1(new_n925), .C2(new_n927), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n909), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n942), .B1(new_n867), .B2(new_n943), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(G63));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT123), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT60), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n863), .B2(new_n865), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n645), .A3(new_n644), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n909), .B1(new_n953), .B2(new_n252), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n948), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n953), .A2(new_n252), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n958), .A2(KEYINPUT61), .A3(new_n909), .A4(new_n954), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(G66));
  OAI21_X1  g774(.A(G953), .B1(new_n500), .B2(new_n468), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n864), .B2(G953), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n912), .B1(G898), .B2(new_n218), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT124), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n962), .B(new_n964), .ZN(G69));
  OAI21_X1  g779(.A(new_n334), .B1(new_n324), .B2(new_n325), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n538), .B1(new_n223), .B2(new_n537), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n844), .B1(new_n602), .B2(new_n610), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT125), .Z(new_n970));
  AND4_X1   g784(.A1(new_n378), .A2(new_n970), .A3(new_n689), .A4(new_n749), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n743), .A2(new_n810), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n694), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n694), .A2(KEYINPUT62), .A3(new_n973), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n971), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n790), .A3(new_n798), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n968), .B1(new_n979), .B2(new_n218), .ZN(new_n980));
  OR3_X1    g794(.A1(new_n780), .A2(new_n746), .A3(new_n811), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n762), .A2(new_n829), .A3(new_n972), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n790), .A2(new_n981), .A3(new_n798), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n983), .A2(G953), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n968), .B1(new_n664), .B2(new_n218), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n980), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(G227), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n988), .B2(new_n664), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n987), .B(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  INV_X1    g806(.A(new_n864), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n992), .B1(new_n983), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n366), .A2(new_n318), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT126), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n978), .A2(new_n790), .A3(new_n798), .A4(new_n864), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n998), .A2(new_n992), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n909), .B(new_n997), .C1(new_n999), .C2(new_n677), .ZN(new_n1000));
  OR2_X1    g814(.A1(new_n854), .A2(new_n861), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n677), .A2(new_n992), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1003), .A2(new_n995), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(KEYINPUT127), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1000), .B1(new_n1005), .B2(new_n1007), .ZN(G57));
endmodule


