//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1307, new_n1308, new_n1309,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT64), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(KEYINPUT64), .A2(G20), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AND2_X1   g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI22_X1  g0021(.A1(new_n203), .A2(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n222), .B1(new_n228), .B2(KEYINPUT66), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT65), .Z(new_n231));
  OAI211_X1 g0031(.A(new_n229), .B(new_n231), .C1(KEYINPUT66), .C2(new_n228), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(new_n207), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n210), .B1(new_n217), .B2(new_n218), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT68), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n240), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT69), .ZN(new_n247));
  XOR2_X1   g0047(.A(G58), .B(G77), .Z(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT70), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n249), .B(new_n253), .Z(G351));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n216), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(G226), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n256), .A2(G274), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n256), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  OAI211_X1 g0068(.A(G222), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n268), .ZN(new_n270));
  NAND2_X1  g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G77), .A3(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(G223), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n269), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n264), .B1(new_n265), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G169), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT8), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G58), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n281), .A3(KEYINPUT71), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT64), .A2(G20), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT64), .A2(G20), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT71), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n282), .A2(G33), .A3(new_n285), .A4(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G1), .A2(G13), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n292), .A2(new_n293), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(KEYINPUT72), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT72), .ZN(new_n299));
  INV_X1    g0099(.A(new_n297), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n294), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT73), .B1(new_n212), .B2(G1), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT73), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(new_n257), .A3(G20), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G50), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n297), .A2(G50), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n295), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n275), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n278), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n267), .A2(new_n268), .ZN(new_n316));
  INV_X1    g0116(.A(G107), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n256), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(G232), .A2(G1698), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n219), .B2(G1698), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n318), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n256), .A2(new_n258), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G244), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(new_n263), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G190), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n306), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n220), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n297), .A2(new_n293), .A3(new_n292), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n329), .A2(new_n330), .B1(new_n220), .B2(new_n300), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n285), .A2(G33), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT15), .B(G87), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n279), .A2(new_n281), .ZN(new_n335));
  INV_X1    g0135(.A(new_n289), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n335), .A2(new_n336), .B1(new_n285), .B2(new_n220), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n294), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n327), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n325), .A2(G200), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n325), .A2(new_n277), .B1(new_n331), .B2(new_n338), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n325), .A2(G179), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n340), .A2(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n312), .A2(KEYINPUT9), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n296), .B1(new_n288), .B2(new_n290), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(new_n310), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT9), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n348), .A3(new_n309), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G200), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n275), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n274), .A2(new_n265), .ZN(new_n353));
  INV_X1    g0153(.A(new_n264), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n354), .A3(G190), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT74), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT74), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n275), .A2(new_n357), .A3(G190), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n352), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT10), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n350), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(new_n350), .B2(new_n359), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n315), .B(new_n344), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT75), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n348), .B1(new_n347), .B2(new_n309), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n307), .B1(new_n301), .B2(new_n298), .ZN(new_n367));
  NOR4_X1   g0167(.A1(new_n346), .A2(new_n367), .A3(KEYINPUT9), .A4(new_n310), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n276), .A2(G200), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n355), .A2(KEYINPUT74), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n357), .B1(new_n275), .B2(G190), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT10), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n350), .A2(new_n359), .A3(new_n360), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n376), .A2(KEYINPUT75), .A3(new_n315), .A4(new_n344), .ZN(new_n377));
  INV_X1    g0177(.A(G226), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n266), .ZN(new_n379));
  INV_X1    g0179(.A(G232), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G1698), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n379), .B(new_n381), .C1(new_n267), .C2(new_n268), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT76), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT76), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n382), .A2(new_n386), .A3(new_n383), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n265), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n263), .B1(new_n322), .B2(new_n219), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT13), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n256), .B1(new_n384), .B2(KEYINPUT76), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n389), .B1(new_n393), .B2(new_n387), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT13), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT14), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n398), .A3(G169), .ZN(new_n399));
  AOI211_X1 g0199(.A(KEYINPUT13), .B(new_n389), .C1(new_n393), .C2(new_n387), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n395), .B1(new_n388), .B2(new_n390), .ZN(new_n401));
  OAI21_X1  g0201(.A(G169), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT14), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n400), .A2(new_n313), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT77), .B1(new_n394), .B2(new_n395), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT77), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n399), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n289), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n332), .B2(new_n220), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n294), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT11), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(KEYINPUT11), .A3(new_n294), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n328), .A2(new_n203), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT12), .B1(new_n297), .B2(G68), .ZN(new_n417));
  OR3_X1    g0217(.A1(new_n297), .A2(KEYINPUT12), .A3(G68), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n416), .A2(new_n330), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n407), .A2(new_n405), .A3(G190), .A4(new_n396), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n420), .B1(new_n397), .B2(G200), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n409), .A2(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(G58), .B(G68), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(G20), .B1(G159), .B2(new_n289), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n267), .A2(new_n268), .A3(G20), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT7), .ZN(new_n427));
  OAI21_X1  g0227(.A(G68), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT3), .B(G33), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n215), .A2(new_n429), .A3(KEYINPUT7), .ZN(new_n430));
  OAI211_X1 g0230(.A(KEYINPUT16), .B(new_n425), .C1(new_n428), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n294), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT7), .B1(new_n215), .B2(new_n429), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n316), .A2(new_n427), .A3(new_n212), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(G68), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT16), .B1(new_n435), .B2(new_n425), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT78), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n306), .A2(new_n282), .A3(new_n287), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n301), .B2(new_n298), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n282), .A2(new_n287), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n300), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n438), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n439), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n302), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(KEYINPUT78), .A3(new_n442), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n437), .A2(new_n448), .ZN(new_n449));
  OR2_X1    g0249(.A1(G223), .A2(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n378), .A2(G1698), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n450), .B(new_n451), .C1(new_n267), .C2(new_n268), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G87), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n265), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n256), .A2(G232), .A3(new_n258), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n263), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n457), .A3(G179), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n256), .B1(new_n452), .B2(new_n453), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n263), .A2(new_n456), .ZN(new_n460));
  OAI21_X1  g0260(.A(G169), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT79), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n458), .A2(new_n461), .A3(KEYINPUT79), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT18), .B1(new_n449), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT17), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n444), .B(new_n447), .C1(new_n432), .C2(new_n436), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n459), .A2(new_n460), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n326), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(G200), .B2(new_n470), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n468), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n448), .ZN(new_n475));
  OR2_X1    g0275(.A1(new_n432), .A2(new_n436), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT17), .A4(new_n472), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n458), .A2(KEYINPUT79), .A3(new_n461), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT79), .B1(new_n458), .B2(new_n461), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT18), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(new_n469), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n467), .A2(new_n474), .A3(new_n477), .A4(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n365), .A2(new_n377), .A3(new_n423), .A4(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT21), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT85), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G33), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G97), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  AND4_X1   g0294(.A1(new_n213), .A2(new_n493), .A3(new_n214), .A4(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G116), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G20), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n488), .A2(new_n489), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n294), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n491), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n498), .A2(new_n497), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n213), .A2(new_n493), .A3(new_n214), .A4(new_n494), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(new_n294), .A4(new_n490), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n257), .A2(G33), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n330), .A2(KEYINPUT84), .A3(G116), .A4(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT84), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n297), .A2(new_n505), .A3(new_n293), .A4(new_n292), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n496), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n497), .ZN(new_n511));
  INV_X1    g0311(.A(G13), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(G1), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n504), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n261), .A2(G1), .ZN(new_n516));
  AND2_X1   g0316(.A1(KEYINPUT5), .A2(G41), .ZN(new_n517));
  NOR2_X1   g0317(.A1(KEYINPUT5), .A2(G41), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(G270), .A3(new_n256), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n266), .A2(G264), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G257), .A2(G1698), .ZN(new_n522));
  OAI22_X1  g0322(.A1(new_n521), .A2(new_n522), .B1(new_n267), .B2(new_n268), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n523), .B(new_n265), .C1(G303), .C2(new_n429), .ZN(new_n524));
  AND2_X1   g0324(.A1(G33), .A2(G41), .ZN(new_n525));
  OAI21_X1  g0325(.A(G274), .B1(new_n525), .B2(new_n293), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT81), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n519), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n257), .A2(G45), .ZN(new_n529));
  OR2_X1    g0329(.A1(KEYINPUT5), .A2(G41), .ZN(new_n530));
  NAND2_X1  g0330(.A1(KEYINPUT5), .A2(G41), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G274), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n216), .B2(new_n255), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT81), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n520), .B(new_n524), .C1(new_n528), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G169), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n487), .B1(new_n515), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n504), .A2(new_n510), .A3(new_n514), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n487), .A2(new_n277), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n527), .B1(new_n519), .B2(new_n526), .ZN(new_n542));
  XNOR2_X1  g0342(.A(KEYINPUT5), .B(G41), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n534), .A2(KEYINPUT81), .A3(new_n543), .A4(new_n516), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n543), .A2(new_n516), .B1(new_n216), .B2(new_n255), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n542), .A2(new_n544), .B1(new_n545), .B2(G270), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n541), .B1(new_n546), .B2(new_n524), .ZN(new_n547));
  INV_X1    g0347(.A(G303), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n256), .B1(new_n316), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n313), .B1(new_n549), .B2(new_n523), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n542), .A2(new_n544), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n550), .A2(new_n551), .A3(new_n520), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n539), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n538), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n536), .A2(G200), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n515), .B(new_n555), .C1(new_n326), .C2(new_n536), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT86), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n536), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n539), .B1(new_n559), .B2(G190), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(KEYINPUT86), .A3(new_n555), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n554), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(KEYINPUT23), .A2(G107), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n283), .B2(new_n284), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G116), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT23), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n212), .ZN(new_n568));
  NAND2_X1  g0368(.A1(KEYINPUT23), .A2(G107), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n213), .B(new_n214), .C1(new_n267), .C2(new_n268), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT22), .B1(new_n571), .B2(new_n224), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n285), .A2(new_n429), .A3(new_n573), .A4(G87), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT24), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI211_X1 g0377(.A(KEYINPUT24), .B(new_n570), .C1(new_n572), .C2(new_n574), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n294), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n551), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n519), .A2(G264), .A3(new_n256), .ZN(new_n581));
  NOR2_X1   g0381(.A1(G250), .A2(G1698), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n227), .B2(G1698), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(new_n429), .B1(G33), .B2(G294), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n581), .B1(new_n584), .B2(new_n256), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n351), .B1(new_n580), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n227), .A2(G1698), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G250), .B2(G1698), .ZN(new_n588));
  INV_X1    g0388(.A(G294), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n588), .A2(new_n316), .B1(new_n492), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(new_n265), .B1(new_n545), .B2(G264), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(new_n326), .A3(new_n551), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT80), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n330), .A2(new_n594), .A3(new_n505), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n508), .A2(KEYINPUT80), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(G107), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n297), .A2(G107), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n598), .B(KEYINPUT25), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n579), .A2(new_n593), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n277), .B1(new_n580), .B2(new_n585), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n591), .A2(new_n313), .A3(new_n551), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n579), .B2(new_n600), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT6), .ZN(new_n607));
  AND2_X1   g0407(.A1(G97), .A2(G107), .ZN(new_n608));
  NOR2_X1   g0408(.A1(G97), .A2(G107), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n317), .A2(KEYINPUT6), .A3(G97), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(new_n215), .B1(G77), .B2(new_n289), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n433), .A2(G107), .A3(new_n434), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n296), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n595), .A2(G97), .A3(new_n596), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n297), .A2(G97), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(G244), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT4), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n429), .A2(KEYINPUT4), .A3(G244), .A4(new_n266), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n429), .A2(G250), .A3(G1698), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n494), .A4(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n265), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n542), .A2(new_n544), .B1(new_n545), .B2(G257), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n625), .A2(new_n326), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(G200), .B1(new_n625), .B2(new_n626), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n618), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n613), .A2(new_n614), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n294), .ZN(new_n631));
  INV_X1    g0431(.A(new_n616), .ZN(new_n632));
  INV_X1    g0432(.A(new_n617), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n625), .A2(new_n626), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n277), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n625), .A2(new_n313), .A3(new_n626), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n213), .A2(G33), .A3(G97), .A4(new_n214), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT19), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n213), .A2(new_n214), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT83), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n224), .ZN(new_n645));
  NAND2_X1  g0445(.A1(KEYINPUT83), .A2(G87), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n609), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n285), .A2(new_n429), .A3(G68), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n641), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n294), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n333), .A2(new_n300), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n595), .A2(G87), .A3(new_n596), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OAI22_X1  g0454(.A1(KEYINPUT82), .A2(new_n225), .B1(new_n261), .B2(G1), .ZN(new_n655));
  NAND2_X1  g0455(.A1(KEYINPUT82), .A2(G250), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n656), .A2(new_n257), .A3(G45), .A4(new_n533), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n256), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n565), .ZN(new_n659));
  NOR2_X1   g0459(.A1(G238), .A2(G1698), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n221), .B2(G1698), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n659), .B1(new_n661), .B2(new_n429), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n326), .B(new_n658), .C1(new_n662), .C2(new_n256), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n219), .A2(new_n266), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n221), .A2(G1698), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n664), .B(new_n665), .C1(new_n267), .C2(new_n268), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n256), .B1(new_n666), .B2(new_n565), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n655), .A2(new_n256), .A3(new_n657), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n663), .B1(new_n669), .B2(G200), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n277), .B1(new_n667), .B2(new_n668), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n313), .B(new_n658), .C1(new_n662), .C2(new_n256), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n333), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n595), .A2(new_n674), .A3(new_n596), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n651), .A2(new_n652), .A3(new_n675), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n654), .A2(new_n670), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n629), .A2(new_n638), .A3(new_n677), .ZN(new_n678));
  AND4_X1   g0478(.A1(new_n486), .A2(new_n562), .A3(new_n606), .A4(new_n678), .ZN(G372));
  INV_X1    g0479(.A(KEYINPUT88), .ZN(new_n680));
  INV_X1    g0480(.A(new_n376), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n474), .A2(new_n477), .ZN(new_n682));
  INV_X1    g0482(.A(new_n420), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n406), .B1(new_n391), .B2(KEYINPUT13), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n394), .A2(KEYINPUT77), .A3(new_n395), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n686), .A2(new_n404), .B1(KEYINPUT14), .B2(new_n402), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n683), .B1(new_n687), .B2(new_n399), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n342), .A2(new_n343), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n422), .B2(new_n421), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n682), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n469), .A2(new_n462), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(new_n481), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n681), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n315), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n680), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n693), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n409), .A2(new_n420), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n422), .A2(new_n421), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n689), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n697), .B1(new_n700), .B2(new_n682), .ZN(new_n701));
  OAI211_X1 g0501(.A(KEYINPUT88), .B(new_n315), .C1(new_n701), .C2(new_n681), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT26), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n673), .A2(new_n676), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n650), .A2(new_n294), .B1(new_n300), .B2(new_n333), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n670), .A2(new_n706), .A3(new_n653), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n704), .B1(new_n638), .B2(new_n708), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n625), .A2(new_n313), .A3(new_n626), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n618), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(new_n677), .A3(KEYINPUT26), .A4(new_n636), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n536), .A2(new_n540), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n546), .A2(new_n550), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n500), .A2(new_n503), .B1(new_n513), .B2(new_n511), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n714), .A2(new_n715), .B1(new_n510), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n277), .B1(new_n546), .B2(new_n524), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT21), .B1(new_n718), .B2(new_n539), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT87), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT87), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n538), .A2(new_n721), .A3(new_n553), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n605), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n579), .A2(new_n593), .A3(new_n600), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n629), .A3(new_n638), .A4(new_n677), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n713), .B(new_n705), .C1(new_n723), .C2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n703), .B1(new_n485), .B2(new_n727), .ZN(G369));
  NAND2_X1  g0528(.A1(new_n285), .A2(new_n513), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n729), .A2(KEYINPUT27), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(KEYINPUT27), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(G213), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G343), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n515), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n720), .A2(new_n722), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n562), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n737), .B1(new_n738), .B2(new_n736), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n579), .A2(new_n600), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n606), .B1(new_n741), .B2(new_n735), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n605), .A2(new_n734), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n717), .A2(new_n719), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n734), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n606), .A2(new_n749), .B1(new_n605), .B2(new_n735), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n747), .A2(new_n750), .ZN(G399));
  INV_X1    g0551(.A(new_n208), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G41), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n647), .A2(G116), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n754), .A2(G1), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(new_n218), .B2(new_n754), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT28), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n713), .A2(new_n705), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n605), .A2(new_n554), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n725), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n735), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT29), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT29), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n726), .A2(new_n764), .A3(new_n735), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT30), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n546), .A2(new_n591), .A3(new_n550), .A4(new_n669), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n767), .B1(new_n768), .B2(new_n635), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(KEYINPUT89), .ZN(new_n770));
  OR3_X1    g0570(.A1(new_n768), .A2(new_n635), .A3(new_n767), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT89), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n772), .B(new_n767), .C1(new_n768), .C2(new_n635), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n591), .A2(new_n551), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n669), .A2(G179), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n635), .A2(new_n536), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n770), .A2(new_n771), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n734), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT31), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n562), .A2(new_n678), .A3(new_n606), .A4(new_n735), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n771), .A2(new_n769), .A3(new_n776), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n782), .A2(KEYINPUT31), .A3(new_n734), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G330), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n766), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n758), .B1(new_n787), .B2(G1), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT90), .Z(G364));
  NOR2_X1   g0589(.A1(new_n215), .A2(new_n512), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G45), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(new_n754), .A3(G1), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT91), .ZN(new_n794));
  OR2_X1    g0594(.A1(G355), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(G355), .A2(new_n794), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n795), .A2(new_n208), .A3(new_n429), .A4(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(G116), .B2(new_n208), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n249), .A2(G45), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n752), .A2(new_n429), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n218), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(new_n261), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n798), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n216), .B1(new_n212), .B2(G169), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT92), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(KEYINPUT92), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n793), .B1(new_n804), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n285), .A2(new_n313), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n351), .A2(G190), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(KEYINPUT33), .B(G317), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G190), .A2(G200), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n215), .A2(new_n313), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n818), .A2(new_n819), .B1(G329), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n215), .A2(new_n313), .A3(new_n816), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n326), .A2(G200), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n215), .B1(new_n827), .B2(G179), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n823), .B1(new_n824), .B2(new_n825), .C1(new_n589), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n326), .A2(new_n351), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n831), .A2(G20), .A3(new_n313), .ZN(new_n832));
  INV_X1    g0632(.A(new_n815), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n827), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G322), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n316), .B1(new_n548), .B2(new_n832), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G311), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n815), .A2(new_n820), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n815), .A2(new_n831), .ZN(new_n840));
  XOR2_X1   g0640(.A(KEYINPUT94), .B(G326), .Z(new_n841));
  OAI22_X1  g0641(.A1(new_n838), .A2(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OR3_X1    g0642(.A1(new_n830), .A2(new_n837), .A3(new_n842), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n829), .A2(KEYINPUT93), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n829), .A2(KEYINPUT93), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(G97), .ZN(new_n848));
  INV_X1    g0648(.A(G159), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT32), .B1(new_n821), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n645), .A2(new_n646), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n429), .B1(new_n852), .B2(new_n832), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n821), .A2(KEYINPUT32), .A3(new_n849), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n853), .B(new_n854), .C1(G58), .C2(new_n834), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n201), .A2(new_n840), .B1(new_n817), .B2(new_n203), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n839), .A2(new_n220), .B1(new_n317), .B2(new_n825), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n848), .A2(new_n850), .A3(new_n855), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n843), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n814), .B1(new_n860), .B2(new_n808), .ZN(new_n861));
  INV_X1    g0661(.A(new_n811), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n861), .B1(new_n739), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n740), .A2(new_n792), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n739), .A2(G330), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT95), .ZN(G396));
  NAND2_X1  g0667(.A1(new_n344), .A2(new_n735), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n726), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT97), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT97), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n726), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n342), .A2(new_n735), .A3(new_n343), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n340), .A2(new_n341), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n734), .A2(new_n339), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n876), .B1(new_n879), .B2(new_n689), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n727), .B2(new_n734), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n786), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n874), .A2(new_n785), .A3(new_n882), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(new_n792), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT98), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n825), .A2(new_n203), .B1(new_n201), .B2(new_n832), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n834), .A2(G143), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n818), .A2(G150), .ZN(new_n890));
  INV_X1    g0690(.A(new_n839), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(G159), .ZN(new_n892));
  INV_X1    g0692(.A(new_n840), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(G137), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n889), .A2(new_n890), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n896), .A2(KEYINPUT34), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n888), .B(new_n897), .C1(G58), .C2(new_n828), .ZN(new_n898));
  INV_X1    g0698(.A(G132), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n429), .B1(new_n821), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT96), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n896), .B2(KEYINPUT34), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n835), .A2(new_n589), .B1(new_n496), .B2(new_n839), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n316), .B1(new_n832), .B2(new_n317), .ZN(new_n904));
  INV_X1    g0704(.A(new_n825), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(G87), .B2(new_n905), .ZN(new_n906));
  OAI221_X1 g0706(.A(new_n906), .B1(new_n824), .B2(new_n817), .C1(new_n548), .C2(new_n840), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n903), .B(new_n907), .C1(G311), .C2(new_n822), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n898), .A2(new_n902), .B1(new_n848), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n808), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n810), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n909), .A2(new_n910), .B1(G77), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n880), .A2(new_n810), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n793), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n886), .A2(new_n887), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n887), .B1(new_n886), .B2(new_n914), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(G384));
  AOI211_X1 g0718(.A(new_n496), .B(new_n217), .C1(KEYINPUT35), .C2(new_n612), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(KEYINPUT35), .B2(new_n612), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT36), .ZN(new_n921));
  OAI21_X1  g0721(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n922), .A2(new_n218), .B1(G50), .B2(new_n203), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(G1), .A3(new_n512), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT99), .Z(new_n926));
  NAND2_X1  g0726(.A1(new_n420), .A2(new_n734), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n423), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n420), .B(new_n734), .C1(new_n699), .C2(new_n409), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n424), .A2(G20), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n289), .A2(G159), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n270), .A2(new_n212), .A3(new_n271), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n203), .B1(new_n934), .B2(KEYINPUT7), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n285), .A2(new_n316), .A3(new_n427), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n296), .B1(new_n937), .B2(KEYINPUT16), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(KEYINPUT16), .B2(new_n937), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n475), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n462), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n449), .A2(new_n472), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n732), .B1(new_n475), .B2(new_n939), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT37), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT37), .B1(new_n449), .B2(new_n472), .ZN(new_n946));
  INV_X1    g0746(.A(new_n732), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n469), .B1(new_n480), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n483), .A2(KEYINPUT101), .A3(new_n944), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT101), .B1(new_n483), .B2(new_n944), .ZN(new_n952));
  OAI211_X1 g0752(.A(KEYINPUT38), .B(new_n950), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT38), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n605), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n717), .A2(new_n719), .A3(KEYINPUT87), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n721), .B1(new_n538), .B2(new_n553), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AND4_X1   g0760(.A1(new_n724), .A2(new_n629), .A3(new_n638), .A4(new_n677), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n709), .A2(new_n712), .B1(new_n676), .B2(new_n673), .ZN(new_n963));
  AOI211_X1 g0763(.A(KEYINPUT97), .B(new_n868), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n872), .B1(new_n726), .B2(new_n869), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n875), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT100), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(KEYINPUT100), .B(new_n875), .C1(new_n964), .C2(new_n965), .ZN(new_n969));
  AOI221_X4 g0769(.A(new_n930), .B1(new_n953), .B2(new_n956), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n956), .A2(KEYINPUT39), .A3(new_n953), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n449), .A2(KEYINPUT102), .A3(new_n472), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT102), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n469), .B2(new_n473), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n469), .A2(new_n947), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n972), .A2(new_n974), .A3(new_n692), .A4(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n976), .A2(KEYINPUT37), .B1(new_n946), .B2(new_n948), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n975), .B1(new_n693), .B2(new_n682), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n955), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n953), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT39), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n698), .A2(new_n734), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n971), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n697), .A2(new_n732), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n970), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(KEYINPUT103), .B1(new_n766), .B2(new_n486), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT103), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n989), .B(new_n485), .C1(new_n763), .C2(new_n765), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n703), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n987), .B(new_n991), .Z(new_n992));
  NAND2_X1  g0792(.A1(new_n956), .A2(new_n953), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n928), .A2(new_n929), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n777), .A2(KEYINPUT31), .A3(new_n734), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n780), .A2(new_n781), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n994), .A2(new_n880), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT40), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n953), .A2(new_n979), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n994), .A2(new_n996), .A3(KEYINPUT40), .A4(new_n880), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n486), .A2(new_n996), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1005), .A2(G330), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n992), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n257), .B2(new_n790), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n992), .A2(new_n1007), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n926), .B1(new_n1009), .B2(new_n1010), .ZN(G367));
  NOR2_X1   g0811(.A1(new_n735), .A2(new_n654), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1012), .A2(new_n676), .A3(new_n673), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n708), .B2(new_n1012), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT43), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT106), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n629), .B(new_n638), .C1(new_n618), .C2(new_n735), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n711), .A2(new_n636), .A3(new_n734), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1019), .A2(new_n606), .A3(new_n749), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT105), .Z(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(KEYINPUT42), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n638), .B1(new_n1017), .B2(new_n957), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n735), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1021), .A2(KEYINPUT42), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1016), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n746), .A2(new_n1019), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT104), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1030), .A2(KEYINPUT43), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(KEYINPUT43), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1014), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1029), .B(new_n1033), .Z(new_n1034));
  XOR2_X1   g0834(.A(new_n753), .B(KEYINPUT41), .Z(new_n1035));
  NAND2_X1  g0835(.A1(new_n750), .A2(new_n1019), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT45), .Z(new_n1037));
  NOR2_X1   g0837(.A1(new_n750), .A2(new_n1019), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT44), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(new_n747), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n606), .A2(new_n749), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n744), .B2(new_n749), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(new_n740), .Z(new_n1044));
  NAND3_X1  g0844(.A1(new_n1041), .A2(new_n787), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1035), .B1(new_n1045), .B2(new_n787), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n791), .A2(G1), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT107), .Z(new_n1048));
  OAI21_X1  g0848(.A(new_n1034), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n825), .A2(new_n226), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n818), .B2(G294), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n824), .B2(new_n839), .C1(new_n548), .C2(new_n835), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n832), .A2(new_n496), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT46), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT108), .Z(new_n1055));
  INV_X1    g0855(.A(G317), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n316), .B1(new_n821), .B2(new_n1056), .C1(new_n1053), .C2(KEYINPUT46), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n840), .A2(new_n838), .B1(new_n829), .B2(new_n317), .ZN(new_n1058));
  NOR4_X1   g0858(.A1(new_n1052), .A2(new_n1055), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n847), .A2(G68), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n825), .A2(new_n220), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n817), .A2(new_n849), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(G150), .C2(new_n834), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n429), .B1(new_n832), .B2(new_n202), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n893), .B2(G143), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n891), .A2(G50), .B1(G137), .B2(new_n822), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1059), .B1(new_n1060), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n910), .B1(new_n1068), .B2(KEYINPUT47), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(KEYINPUT47), .B2(new_n1068), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n813), .B1(new_n752), .B2(new_n674), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n244), .A2(new_n800), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n792), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1070), .B(new_n1073), .C1(new_n862), .C2(new_n1014), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1049), .A2(new_n1074), .ZN(G387));
  NAND2_X1  g0875(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n835), .A2(new_n201), .B1(new_n849), .B2(new_n840), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n429), .B1(new_n832), .B2(new_n220), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1077), .A2(new_n1050), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n847), .A2(new_n674), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n203), .A2(new_n839), .B1(new_n817), .B2(new_n441), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G150), .B2(new_n822), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n429), .B1(new_n905), .B2(G116), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n829), .A2(new_n824), .B1(new_n589), .B2(new_n832), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G317), .A2(new_n834), .B1(new_n893), .B2(G322), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n548), .B2(new_n839), .C1(new_n838), .C2(new_n817), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT48), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1088), .B2(new_n1087), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT49), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1084), .B1(new_n821), .B2(new_n841), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1083), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n808), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n755), .ZN(new_n1096));
  AOI211_X1 g0896(.A(G45), .B(new_n1096), .C1(G68), .C2(G77), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT109), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n335), .A2(G50), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT50), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n800), .C1(new_n261), .C2(new_n240), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n429), .A2(new_n208), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1104), .B1(G107), .B2(new_n208), .C1(new_n755), .C2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n792), .B1(new_n1106), .B2(new_n812), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1095), .B(new_n1107), .C1(new_n744), .C2(new_n862), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1044), .A2(new_n787), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(KEYINPUT110), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1044), .A2(new_n787), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1110), .A2(new_n753), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1109), .A2(KEYINPUT110), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1076), .B(new_n1108), .C1(new_n1112), .C2(new_n1113), .ZN(G393));
  INV_X1    g0914(.A(new_n1041), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1111), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n753), .A3(new_n1045), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1017), .A2(new_n811), .A3(new_n1018), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n253), .A2(new_n801), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n812), .B1(new_n226), .B2(new_n208), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n793), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n835), .A2(new_n838), .B1(new_n1056), .B2(new_n840), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT52), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n316), .B1(new_n825), .B2(new_n317), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n839), .A2(new_n589), .B1(new_n829), .B2(new_n496), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(G303), .C2(new_n818), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n821), .A2(new_n836), .B1(new_n824), .B2(new_n832), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT111), .Z(new_n1128));
  NAND3_X1  g0928(.A1(new_n1123), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(G150), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n835), .A2(new_n849), .B1(new_n1130), .B2(new_n840), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT51), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n847), .A2(G77), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n429), .B1(new_n832), .B2(new_n203), .C1(new_n825), .C2(new_n224), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n822), .A2(G143), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n335), .B2(new_n839), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(G50), .C2(new_n818), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1132), .A2(new_n1133), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1129), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1139), .A2(KEYINPUT112), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(new_n910), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(KEYINPUT112), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1121), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1041), .A2(new_n1048), .B1(new_n1118), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1117), .A2(new_n1144), .ZN(G390));
  NAND3_X1  g0945(.A1(new_n996), .A2(G330), .A3(new_n880), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n930), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n994), .A2(new_n784), .A3(G330), .A4(new_n880), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n957), .A2(new_n748), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n961), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n734), .B1(new_n1150), .B2(new_n963), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n879), .A2(new_n689), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n876), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1147), .A2(new_n1148), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n968), .A2(new_n969), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n930), .B1(new_n785), .B2(new_n881), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n994), .A2(new_n996), .A3(G330), .A4(new_n880), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1154), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n486), .A2(G330), .A3(new_n996), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n703), .B(new_n1160), .C1(new_n988), .C2(new_n990), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n971), .A2(new_n982), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n930), .B1(new_n968), .B2(new_n969), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n983), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1153), .A2(new_n930), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n983), .B(KEYINPUT113), .Z(new_n1168));
  NAND3_X1  g0968(.A1(new_n1167), .A2(new_n980), .A3(new_n1168), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1166), .A2(new_n1148), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1157), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1163), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1166), .A2(new_n1148), .A3(new_n1169), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1169), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT100), .B1(new_n874), .B2(new_n875), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n969), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n994), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n983), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1174), .B1(new_n1179), .B2(new_n1164), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1173), .B(new_n1162), .C1(new_n1180), .C2(new_n1157), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1172), .A2(new_n753), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n910), .A2(new_n441), .A3(new_n810), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT54), .B(G143), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n891), .A2(new_n1185), .B1(G50), .B2(new_n905), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n832), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT53), .B1(new_n1187), .B2(G150), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1187), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1186), .B(new_n429), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n893), .A2(G128), .B1(G125), .B2(new_n822), .ZN(new_n1191));
  INV_X1    g0991(.A(G137), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n817), .C1(new_n899), .C2(new_n835), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1190), .B(new_n1193), .C1(G159), .C2(new_n847), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1133), .B1(new_n496), .B2(new_n835), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT114), .Z(new_n1196));
  OAI22_X1  g0996(.A1(new_n317), .A2(new_n817), .B1(new_n840), .B2(new_n824), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n839), .A2(new_n226), .B1(new_n589), .B2(new_n821), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n316), .B1(new_n832), .B2(new_n224), .C1(new_n825), .C2(new_n203), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1194), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n793), .B(new_n1183), .C1(new_n1201), .C2(new_n910), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1164), .B2(new_n809), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n1204), .B2(new_n1048), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1182), .A2(new_n1205), .A3(KEYINPUT115), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT115), .B1(new_n1182), .B2(new_n1205), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(G378));
  INV_X1    g1008(.A(KEYINPUT118), .ZN(new_n1209));
  OAI21_X1  g1009(.A(G330), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1209), .B1(new_n999), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(G330), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1002), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(new_n1213), .B2(new_n980), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n997), .B1(new_n956), .B2(new_n953), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(KEYINPUT118), .C1(KEYINPUT40), .C2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n376), .A2(new_n315), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n312), .A2(new_n947), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1217), .B(new_n1218), .Z(new_n1219));
  XNOR2_X1  g1019(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1219), .B(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1211), .A2(new_n1216), .A3(new_n1222), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1000), .A2(KEYINPUT118), .A3(new_n1214), .A4(new_n1221), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1223), .A2(new_n987), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n987), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1221), .A2(new_n809), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n793), .B1(new_n911), .B2(G50), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n429), .A2(G41), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n220), .B2(new_n832), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n825), .A2(new_n202), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n891), .B2(new_n674), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n824), .B2(new_n821), .C1(new_n317), .C2(new_n835), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1231), .B(new_n1234), .C1(G97), .C2(new_n818), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1060), .B1(new_n496), .B2(new_n840), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1236), .A2(KEYINPUT116), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(KEYINPUT116), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1235), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT58), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n834), .A2(G128), .B1(new_n1187), .B2(new_n1185), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT117), .ZN(new_n1242));
  INV_X1    g1042(.A(G125), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n1243), .A2(new_n840), .B1(new_n839), .B2(new_n1192), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G132), .B2(new_n818), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1242), .B(new_n1245), .C1(new_n1130), .C2(new_n846), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n492), .B(new_n260), .C1(new_n825), .C2(new_n849), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G124), .B2(new_n822), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1240), .B1(new_n1247), .B2(new_n1251), .C1(new_n1230), .C2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1229), .B1(new_n1253), .B2(new_n808), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1227), .A2(new_n1048), .B1(new_n1228), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1161), .B1(new_n1204), .B2(new_n1162), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n987), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1223), .A2(new_n987), .A3(new_n1224), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(KEYINPUT57), .A3(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n753), .B1(new_n1256), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1161), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1181), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1255), .B1(new_n1262), .B2(new_n1265), .ZN(G375));
  INV_X1    g1066(.A(new_n1035), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1158), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1154), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1161), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1163), .A2(new_n1267), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n930), .A2(new_n809), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n793), .B1(new_n911), .B2(G68), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n835), .A2(new_n824), .B1(new_n317), .B2(new_n839), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(G294), .B2(new_n893), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n429), .B(new_n1061), .C1(G97), .C2(new_n1187), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n818), .A2(G116), .B1(G303), .B2(new_n822), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1276), .A2(new_n1080), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n835), .A2(new_n1192), .B1(new_n1130), .B2(new_n839), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(G132), .B2(new_n893), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n316), .B(new_n1232), .C1(G159), .C2(new_n1187), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n818), .A2(new_n1185), .B1(G128), .B2(new_n822), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n846), .A2(new_n201), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1279), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1274), .B1(new_n1286), .B2(new_n808), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1272), .A2(new_n1048), .B1(new_n1273), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1271), .A2(new_n1288), .ZN(G381));
  INV_X1    g1089(.A(G390), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1049), .A2(new_n1074), .A3(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1182), .A2(new_n1205), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1228), .A2(new_n1254), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1048), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT57), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1225), .A2(new_n1226), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n754), .B1(new_n1300), .B2(new_n1264), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1299), .B1(new_n1256), .B2(new_n1296), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1298), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  OR2_X1    g1103(.A1(G393), .A2(G396), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1304), .A2(G384), .A3(G381), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1292), .A2(new_n1294), .A3(new_n1303), .A4(new_n1305), .ZN(G407));
  NAND2_X1  g1106(.A1(new_n733), .A2(G213), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1303), .A2(new_n1294), .A3(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(G407), .A2(G213), .A3(new_n1309), .ZN(G409));
  INV_X1    g1110(.A(KEYINPUT125), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT115), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1293), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1182), .A2(new_n1205), .A3(KEYINPUT115), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1312), .A2(new_n1314), .A3(new_n1315), .A4(new_n1255), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1227), .A2(new_n1264), .A3(new_n1267), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1255), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1294), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1308), .B1(new_n1316), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1308), .A2(G2897), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n754), .B1(new_n1263), .B2(new_n1272), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT60), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1270), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1159), .A2(KEYINPUT60), .A3(new_n1161), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1323), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1327), .A2(G384), .A3(new_n1288), .ZN(new_n1328));
  AOI21_X1  g1128(.A(G384), .B1(new_n1327), .B2(new_n1288), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1322), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT121), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  OAI211_X1 g1132(.A(KEYINPUT121), .B(new_n1322), .C1(new_n1328), .C2(new_n1329), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(G384), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1159), .A2(KEYINPUT60), .A3(new_n1161), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n753), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT60), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1336), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1288), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1335), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1327), .A2(G384), .A3(new_n1288), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1341), .A2(new_n1342), .A3(new_n1321), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT120), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1341), .A2(KEYINPUT120), .A3(new_n1342), .A4(new_n1321), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT122), .ZN(new_n1348));
  AND3_X1   g1148(.A1(new_n1334), .A2(new_n1347), .A3(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1348), .B1(new_n1334), .B2(new_n1347), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1320), .A2(new_n1349), .A3(new_n1350), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1311), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1352), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1350), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1334), .A2(new_n1347), .A3(new_n1348), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  OAI211_X1 g1157(.A(KEYINPUT125), .B(new_n1354), .C1(new_n1357), .C2(new_n1320), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1353), .A2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(G387), .A2(G390), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1304), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(G393), .A2(G396), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1362), .ZN(new_n1363));
  OAI21_X1  g1163(.A(KEYINPUT123), .B1(new_n1361), .B2(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1360), .A2(new_n1291), .A3(new_n1364), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(new_n1361), .A2(new_n1363), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT123), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1366), .A2(new_n1367), .ZN(new_n1368));
  XNOR2_X1  g1168(.A(new_n1365), .B(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n1319), .B1(new_n1370), .B2(G375), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1371), .A2(new_n1307), .A3(new_n1372), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1373), .A2(KEYINPUT62), .ZN(new_n1374));
  INV_X1    g1174(.A(KEYINPUT62), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1375), .B1(new_n1320), .B2(new_n1372), .ZN(new_n1376));
  NOR3_X1   g1176(.A1(new_n1369), .A2(new_n1374), .A3(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1373), .A2(KEYINPUT63), .ZN(new_n1378));
  INV_X1    g1178(.A(KEYINPUT63), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n1320), .A2(new_n1379), .A3(new_n1372), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1378), .A2(new_n1380), .ZN(new_n1381));
  AOI21_X1  g1181(.A(new_n1293), .B1(new_n1255), .B2(new_n1317), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1382), .B1(G378), .B2(new_n1303), .ZN(new_n1383));
  OAI21_X1  g1183(.A(KEYINPUT119), .B1(new_n1383), .B2(new_n1308), .ZN(new_n1384));
  INV_X1    g1184(.A(KEYINPUT119), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1371), .A2(new_n1385), .A3(new_n1307), .ZN(new_n1386));
  NAND4_X1  g1186(.A1(new_n1384), .A2(new_n1386), .A3(new_n1356), .A4(new_n1355), .ZN(new_n1387));
  INV_X1    g1187(.A(KEYINPUT61), .ZN(new_n1388));
  NAND3_X1  g1188(.A1(new_n1381), .A2(new_n1387), .A3(new_n1388), .ZN(new_n1389));
  AOI22_X1  g1189(.A1(new_n1359), .A2(new_n1377), .B1(new_n1369), .B2(new_n1389), .ZN(G405));
  NOR2_X1   g1190(.A1(new_n1372), .A2(KEYINPUT126), .ZN(new_n1391));
  NOR2_X1   g1191(.A1(new_n1370), .A2(G375), .ZN(new_n1392));
  AND2_X1   g1192(.A1(new_n1372), .A2(KEYINPUT126), .ZN(new_n1393));
  OR2_X1    g1193(.A1(new_n1392), .A2(new_n1393), .ZN(new_n1394));
  NOR2_X1   g1194(.A1(new_n1303), .A2(new_n1293), .ZN(new_n1395));
  OAI21_X1  g1195(.A(new_n1391), .B1(new_n1394), .B2(new_n1395), .ZN(new_n1396));
  OR4_X1    g1196(.A1(new_n1392), .A2(new_n1395), .A3(new_n1391), .A4(new_n1393), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1396), .A2(new_n1397), .ZN(new_n1398));
  XNOR2_X1  g1198(.A(new_n1398), .B(new_n1369), .ZN(G402));
endmodule


