//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  OAI21_X1  g000(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT0), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n194), .A2(new_n196), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G143), .B(G146), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n192), .A2(new_n199), .B1(new_n191), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT4), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT74), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT3), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT74), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n205), .A2(new_n207), .B1(G104), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G107), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(KEYINPUT74), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n203), .B(G101), .C1(new_n209), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT76), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n205), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n213), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n208), .A2(G104), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n210), .A2(G107), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(new_n205), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT76), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n222), .A2(new_n223), .A3(new_n203), .A4(G101), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n202), .B1(new_n216), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT75), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n209), .A2(new_n214), .ZN(new_n227));
  INV_X1    g041(.A(G101), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n203), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(G101), .B1(new_n209), .B2(new_n214), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n218), .A2(new_n221), .A3(new_n228), .ZN(new_n232));
  AND4_X1   g046(.A1(new_n226), .A2(new_n230), .A3(new_n232), .A4(KEYINPUT4), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n225), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n235));
  INV_X1    g049(.A(G134), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G137), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT11), .A3(G134), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(G137), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G131), .ZN(new_n242));
  INV_X1    g056(.A(G131), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n237), .A2(new_n239), .A3(new_n243), .A4(new_n240), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n194), .B(new_n196), .C1(KEYINPUT1), .C2(new_n190), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n194), .A2(new_n196), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT1), .B1(new_n195), .B2(G146), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(G128), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n228), .B1(new_n213), .B2(new_n211), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n232), .A2(new_n247), .A3(new_n250), .A4(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT10), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n250), .A2(new_n247), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT10), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n256), .A2(new_n257), .A3(new_n232), .A4(new_n252), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n234), .A2(new_n246), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT77), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(KEYINPUT12), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n209), .A2(new_n214), .A3(G101), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n263), .A2(new_n255), .A3(new_n251), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n232), .A2(new_n252), .B1(new_n247), .B2(new_n250), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n245), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT12), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(KEYINPUT77), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n262), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n255), .B1(new_n263), .B2(new_n251), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n246), .B1(new_n271), .B2(new_n253), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n272), .A2(new_n261), .A3(KEYINPUT12), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n260), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  INV_X1    g089(.A(G227), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G953), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n275), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G469), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n234), .A2(new_n259), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n245), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n278), .A3(new_n260), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n280), .A2(new_n281), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n281), .A2(new_n285), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n262), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(new_n272), .B2(new_n268), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n266), .A2(KEYINPUT77), .A3(new_n267), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n279), .B1(new_n292), .B2(new_n260), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n283), .A2(new_n279), .A3(new_n260), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n286), .B(new_n288), .C1(new_n296), .C2(new_n281), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  OAI21_X1  g112(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G140), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G125), .ZN(new_n302));
  INV_X1    g116(.A(G125), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G140), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n304), .A3(KEYINPUT16), .ZN(new_n305));
  OR3_X1    g119(.A1(new_n303), .A2(KEYINPUT16), .A3(G140), .ZN(new_n306));
  AOI21_X1  g120(.A(G146), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n305), .A2(G146), .A3(new_n306), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n305), .A2(new_n306), .A3(G146), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT69), .ZN(new_n312));
  INV_X1    g126(.A(G237), .ZN(new_n313));
  INV_X1    g127(.A(G953), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(G214), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(new_n195), .ZN(new_n316));
  NOR2_X1   g130(.A1(G237), .A2(G953), .ZN(new_n317));
  AOI21_X1  g131(.A(G143), .B1(new_n317), .B2(G214), .ZN(new_n318));
  OAI21_X1  g132(.A(G131), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT17), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n195), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n317), .A2(G143), .A3(G214), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n243), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(KEYINPUT17), .B(G131), .C1(new_n316), .C2(new_n318), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n310), .A2(new_n312), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(G113), .B(G122), .Z(new_n327));
  XOR2_X1   g141(.A(KEYINPUT82), .B(G104), .Z(new_n328));
  XOR2_X1   g142(.A(new_n327), .B(new_n328), .Z(new_n329));
  OAI211_X1 g143(.A(KEYINPUT18), .B(G131), .C1(new_n316), .C2(new_n318), .ZN(new_n330));
  NAND2_X1  g144(.A1(KEYINPUT18), .A2(G131), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n321), .A2(new_n322), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n302), .A2(new_n304), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G146), .ZN(new_n334));
  XNOR2_X1  g148(.A(G125), .B(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n193), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n330), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n326), .A2(new_n329), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n329), .B1(new_n326), .B2(new_n338), .ZN(new_n341));
  OAI211_X1 g155(.A(KEYINPUT83), .B(new_n285), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G475), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n324), .A2(new_n325), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n305), .A2(new_n306), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n193), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n305), .A2(new_n306), .A3(new_n309), .A4(G146), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n312), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n338), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n329), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(G902), .B1(new_n351), .B2(new_n339), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(KEYINPUT83), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n319), .A2(new_n323), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT19), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n335), .B(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n354), .B(new_n311), .C1(G146), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n338), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n350), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n339), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT20), .ZN(new_n361));
  NOR2_X1   g175(.A1(G475), .A2(G902), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n361), .B1(new_n360), .B2(new_n362), .ZN(new_n365));
  OAI22_X1  g179(.A1(new_n343), .A2(new_n353), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(G234), .A2(G237), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(G952), .A3(new_n314), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(KEYINPUT87), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n367), .A2(G902), .A3(G953), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT21), .B(G898), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G116), .B(G122), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT14), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n378));
  INV_X1    g192(.A(G122), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G116), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n208), .B1(new_n380), .B2(KEYINPUT14), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n378), .B1(new_n377), .B2(new_n381), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n375), .A2(new_n208), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT84), .B1(new_n190), .B2(G143), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT84), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n195), .A3(G128), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n195), .A2(G128), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n236), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n236), .B1(new_n389), .B2(new_n391), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n385), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT13), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n390), .B1(new_n389), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n386), .A2(new_n388), .A3(KEYINPUT13), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n236), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n375), .B(new_n208), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n392), .ZN(new_n401));
  OAI22_X1  g215(.A1(new_n384), .A2(new_n395), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G217), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n298), .A2(new_n403), .A3(G953), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n404), .ZN(new_n406));
  OAI221_X1 g220(.A(new_n406), .B1(new_n401), .B2(new_n399), .C1(new_n395), .C2(new_n384), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n407), .A3(new_n285), .ZN(new_n408));
  INV_X1    g222(.A(G478), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(KEYINPUT15), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n410), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n405), .A2(new_n407), .A3(new_n285), .A4(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(KEYINPUT86), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT86), .B1(new_n411), .B2(new_n413), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n374), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n300), .A2(new_n366), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT73), .ZN(new_n419));
  INV_X1    g233(.A(G234), .ZN(new_n420));
  OAI21_X1  g234(.A(G217), .B1(new_n420), .B2(G902), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT67), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT25), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n314), .A2(G221), .A3(G234), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT71), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT22), .B(G137), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT68), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n190), .A2(G119), .ZN(new_n430));
  INV_X1    g244(.A(G119), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G128), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT24), .B(G110), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G110), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT24), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT24), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G110), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G119), .B(G128), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT68), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n431), .A2(G128), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n443), .B(new_n432), .C1(new_n444), .C2(KEYINPUT23), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n435), .A2(new_n442), .B1(G110), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n348), .A2(new_n446), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n311), .A2(new_n336), .ZN(new_n448));
  OAI22_X1  g262(.A1(new_n445), .A2(G110), .B1(new_n441), .B2(new_n440), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n428), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT70), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n445), .A2(G110), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n433), .A2(new_n434), .A3(new_n429), .ZN(new_n454));
  AOI21_X1  g268(.A(KEYINPUT68), .B1(new_n440), .B2(new_n441), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(new_n310), .B2(new_n312), .ZN(new_n457));
  INV_X1    g271(.A(new_n450), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n452), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n447), .A2(KEYINPUT70), .A3(new_n450), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n451), .B1(new_n461), .B2(new_n428), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n423), .B1(new_n462), .B2(G902), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n447), .A2(KEYINPUT70), .A3(new_n450), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT70), .B1(new_n447), .B2(new_n450), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n428), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n451), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(KEYINPUT25), .A3(new_n285), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n422), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(G902), .B1(new_n420), .B2(G217), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT72), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n462), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n419), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n422), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT25), .B1(new_n468), .B2(new_n285), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n423), .B(G902), .C1(new_n466), .C2(new_n467), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n474), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(KEYINPUT73), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G472), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n431), .A2(G116), .ZN(new_n484));
  INV_X1    g298(.A(G116), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G119), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT2), .B(G113), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n488), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n245), .A2(new_n201), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n494));
  INV_X1    g308(.A(new_n240), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n236), .A2(G137), .ZN(new_n496));
  OAI21_X1  g310(.A(G131), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n250), .A2(new_n497), .A3(new_n244), .A4(new_n247), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n494), .B1(new_n493), .B2(new_n498), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n492), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT31), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n317), .A2(G210), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT27), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT26), .B(G101), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n497), .A2(new_n244), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n256), .A2(new_n507), .B1(new_n245), .B2(new_n201), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n491), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n501), .A2(new_n502), .A3(new_n506), .A4(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT28), .B1(new_n508), .B2(new_n491), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n493), .A2(new_n498), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n492), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n511), .B1(new_n514), .B2(KEYINPUT28), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n506), .B(KEYINPUT65), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n512), .A2(new_n492), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n512), .A2(KEYINPUT30), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n518), .B1(new_n521), .B2(new_n492), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n502), .B1(new_n522), .B2(new_n506), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n483), .B(new_n285), .C1(new_n517), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT32), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n501), .A2(new_n506), .A3(new_n509), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT31), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(new_n510), .C1(new_n515), .C2(new_n516), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT32), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n483), .A4(new_n285), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n515), .A2(KEYINPUT29), .A3(new_n506), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT66), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n522), .B2(new_n506), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n501), .A2(new_n509), .ZN(new_n534));
  INV_X1    g348(.A(new_n506), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(KEYINPUT66), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n515), .A2(new_n516), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n285), .B(new_n531), .C1(new_n537), .C2(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n525), .A2(new_n530), .B1(new_n541), .B2(G472), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n482), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G214), .B1(G237), .B2(G902), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT78), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n255), .A2(new_n303), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n303), .B2(new_n201), .ZN(new_n547));
  INV_X1    g361(.A(G224), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(G953), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n547), .B(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n491), .B1(new_n216), .B2(new_n224), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n231), .B2(new_n233), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n484), .A2(new_n486), .A3(KEYINPUT5), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n553), .B(G113), .C1(KEYINPUT5), .C2(new_n484), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n232), .A2(new_n489), .A3(new_n554), .A4(new_n252), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT6), .ZN(new_n557));
  XNOR2_X1  g371(.A(G110), .B(G122), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT79), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n556), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n552), .A2(new_n555), .A3(new_n558), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT6), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n552), .B2(new_n555), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n550), .B(new_n562), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT7), .B1(new_n548), .B2(G953), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n547), .B(new_n567), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n555), .A2(KEYINPUT80), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n554), .A2(new_n489), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n263), .B2(new_n251), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n555), .A2(KEYINPUT80), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n558), .B(KEYINPUT8), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n568), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(G902), .B1(new_n575), .B2(new_n563), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n566), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G210), .B1(G237), .B2(G902), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT81), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n579), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n566), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n545), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n418), .A2(new_n543), .A3(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT88), .B(G101), .Z(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(G3));
  OAI21_X1  g400(.A(new_n285), .B1(new_n517), .B2(new_n523), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G472), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n524), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n482), .A2(new_n300), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n580), .A2(KEYINPUT89), .A3(new_n582), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n405), .A2(new_n407), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT90), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT90), .A4(new_n592), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n404), .A2(KEYINPUT91), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n592), .B1(new_n402), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n402), .B2(new_n597), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n409), .A2(G902), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n595), .A2(new_n596), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n408), .A2(new_n409), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n366), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n544), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n581), .B1(new_n566), .B2(new_n576), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT89), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND4_X1   g423(.A1(new_n374), .A2(new_n591), .A3(new_n605), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n590), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  NOR3_X1   g427(.A1(new_n366), .A2(new_n415), .A3(new_n416), .ZN(new_n614));
  AND4_X1   g428(.A1(new_n374), .A2(new_n591), .A3(new_n609), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n590), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  INV_X1    g432(.A(new_n589), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT36), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n427), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(KEYINPUT92), .Z(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n461), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n459), .A3(new_n460), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n473), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n479), .A3(KEYINPUT93), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT93), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n470), .B2(new_n626), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n418), .A2(new_n583), .A3(new_n619), .A4(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT37), .B(G110), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G12));
  NAND2_X1  g448(.A1(new_n525), .A2(new_n530), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n541), .A2(G472), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n630), .A2(new_n628), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n591), .A2(new_n609), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT94), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n640), .A2(KEYINPUT94), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n370), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n369), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT95), .ZN(new_n645));
  NOR4_X1   g459(.A1(new_n366), .A2(new_n415), .A3(new_n416), .A4(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n646), .A2(new_n299), .A3(new_n297), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n639), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  INV_X1    g463(.A(new_n582), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n607), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n526), .ZN(new_n654));
  INV_X1    g468(.A(new_n516), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n514), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n656), .B2(G902), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n635), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n352), .A2(KEYINPUT83), .ZN(new_n660));
  INV_X1    g474(.A(G475), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n352), .B2(KEYINPUT83), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n360), .A2(new_n362), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT20), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n660), .A2(new_n662), .B1(new_n664), .B2(new_n363), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n665), .A2(new_n415), .A3(new_n416), .ZN(new_n666));
  AND4_X1   g480(.A1(new_n544), .A2(new_n630), .A3(new_n628), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT97), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n659), .A2(KEYINPUT97), .A3(new_n667), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT98), .B(KEYINPUT39), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n645), .B(new_n672), .Z(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n297), .A2(new_n299), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT40), .Z(new_n676));
  NAND3_X1  g490(.A1(new_n670), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G143), .ZN(G45));
  INV_X1    g492(.A(new_n645), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n366), .A2(new_n603), .A3(new_n679), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n680), .A2(new_n297), .A3(new_n299), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n639), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  NAND2_X1  g497(.A1(new_n286), .A2(new_n299), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n280), .A2(new_n285), .A3(new_n284), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n686), .A2(new_n687), .A3(G469), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n687), .B1(new_n686), .B2(G469), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n685), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT100), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n234), .A2(new_n246), .A3(new_n259), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n246), .B1(new_n234), .B2(new_n259), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n692), .A2(new_n693), .A3(new_n279), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n278), .B1(new_n292), .B2(new_n260), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n694), .A2(new_n695), .A3(G902), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT99), .B1(new_n696), .B2(new_n281), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n686), .A2(new_n687), .A3(G469), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n684), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n610), .A2(new_n543), .A3(new_n691), .A4(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n697), .A2(new_n698), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n700), .B1(new_n705), .B2(new_n685), .ZN(new_n706));
  AOI211_X1 g520(.A(KEYINPUT100), .B(new_n684), .C1(new_n697), .C2(new_n698), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(KEYINPUT101), .A3(new_n543), .A4(new_n610), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND4_X1  g526(.A1(new_n615), .A2(new_n543), .A3(new_n691), .A4(new_n701), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n708), .A2(KEYINPUT102), .A3(new_n543), .A4(new_n615), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  NOR2_X1   g532(.A1(new_n417), .A2(new_n366), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n705), .A2(new_n719), .A3(new_n685), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n638), .A3(new_n637), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  NAND3_X1  g537(.A1(new_n701), .A2(new_n691), .A3(new_n374), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n591), .A2(new_n609), .A3(new_n666), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n479), .A2(new_n480), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n588), .A2(new_n727), .A3(new_n524), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n587), .A2(KEYINPUT103), .A3(G472), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n724), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT104), .B(G122), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G24));
  AOI22_X1  g548(.A1(new_n630), .A2(new_n628), .B1(new_n728), .B2(new_n729), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n638), .A3(new_n680), .A4(new_n699), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT105), .B(G125), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G27));
  INV_X1    g552(.A(new_n299), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n286), .A2(new_n288), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n692), .A2(new_n693), .A3(new_n278), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT106), .B1(new_n741), .B2(new_n293), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n295), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(G469), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n739), .B1(new_n740), .B2(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n650), .A2(new_n607), .A3(new_n606), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(new_n543), .ZN(new_n749));
  INV_X1    g563(.A(new_n680), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(KEYINPUT42), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n542), .A2(new_n726), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n746), .A3(new_n680), .A4(new_n747), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n749), .A2(new_n751), .B1(KEYINPUT42), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  NAND3_X1  g569(.A1(new_n748), .A2(new_n543), .A3(new_n646), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  NAND2_X1  g571(.A1(new_n665), .A2(new_n603), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n589), .A3(new_n631), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n747), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n742), .A2(KEYINPUT45), .A3(new_n744), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n296), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(G469), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n288), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n288), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n286), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n299), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT108), .B1(new_n777), .B2(new_n673), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n776), .A2(new_n779), .A3(new_n299), .A4(new_n674), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n765), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n238), .ZN(G39));
  AND4_X1   g596(.A1(new_n542), .A2(new_n482), .A3(new_n680), .A4(new_n747), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT47), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n777), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n776), .A2(KEYINPUT47), .A3(new_n299), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n301), .ZN(G42));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n790));
  INV_X1    g604(.A(new_n369), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n760), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n730), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n793), .A2(new_n544), .A3(new_n653), .A4(new_n690), .ZN(new_n794));
  OR2_X1    g608(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n747), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n797), .A2(new_n690), .A3(new_n658), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(new_n475), .A3(new_n481), .A4(new_n791), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n366), .A3(new_n603), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT116), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n792), .A2(new_n699), .A3(new_n735), .A4(new_n747), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n796), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT117), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n786), .A2(new_n787), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n705), .A2(new_n286), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n299), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n793), .A2(new_n797), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT114), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n803), .A2(KEYINPUT117), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n804), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n808), .A2(KEYINPUT114), .A3(new_n810), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n790), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n792), .A2(new_n699), .A3(new_n752), .A4(new_n747), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT48), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n638), .A2(new_n792), .A3(new_n699), .A4(new_n730), .ZN(new_n818));
  INV_X1    g632(.A(G952), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n818), .A2(new_n819), .A3(G953), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n817), .B(new_n820), .C1(new_n604), .C2(new_n799), .ZN(new_n821));
  AND4_X1   g635(.A1(KEYINPUT51), .A2(new_n796), .A3(new_n801), .A4(new_n802), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n808), .B2(new_n810), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n822), .B(KEYINPUT118), .C1(new_n808), .C2(new_n810), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n821), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n815), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n637), .B(new_n638), .C1(new_n647), .C2(new_n681), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n470), .A2(new_n626), .A3(new_n645), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n725), .A2(new_n746), .A3(new_n658), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n829), .A2(new_n736), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n829), .A2(new_n736), .A3(new_n831), .A4(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT111), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n583), .A2(new_n837), .A3(new_n374), .A4(new_n605), .ZN(new_n838));
  INV_X1    g652(.A(new_n545), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n839), .B(new_n374), .C1(new_n650), .C2(new_n607), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT111), .B1(new_n840), .B2(new_n604), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n590), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n411), .A2(new_n413), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n665), .A2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n583), .A2(new_n374), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n590), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n842), .A2(new_n632), .A3(new_n846), .A4(new_n584), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n748), .A2(new_n680), .A3(new_n735), .ZN(new_n848));
  INV_X1    g662(.A(new_n300), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n366), .A2(new_n843), .A3(new_n645), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n637), .A2(new_n849), .A3(new_n747), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n756), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n836), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n706), .A2(new_n707), .A3(new_n373), .ZN(new_n855));
  INV_X1    g669(.A(new_n731), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n855), .A2(new_n856), .B1(new_n639), .B2(new_n721), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n710), .A2(new_n717), .A3(new_n754), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n854), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n854), .B2(new_n858), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n860), .B1(KEYINPUT112), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(KEYINPUT112), .B2(new_n861), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n836), .A2(KEYINPUT53), .A3(new_n853), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n858), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n722), .B1(new_n724), .B2(new_n731), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n704), .B2(new_n709), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(KEYINPUT113), .A3(new_n717), .A4(new_n754), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n865), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n872), .A3(new_n861), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  OAI22_X1  g688(.A1(new_n828), .A2(new_n874), .B1(G952), .B2(G953), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n665), .A2(new_n603), .A3(new_n839), .A4(new_n299), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n726), .B(new_n876), .C1(new_n806), .C2(KEYINPUT49), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT109), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n653), .A2(new_n658), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n878), .B(new_n879), .C1(KEYINPUT49), .C2(new_n806), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT110), .Z(new_n881));
  NAND2_X1  g695(.A1(new_n875), .A2(new_n881), .ZN(G75));
  INV_X1    g696(.A(KEYINPUT56), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n871), .A2(new_n861), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(G902), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n885), .B2(new_n581), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(new_n550), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT55), .Z(new_n889));
  AND2_X1   g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n886), .A2(new_n889), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n314), .A2(G952), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G51));
  NOR2_X1   g707(.A1(new_n885), .A2(new_n771), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n694), .A2(new_n695), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  XNOR2_X1  g710(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n287), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n871), .A2(new_n872), .A3(new_n861), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n872), .B1(new_n871), .B2(new_n861), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n896), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI211_X1 g717(.A(KEYINPUT120), .B(new_n898), .C1(new_n899), .C2(new_n900), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n894), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT121), .B1(new_n905), .B2(new_n892), .ZN(new_n906));
  INV_X1    g720(.A(new_n894), .ZN(new_n907));
  INV_X1    g721(.A(new_n898), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(new_n873), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n895), .B1(new_n910), .B2(KEYINPUT120), .ZN(new_n911));
  INV_X1    g725(.A(new_n904), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n907), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n914));
  INV_X1    g728(.A(new_n892), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n906), .A2(new_n916), .ZN(G54));
  NAND2_X1  g731(.A1(KEYINPUT58), .A2(G475), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT122), .Z(new_n919));
  NOR2_X1   g733(.A1(new_n885), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n915), .B1(new_n920), .B2(new_n360), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n360), .B2(new_n920), .ZN(G60));
  NAND3_X1  g736(.A1(new_n595), .A2(new_n596), .A3(new_n599), .ZN(new_n923));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT59), .Z(new_n925));
  AOI211_X1 g739(.A(new_n923), .B(new_n925), .C1(new_n909), .C2(new_n873), .ZN(new_n926));
  INV_X1    g740(.A(new_n925), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n874), .A2(new_n927), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n892), .B(new_n926), .C1(new_n928), .C2(new_n923), .ZN(G63));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT60), .Z(new_n931));
  AND2_X1   g745(.A1(new_n884), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n915), .B1(new_n932), .B2(new_n468), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n624), .A2(new_n625), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n934), .B2(new_n932), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g750(.A(new_n371), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n314), .B1(new_n937), .B2(G224), .ZN(new_n938));
  INV_X1    g752(.A(new_n847), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n869), .A2(new_n717), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n940), .B2(new_n314), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n887), .B1(G898), .B2(new_n314), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n941), .B(new_n942), .Z(G69));
  XOR2_X1   g757(.A(new_n521), .B(new_n356), .Z(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n640), .B2(new_n314), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n778), .A2(new_n780), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n725), .A3(new_n752), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n754), .A2(new_n756), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n788), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n765), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n829), .A2(new_n736), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n954), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT124), .B1(new_n781), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n950), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n945), .B1(new_n958), .B2(new_n314), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n314), .B1(G227), .B2(G900), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n677), .A2(new_n954), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT123), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n605), .A2(new_n844), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n797), .A2(new_n965), .A3(new_n675), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n543), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n961), .B2(KEYINPUT62), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n781), .A2(new_n968), .A3(new_n788), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n944), .B1(new_n970), .B2(new_n314), .ZN(new_n971));
  OR3_X1    g785(.A1(new_n959), .A2(new_n960), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n960), .B1(new_n959), .B2(new_n971), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(G72));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT125), .Z(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n970), .B2(new_n940), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(new_n506), .A3(new_n534), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n863), .B(new_n976), .C1(new_n654), .C2(new_n537), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n522), .A2(new_n535), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT126), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n955), .A2(new_n957), .ZN(new_n985));
  INV_X1    g799(.A(new_n950), .ZN(new_n986));
  INV_X1    g800(.A(new_n940), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n984), .B1(new_n988), .B2(new_n978), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT127), .B1(new_n989), .B2(new_n892), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n977), .B1(new_n958), .B2(new_n987), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n991), .B(new_n915), .C1(new_n992), .C2(new_n984), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n982), .B1(new_n990), .B2(new_n993), .ZN(G57));
endmodule


