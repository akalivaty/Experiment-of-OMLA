

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752;

  AND2_X1 U371 ( .A1(n723), .A2(G210), .ZN(n633) );
  AND2_X1 U372 ( .A1(n375), .A2(n377), .ZN(n349) );
  XNOR2_X1 U373 ( .A(n450), .B(KEYINPUT3), .ZN(n451) );
  BUF_X1 U374 ( .A(G143), .Z(n350) );
  NAND2_X1 U375 ( .A1(n349), .A2(n373), .ZN(n550) );
  INV_X1 U376 ( .A(KEYINPUT18), .ZN(n391) );
  NOR2_X1 U377 ( .A1(G953), .A2(G237), .ZN(n481) );
  XNOR2_X1 U378 ( .A(n526), .B(n385), .ZN(n406) );
  XNOR2_X1 U379 ( .A(n593), .B(n532), .ZN(n596) );
  AND2_X1 U380 ( .A1(n516), .A2(n515), .ZN(n665) );
  NAND2_X2 U381 ( .A1(n550), .A2(n669), .ZN(n384) );
  XNOR2_X2 U382 ( .A(n384), .B(KEYINPUT40), .ZN(n636) );
  OR2_X2 U383 ( .A1(n638), .A2(G902), .ZN(n393) );
  XNOR2_X2 U384 ( .A(n490), .B(n489), .ZN(n523) );
  NOR2_X1 U385 ( .A1(n715), .A2(n591), .ZN(n576) );
  NOR2_X1 U386 ( .A1(n530), .A2(n566), .ZN(n458) );
  INV_X1 U387 ( .A(n703), .ZN(n403) );
  NOR2_X1 U388 ( .A1(n502), .A2(n517), .ZN(n503) );
  AND2_X1 U389 ( .A1(n514), .A2(n524), .ZN(n669) );
  AND2_X1 U390 ( .A1(n383), .A2(n382), .ZN(n381) );
  XNOR2_X1 U391 ( .A(n407), .B(KEYINPUT108), .ZN(n521) );
  XNOR2_X1 U392 ( .A(n503), .B(KEYINPUT30), .ZN(n392) );
  BUF_X1 U393 ( .A(n502), .Z(n566) );
  XNOR2_X1 U394 ( .A(n531), .B(KEYINPUT104), .ZN(n502) );
  XNOR2_X1 U395 ( .A(n387), .B(n386), .ZN(n725) );
  XNOR2_X1 U396 ( .A(n391), .B(G125), .ZN(n390) );
  XNOR2_X1 U397 ( .A(KEYINPUT84), .B(KEYINPUT17), .ZN(n389) );
  XNOR2_X2 U398 ( .A(n462), .B(n461), .ZN(n737) );
  XNOR2_X1 U399 ( .A(n351), .B(KEYINPUT48), .ZN(n367) );
  NAND2_X1 U400 ( .A1(n542), .A2(n541), .ZN(n351) );
  XNOR2_X2 U401 ( .A(n465), .B(G134), .ZN(n447) );
  XNOR2_X1 U402 ( .A(KEYINPUT79), .B(KEYINPUT46), .ZN(n512) );
  NAND2_X1 U403 ( .A1(n367), .A2(KEYINPUT78), .ZN(n365) );
  NOR2_X1 U404 ( .A1(n549), .A2(n361), .ZN(n368) );
  NOR2_X1 U405 ( .A1(n406), .A2(n504), .ZN(n404) );
  XNOR2_X1 U406 ( .A(n397), .B(n396), .ZN(n741) );
  INV_X1 U407 ( .A(G140), .ZN(n396) );
  XNOR2_X1 U408 ( .A(KEYINPUT10), .B(G125), .ZN(n397) );
  XNOR2_X1 U409 ( .A(n429), .B(n428), .ZN(n388) );
  XNOR2_X1 U410 ( .A(n741), .B(G146), .ZN(n480) );
  XOR2_X1 U411 ( .A(n574), .B(n573), .Z(n715) );
  AND2_X1 U412 ( .A1(n400), .A2(n399), .ZN(n398) );
  XNOR2_X1 U413 ( .A(n659), .B(KEYINPUT102), .ZN(n551) );
  OR2_X2 U414 ( .A1(n526), .A2(n517), .ZN(n535) );
  NAND2_X1 U415 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U416 ( .A(G237), .ZN(n470) );
  XNOR2_X1 U417 ( .A(G128), .B(KEYINPUT90), .ZN(n427) );
  XNOR2_X1 U418 ( .A(G101), .B(G104), .ZN(n494) );
  AND2_X1 U419 ( .A1(n551), .A2(n663), .ZN(n705) );
  NAND2_X1 U420 ( .A1(n366), .A2(n365), .ZN(n364) );
  NAND2_X1 U421 ( .A1(n549), .A2(n361), .ZN(n363) );
  INV_X1 U422 ( .A(KEYINPUT38), .ZN(n385) );
  XOR2_X1 U423 ( .A(KEYINPUT70), .B(KEYINPUT22), .Z(n560) );
  XNOR2_X1 U424 ( .A(n742), .B(n394), .ZN(n638) );
  XOR2_X1 U425 ( .A(G122), .B(G104), .Z(n483) );
  INV_X1 U426 ( .A(G128), .ZN(n419) );
  INV_X1 U427 ( .A(n521), .ZN(n405) );
  XNOR2_X1 U428 ( .A(n395), .B(KEYINPUT101), .ZN(n659) );
  XNOR2_X1 U429 ( .A(n480), .B(n353), .ZN(n386) );
  XNOR2_X1 U430 ( .A(n431), .B(n388), .ZN(n387) );
  XNOR2_X1 U431 ( .A(n370), .B(n358), .ZN(n750) );
  NOR2_X1 U432 ( .A1(n543), .A2(n535), .ZN(n537) );
  NAND2_X1 U433 ( .A1(n578), .A2(n577), .ZN(n369) );
  NAND2_X1 U434 ( .A1(n600), .A2(n563), .ZN(n565) );
  NOR2_X1 U435 ( .A1(n663), .A2(n408), .ZN(n664) );
  AND2_X1 U436 ( .A1(n392), .A2(n355), .ZN(n352) );
  XOR2_X1 U437 ( .A(n424), .B(n423), .Z(n353) );
  NAND2_X1 U438 ( .A1(n701), .A2(n491), .ZN(n354) );
  AND2_X1 U439 ( .A1(n404), .A2(n374), .ZN(n355) );
  NOR2_X1 U440 ( .A1(n406), .A2(n354), .ZN(n356) );
  NOR2_X1 U441 ( .A1(n372), .A2(G900), .ZN(n357) );
  XOR2_X1 U442 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n358) );
  NOR2_X1 U443 ( .A1(n659), .A2(n408), .ZN(n359) );
  INV_X1 U444 ( .A(KEYINPUT41), .ZN(n491) );
  INV_X1 U445 ( .A(KEYINPUT78), .ZN(n361) );
  XOR2_X1 U446 ( .A(n632), .B(n631), .Z(n360) );
  NOR2_X2 U447 ( .A1(n364), .A2(n362), .ZN(n679) );
  NOR2_X1 U448 ( .A1(n363), .A2(n367), .ZN(n362) );
  NOR2_X1 U449 ( .A1(n368), .A2(n627), .ZN(n366) );
  XNOR2_X2 U450 ( .A(n369), .B(n579), .ZN(n751) );
  NOR2_X1 U451 ( .A1(n588), .A2(n596), .ZN(n572) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n410) );
  NAND2_X2 U453 ( .A1(n381), .A2(n378), .ZN(n600) );
  XNOR2_X2 U454 ( .A(n449), .B(n448), .ZN(n452) );
  XNOR2_X2 U455 ( .A(n452), .B(n451), .ZN(n462) );
  NAND2_X1 U456 ( .A1(n501), .A2(n516), .ZN(n370) );
  NAND2_X1 U457 ( .A1(n675), .A2(n626), .ZN(n539) );
  NAND2_X1 U458 ( .A1(n538), .A2(n687), .ZN(n675) );
  NAND2_X1 U459 ( .A1(n521), .A2(n509), .ZN(n377) );
  NAND2_X1 U460 ( .A1(n372), .A2(G234), .ZN(n412) );
  NAND2_X1 U461 ( .A1(n372), .A2(G224), .ZN(n464) );
  NAND2_X1 U462 ( .A1(n372), .A2(G227), .ZN(n492) );
  OR2_X1 U463 ( .A1(n372), .A2(G952), .ZN(n647) );
  NAND2_X1 U464 ( .A1(n743), .A2(n372), .ZN(n749) );
  XNOR2_X2 U465 ( .A(n411), .B(G953), .ZN(n372) );
  NAND2_X1 U466 ( .A1(n405), .A2(n352), .ZN(n373) );
  INV_X1 U467 ( .A(n509), .ZN(n374) );
  NAND2_X1 U468 ( .A1(n376), .A2(n509), .ZN(n375) );
  NAND2_X1 U469 ( .A1(n392), .A2(n404), .ZN(n376) );
  NOR2_X1 U470 ( .A1(n559), .A2(n560), .ZN(n379) );
  INV_X1 U471 ( .A(n575), .ZN(n380) );
  NAND2_X1 U472 ( .A1(n559), .A2(n560), .ZN(n382) );
  NAND2_X1 U473 ( .A1(n575), .A2(n560), .ZN(n383) );
  XNOR2_X2 U474 ( .A(n558), .B(KEYINPUT0), .ZN(n575) );
  NAND2_X1 U475 ( .A1(n636), .A2(n511), .ZN(n513) );
  NAND2_X1 U476 ( .A1(n406), .A2(KEYINPUT41), .ZN(n399) );
  AND2_X1 U477 ( .A1(n406), .A2(n517), .ZN(n702) );
  OR2_X1 U478 ( .A1(n406), .A2(n517), .ZN(n704) );
  NAND2_X1 U479 ( .A1(n392), .A2(n505), .ZN(n522) );
  XNOR2_X2 U480 ( .A(n393), .B(n457), .ZN(n531) );
  XNOR2_X1 U481 ( .A(n462), .B(n456), .ZN(n394) );
  XNOR2_X2 U482 ( .A(n447), .B(n446), .ZN(n742) );
  NOR2_X1 U483 ( .A1(n514), .A2(n524), .ZN(n395) );
  NAND2_X1 U484 ( .A1(n398), .A2(n401), .ZN(n685) );
  NAND2_X1 U485 ( .A1(n402), .A2(KEYINPUT41), .ZN(n400) );
  NAND2_X1 U486 ( .A1(n403), .A2(n701), .ZN(n402) );
  NAND2_X1 U487 ( .A1(n356), .A2(n403), .ZN(n401) );
  NAND2_X1 U488 ( .A1(n508), .A2(n597), .ZN(n407) );
  INV_X1 U489 ( .A(n518), .ZN(n408) );
  XNOR2_X2 U490 ( .A(n535), .B(KEYINPUT19), .ZN(n518) );
  XNOR2_X2 U491 ( .A(n420), .B(n419), .ZN(n465) );
  BUF_X1 U492 ( .A(n575), .Z(n591) );
  XNOR2_X2 U493 ( .A(G119), .B(G116), .ZN(n449) );
  XNOR2_X2 U494 ( .A(KEYINPUT67), .B(KEYINPUT83), .ZN(n448) );
  BUF_X1 U495 ( .A(n609), .Z(n730) );
  OR2_X1 U496 ( .A1(n557), .A2(n556), .ZN(n409) );
  AND2_X1 U497 ( .A1(n609), .A2(n679), .ZN(n610) );
  INV_X1 U498 ( .A(G137), .ZN(n426) );
  XNOR2_X1 U499 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U500 ( .A(n497), .B(n496), .ZN(n498) );
  NAND2_X1 U501 ( .A1(n687), .A2(n572), .ZN(n573) );
  XNOR2_X1 U502 ( .A(n416), .B(n415), .ZN(n417) );
  AND2_X1 U503 ( .A1(n589), .A2(n507), .ZN(n508) );
  INV_X2 U504 ( .A(KEYINPUT64), .ZN(n411) );
  XOR2_X1 U505 ( .A(KEYINPUT8), .B(n412), .Z(n430) );
  NAND2_X1 U506 ( .A1(G217), .A2(n430), .ZN(n418) );
  XOR2_X1 U507 ( .A(KEYINPUT9), .B(G116), .Z(n414) );
  XNOR2_X1 U508 ( .A(G122), .B(G107), .ZN(n413) );
  XNOR2_X1 U509 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U510 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n415) );
  XNOR2_X1 U511 ( .A(n418), .B(n417), .ZN(n422) );
  XNOR2_X2 U512 ( .A(KEYINPUT72), .B(G143), .ZN(n420) );
  INV_X1 U513 ( .A(n447), .ZN(n421) );
  XNOR2_X1 U514 ( .A(n422), .B(n421), .ZN(n616) );
  XOR2_X1 U515 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n424) );
  XNOR2_X1 U516 ( .A(KEYINPUT75), .B(KEYINPUT24), .ZN(n423) );
  XNOR2_X1 U517 ( .A(G110), .B(G119), .ZN(n425) );
  XNOR2_X1 U518 ( .A(n425), .B(KEYINPUT23), .ZN(n429) );
  NAND2_X1 U519 ( .A1(G221), .A2(n430), .ZN(n431) );
  NOR2_X1 U520 ( .A1(n725), .A2(G902), .ZN(n436) );
  XNOR2_X1 U521 ( .A(G902), .B(KEYINPUT15), .ZN(n611) );
  NAND2_X1 U522 ( .A1(G234), .A2(n611), .ZN(n432) );
  XNOR2_X1 U523 ( .A(KEYINPUT20), .B(n432), .ZN(n437) );
  NAND2_X1 U524 ( .A1(n437), .A2(G217), .ZN(n434) );
  XNOR2_X1 U525 ( .A(KEYINPUT25), .B(KEYINPUT71), .ZN(n433) );
  XNOR2_X1 U526 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U527 ( .A(n436), .B(n435), .ZN(n571) );
  NAND2_X1 U528 ( .A1(G221), .A2(n437), .ZN(n438) );
  XNOR2_X1 U529 ( .A(n438), .B(KEYINPUT21), .ZN(n690) );
  NAND2_X1 U530 ( .A1(G237), .A2(G234), .ZN(n439) );
  XNOR2_X1 U531 ( .A(n439), .B(KEYINPUT14), .ZN(n441) );
  NAND2_X1 U532 ( .A1(G952), .A2(n441), .ZN(n440) );
  XOR2_X1 U533 ( .A(KEYINPUT85), .B(n440), .Z(n714) );
  NOR2_X1 U534 ( .A1(n714), .A2(G953), .ZN(n557) );
  AND2_X1 U535 ( .A1(G902), .A2(n441), .ZN(n554) );
  AND2_X1 U536 ( .A1(n554), .A2(n357), .ZN(n442) );
  NOR2_X1 U537 ( .A1(n557), .A2(n442), .ZN(n504) );
  NOR2_X1 U538 ( .A1(n690), .A2(n504), .ZN(n443) );
  XNOR2_X1 U539 ( .A(KEYINPUT66), .B(n443), .ZN(n444) );
  NAND2_X1 U540 ( .A1(n571), .A2(n444), .ZN(n530) );
  XNOR2_X1 U541 ( .A(KEYINPUT4), .B(G146), .ZN(n463) );
  XNOR2_X1 U542 ( .A(G137), .B(G131), .ZN(n445) );
  XNOR2_X1 U543 ( .A(n463), .B(n445), .ZN(n446) );
  XNOR2_X2 U544 ( .A(G113), .B(G101), .ZN(n450) );
  NAND2_X1 U545 ( .A1(n481), .A2(G210), .ZN(n453) );
  XNOR2_X1 U546 ( .A(n453), .B(KEYINPUT5), .ZN(n455) );
  XNOR2_X1 U547 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n454) );
  XNOR2_X1 U548 ( .A(n455), .B(n454), .ZN(n456) );
  INV_X1 U549 ( .A(G472), .ZN(n457) );
  XNOR2_X1 U550 ( .A(n458), .B(KEYINPUT28), .ZN(n516) );
  XNOR2_X1 U551 ( .A(G122), .B(G104), .ZN(n459) );
  XNOR2_X1 U552 ( .A(n459), .B(KEYINPUT16), .ZN(n460) );
  XNOR2_X1 U553 ( .A(G110), .B(G107), .ZN(n495) );
  XNOR2_X1 U554 ( .A(n460), .B(n495), .ZN(n461) );
  XNOR2_X1 U555 ( .A(n464), .B(n463), .ZN(n467) );
  XNOR2_X1 U556 ( .A(n465), .B(n410), .ZN(n466) );
  XNOR2_X1 U557 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U558 ( .A(n737), .B(n468), .ZN(n632) );
  INV_X1 U559 ( .A(n611), .ZN(n469) );
  OR2_X2 U560 ( .A1(n632), .A2(n469), .ZN(n472) );
  INV_X1 U561 ( .A(G902), .ZN(n487) );
  NAND2_X1 U562 ( .A1(n487), .A2(n470), .ZN(n473) );
  NAND2_X1 U563 ( .A1(n473), .A2(G210), .ZN(n471) );
  XNOR2_X2 U564 ( .A(n472), .B(n471), .ZN(n526) );
  AND2_X1 U565 ( .A1(n473), .A2(G214), .ZN(n517) );
  INV_X1 U566 ( .A(n517), .ZN(n701) );
  NAND2_X1 U567 ( .A1(n616), .A2(n487), .ZN(n476) );
  INV_X1 U568 ( .A(KEYINPUT100), .ZN(n474) );
  XNOR2_X1 U569 ( .A(n474), .B(G478), .ZN(n475) );
  XNOR2_X2 U570 ( .A(n476), .B(n475), .ZN(n524) );
  XOR2_X1 U571 ( .A(KEYINPUT11), .B(G113), .Z(n478) );
  XNOR2_X1 U572 ( .A(n350), .B(G131), .ZN(n477) );
  XNOR2_X1 U573 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U574 ( .A(n480), .B(n479), .ZN(n486) );
  NAND2_X1 U575 ( .A1(n481), .A2(G214), .ZN(n482) );
  XNOR2_X1 U576 ( .A(n482), .B(KEYINPUT12), .ZN(n484) );
  XOR2_X1 U577 ( .A(n484), .B(n483), .Z(n485) );
  XNOR2_X1 U578 ( .A(n486), .B(n485), .ZN(n644) );
  NAND2_X1 U579 ( .A1(n644), .A2(n487), .ZN(n490) );
  XNOR2_X1 U580 ( .A(G475), .B(KEYINPUT13), .ZN(n488) );
  XOR2_X1 U581 ( .A(n488), .B(KEYINPUT97), .Z(n489) );
  NAND2_X1 U582 ( .A1(n524), .A2(n523), .ZN(n703) );
  XOR2_X1 U583 ( .A(G140), .B(KEYINPUT87), .Z(n493) );
  XNOR2_X1 U584 ( .A(n493), .B(n492), .ZN(n497) );
  XNOR2_X1 U585 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U586 ( .A(n742), .B(n498), .ZN(n619) );
  NOR2_X1 U587 ( .A1(n619), .A2(G902), .ZN(n500) );
  INV_X1 U588 ( .A(G469), .ZN(n499) );
  XNOR2_X2 U589 ( .A(n500), .B(n499), .ZN(n589) );
  XOR2_X1 U590 ( .A(n589), .B(KEYINPUT109), .Z(n515) );
  AND2_X1 U591 ( .A1(n685), .A2(n515), .ZN(n501) );
  INV_X1 U592 ( .A(n750), .ZN(n511) );
  INV_X1 U593 ( .A(n504), .ZN(n505) );
  INV_X1 U594 ( .A(n571), .ZN(n597) );
  INV_X1 U595 ( .A(KEYINPUT91), .ZN(n506) );
  XNOR2_X1 U596 ( .A(n690), .B(n506), .ZN(n570) );
  INV_X1 U597 ( .A(n570), .ZN(n507) );
  XOR2_X1 U598 ( .A(KEYINPUT69), .B(KEYINPUT39), .Z(n509) );
  INV_X1 U599 ( .A(KEYINPUT98), .ZN(n510) );
  XNOR2_X1 U600 ( .A(n523), .B(n510), .ZN(n514) );
  XNOR2_X1 U601 ( .A(n513), .B(n512), .ZN(n542) );
  INV_X1 U602 ( .A(n669), .ZN(n663) );
  NAND2_X1 U603 ( .A1(n665), .A2(n518), .ZN(n519) );
  OR2_X2 U604 ( .A1(n705), .A2(n519), .ZN(n520) );
  XNOR2_X1 U605 ( .A(n520), .B(KEYINPUT47), .ZN(n540) );
  OR2_X1 U606 ( .A1(n522), .A2(n521), .ZN(n529) );
  NOR2_X1 U607 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U608 ( .A(n525), .B(KEYINPUT106), .ZN(n577) );
  BUF_X1 U609 ( .A(n526), .Z(n527) );
  INV_X1 U610 ( .A(n527), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n577), .A2(n548), .ZN(n528) );
  OR2_X1 U612 ( .A1(n529), .A2(n528), .ZN(n626) );
  NOR2_X1 U613 ( .A1(n530), .A2(n663), .ZN(n534) );
  BUF_X2 U614 ( .A(n531), .Z(n593) );
  XNOR2_X1 U615 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n532) );
  INV_X1 U616 ( .A(n596), .ZN(n533) );
  NAND2_X1 U617 ( .A1(n534), .A2(n533), .ZN(n543) );
  XOR2_X1 U618 ( .A(KEYINPUT111), .B(KEYINPUT36), .Z(n536) );
  XNOR2_X1 U619 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X2 U620 ( .A(n589), .B(KEYINPUT1), .ZN(n687) );
  NOR2_X1 U621 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U622 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n546) );
  NOR2_X1 U623 ( .A1(n687), .A2(n543), .ZN(n544) );
  NAND2_X1 U624 ( .A1(n701), .A2(n544), .ZN(n545) );
  XOR2_X1 U625 ( .A(n546), .B(n545), .Z(n547) );
  NOR2_X1 U626 ( .A1(n548), .A2(n547), .ZN(n628) );
  INV_X1 U627 ( .A(n628), .ZN(n549) );
  INV_X1 U628 ( .A(n550), .ZN(n552) );
  NOR2_X1 U629 ( .A1(n552), .A2(n551), .ZN(n627) );
  NAND2_X1 U630 ( .A1(n679), .A2(KEYINPUT2), .ZN(n553) );
  XNOR2_X1 U631 ( .A(n553), .B(KEYINPUT77), .ZN(n608) );
  INV_X1 U632 ( .A(G953), .ZN(n729) );
  NOR2_X1 U633 ( .A1(G898), .A2(n729), .ZN(n736) );
  NAND2_X1 U634 ( .A1(n736), .A2(n554), .ZN(n555) );
  XOR2_X1 U635 ( .A(n555), .B(KEYINPUT86), .Z(n556) );
  NAND2_X1 U636 ( .A1(n518), .A2(n409), .ZN(n558) );
  OR2_X1 U637 ( .A1(n703), .A2(n570), .ZN(n559) );
  INV_X1 U638 ( .A(n687), .ZN(n562) );
  INV_X1 U639 ( .A(n597), .ZN(n689) );
  NAND2_X1 U640 ( .A1(n689), .A2(n596), .ZN(n561) );
  NOR2_X1 U641 ( .A1(n562), .A2(n561), .ZN(n563) );
  INV_X1 U642 ( .A(KEYINPUT32), .ZN(n564) );
  XNOR2_X2 U643 ( .A(n565), .B(n564), .ZN(n629) );
  NAND2_X1 U644 ( .A1(n689), .A2(n566), .ZN(n567) );
  NOR2_X1 U645 ( .A1(n687), .A2(n567), .ZN(n568) );
  AND2_X1 U646 ( .A1(n600), .A2(n568), .ZN(n658) );
  NOR2_X2 U647 ( .A1(n629), .A2(n658), .ZN(n569) );
  XNOR2_X1 U648 ( .A(n569), .B(KEYINPUT80), .ZN(n580) );
  XOR2_X1 U649 ( .A(KEYINPUT105), .B(KEYINPUT33), .Z(n574) );
  OR2_X1 U650 ( .A1(n571), .A2(n570), .ZN(n588) );
  XNOR2_X1 U651 ( .A(n576), .B(KEYINPUT34), .ZN(n578) );
  INV_X1 U652 ( .A(KEYINPUT35), .ZN(n579) );
  NAND2_X1 U653 ( .A1(n580), .A2(n751), .ZN(n583) );
  INV_X1 U654 ( .A(KEYINPUT68), .ZN(n581) );
  NOR2_X1 U655 ( .A1(n581), .A2(KEYINPUT44), .ZN(n582) );
  XNOR2_X1 U656 ( .A(n583), .B(n582), .ZN(n606) );
  NOR2_X1 U657 ( .A1(n588), .A2(n593), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n687), .A2(n584), .ZN(n697) );
  NOR2_X1 U659 ( .A1(n697), .A2(n591), .ZN(n587) );
  XOR2_X1 U660 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n585) );
  XOR2_X1 U661 ( .A(KEYINPUT95), .B(n585), .Z(n586) );
  XNOR2_X1 U662 ( .A(n587), .B(n586), .ZN(n672) );
  INV_X1 U663 ( .A(n588), .ZN(n686) );
  NAND2_X1 U664 ( .A1(n686), .A2(n589), .ZN(n590) );
  NOR2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U666 ( .A(KEYINPUT92), .B(n592), .Z(n594) );
  INV_X1 U667 ( .A(n593), .ZN(n692) );
  NOR2_X1 U668 ( .A1(n594), .A2(n692), .ZN(n654) );
  NOR2_X1 U669 ( .A1(n672), .A2(n654), .ZN(n595) );
  NOR2_X1 U670 ( .A1(n595), .A2(n705), .ZN(n604) );
  NAND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U672 ( .A1(n687), .A2(n598), .ZN(n599) );
  AND2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n651) );
  INV_X1 U674 ( .A(KEYINPUT44), .ZN(n601) );
  NOR2_X1 U675 ( .A1(n601), .A2(KEYINPUT68), .ZN(n602) );
  OR2_X1 U676 ( .A1(n651), .A2(n602), .ZN(n603) );
  NOR2_X1 U677 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT45), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n608), .A2(n730), .ZN(n677) );
  NOR2_X1 U681 ( .A1(n610), .A2(KEYINPUT2), .ZN(n612) );
  NOR2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n677), .A2(n613), .ZN(n614) );
  XNOR2_X2 U684 ( .A(n614), .B(KEYINPUT65), .ZN(n723) );
  NAND2_X1 U685 ( .A1(n723), .A2(G478), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n615), .B(n616), .ZN(n617) );
  AND2_X1 U687 ( .A1(n617), .A2(n647), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n618), .B(KEYINPUT122), .ZN(G63) );
  NAND2_X1 U689 ( .A1(n723), .A2(G469), .ZN(n623) );
  XNOR2_X1 U690 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n621) );
  XNOR2_X1 U691 ( .A(n619), .B(KEYINPUT57), .ZN(n620) );
  XNOR2_X1 U692 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U693 ( .A(n623), .B(n622), .ZN(n624) );
  INV_X1 U694 ( .A(n647), .ZN(n728) );
  NOR2_X2 U695 ( .A1(n624), .A2(n728), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n625), .B(KEYINPUT120), .ZN(G54) );
  XNOR2_X1 U697 ( .A(n626), .B(n350), .ZN(G45) );
  XOR2_X1 U698 ( .A(G134), .B(n627), .Z(G36) );
  XOR2_X1 U699 ( .A(G140), .B(n628), .Z(G42) );
  XOR2_X1 U700 ( .A(n629), .B(G119), .Z(G21) );
  XNOR2_X1 U701 ( .A(KEYINPUT73), .B(KEYINPUT54), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n630), .B(KEYINPUT55), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n633), .B(n360), .ZN(n634) );
  NOR2_X1 U704 ( .A1(n634), .A2(n728), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n635), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U706 ( .A(n636), .B(G131), .ZN(G33) );
  NAND2_X1 U707 ( .A1(n723), .A2(G472), .ZN(n640) );
  XOR2_X1 U708 ( .A(KEYINPUT82), .B(KEYINPUT62), .Z(n637) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(n641) );
  NAND2_X1 U711 ( .A1(n641), .A2(n647), .ZN(n643) );
  XOR2_X1 U712 ( .A(KEYINPUT81), .B(KEYINPUT63), .Z(n642) );
  XNOR2_X1 U713 ( .A(n643), .B(n642), .ZN(G57) );
  NAND2_X1 U714 ( .A1(n723), .A2(G475), .ZN(n646) );
  XOR2_X1 U715 ( .A(n644), .B(KEYINPUT59), .Z(n645) );
  XNOR2_X1 U716 ( .A(n646), .B(n645), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X1 U718 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(G60) );
  XOR2_X1 U720 ( .A(G101), .B(n651), .Z(G3) );
  NAND2_X1 U721 ( .A1(n654), .A2(n669), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n652), .B(KEYINPUT112), .ZN(n653) );
  XNOR2_X1 U723 ( .A(G104), .B(n653), .ZN(G6) );
  XOR2_X1 U724 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n656) );
  INV_X1 U725 ( .A(n659), .ZN(n671) );
  NAND2_X1 U726 ( .A1(n654), .A2(n671), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U728 ( .A(G107), .B(n657), .ZN(G9) );
  XOR2_X1 U729 ( .A(G110), .B(n658), .Z(G12) );
  AND2_X1 U730 ( .A1(n359), .A2(n665), .ZN(n661) );
  XNOR2_X1 U731 ( .A(KEYINPUT113), .B(KEYINPUT29), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(n662) );
  XOR2_X1 U733 ( .A(G128), .B(n662), .Z(G30) );
  AND2_X1 U734 ( .A1(n665), .A2(n664), .ZN(n667) );
  XNOR2_X1 U735 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U737 ( .A(G146), .B(n668), .ZN(G48) );
  NAND2_X1 U738 ( .A1(n672), .A2(n669), .ZN(n670) );
  XNOR2_X1 U739 ( .A(n670), .B(G113), .ZN(G15) );
  NAND2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U741 ( .A(n673), .B(G116), .ZN(G18) );
  XOR2_X1 U742 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n674) );
  XNOR2_X1 U743 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U744 ( .A(G125), .B(n676), .ZN(G27) );
  XNOR2_X1 U745 ( .A(KEYINPUT2), .B(KEYINPUT74), .ZN(n681) );
  NOR2_X1 U746 ( .A1(n730), .A2(n681), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n678), .B(KEYINPUT76), .ZN(n683) );
  BUF_X1 U748 ( .A(n679), .Z(n680) );
  NOR2_X1 U749 ( .A1(n680), .A2(n681), .ZN(n682) );
  NOR2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U751 ( .A1(n677), .A2(n684), .ZN(n720) );
  INV_X1 U752 ( .A(n685), .ZN(n716) );
  OR2_X1 U753 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U754 ( .A(n688), .B(KEYINPUT50), .ZN(n695) );
  NAND2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U756 ( .A(KEYINPUT49), .B(n691), .ZN(n693) );
  NOR2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U758 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U759 ( .A(n696), .B(KEYINPUT117), .Z(n698) );
  AND2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U761 ( .A(KEYINPUT51), .B(n699), .Z(n700) );
  NOR2_X1 U762 ( .A1(n716), .A2(n700), .ZN(n710) );
  NOR2_X1 U763 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U764 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U765 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U766 ( .A1(n708), .A2(n715), .ZN(n709) );
  NOR2_X1 U767 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U768 ( .A(n711), .B(KEYINPUT118), .ZN(n712) );
  XNOR2_X1 U769 ( .A(KEYINPUT52), .B(n712), .ZN(n713) );
  NOR2_X1 U770 ( .A1(n714), .A2(n713), .ZN(n718) );
  NOR2_X1 U771 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U772 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U773 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U774 ( .A1(n721), .A2(G953), .ZN(n722) );
  XNOR2_X1 U775 ( .A(n722), .B(KEYINPUT53), .ZN(G75) );
  BUF_X1 U776 ( .A(n723), .Z(n724) );
  NAND2_X1 U777 ( .A1(n724), .A2(G217), .ZN(n726) );
  XNOR2_X1 U778 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U779 ( .A1(n728), .A2(n727), .ZN(G66) );
  NAND2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n735) );
  XOR2_X1 U781 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n732) );
  NAND2_X1 U782 ( .A1(G224), .A2(G953), .ZN(n731) );
  XNOR2_X1 U783 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U784 ( .A1(n733), .A2(G898), .ZN(n734) );
  NAND2_X1 U785 ( .A1(n735), .A2(n734), .ZN(n739) );
  NOR2_X1 U786 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U787 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U788 ( .A(KEYINPUT124), .B(n740), .ZN(G69) );
  XNOR2_X1 U789 ( .A(n742), .B(n741), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n680), .B(n744), .ZN(n743) );
  XOR2_X1 U791 ( .A(G227), .B(n744), .Z(n745) );
  NAND2_X1 U792 ( .A1(n745), .A2(G900), .ZN(n746) );
  XOR2_X1 U793 ( .A(KEYINPUT125), .B(n746), .Z(n747) );
  NAND2_X1 U794 ( .A1(n747), .A2(G953), .ZN(n748) );
  NAND2_X1 U795 ( .A1(n749), .A2(n748), .ZN(G72) );
  XOR2_X1 U796 ( .A(n750), .B(G137), .Z(G39) );
  XNOR2_X1 U797 ( .A(G122), .B(KEYINPUT126), .ZN(n752) );
  XNOR2_X1 U798 ( .A(n752), .B(n751), .ZN(G24) );
endmodule

