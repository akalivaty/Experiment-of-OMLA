//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1217, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n218), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  NAND2_X1  g0051(.A1(new_n208), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n213), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT71), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G58), .ZN(new_n259));
  OR3_X1    g0059(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT8), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n207), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT72), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n255), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n207), .A2(G1), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n254), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G50), .ZN(new_n272));
  INV_X1    g0072(.A(G13), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G1), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G20), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n272), .B1(G50), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT78), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT9), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n279), .B1(new_n278), .B2(new_n280), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT10), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(KEYINPUT79), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n213), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT3), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT3), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G33), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G1698), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(G222), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT70), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(G1698), .ZN(new_n298));
  INV_X1    g0098(.A(G223), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n298), .A2(new_n299), .B1(new_n224), .B2(new_n294), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n289), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n213), .B2(new_n287), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT68), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT68), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G41), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n303), .B(new_n206), .C1(new_n308), .C2(G45), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n288), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g0112(.A(new_n312), .B(KEYINPUT69), .Z(new_n313));
  AOI21_X1  g0113(.A(new_n310), .B1(new_n313), .B2(G226), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n301), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n286), .B1(new_n316), .B2(G190), .ZN(new_n317));
  XOR2_X1   g0117(.A(KEYINPUT77), .B(G200), .Z(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n315), .A2(new_n319), .B1(new_n277), .B2(KEYINPUT9), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n284), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(KEYINPUT79), .A3(new_n285), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n285), .A2(KEYINPUT79), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n284), .A2(new_n323), .A3(new_n317), .A4(new_n320), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n277), .B1(new_n315), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(G179), .B2(new_n315), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n322), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n310), .B1(new_n313), .B2(G238), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  INV_X1    g0130(.A(G232), .ZN(new_n331));
  INV_X1    g0131(.A(G97), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n298), .A2(new_n331), .B1(new_n290), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n291), .A2(new_n293), .ZN(new_n334));
  INV_X1    g0134(.A(G226), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n334), .A2(new_n335), .A3(G1698), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n289), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n329), .A2(new_n330), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n330), .B1(new_n329), .B2(new_n337), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT14), .B1(new_n341), .B2(new_n325), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(G179), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(G169), .C1(new_n339), .C2(new_n340), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT80), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n275), .A2(KEYINPUT74), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n273), .A2(new_n207), .A3(G1), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT74), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n255), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n270), .A2(new_n218), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n347), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR4_X1   g0156(.A1(new_n353), .A2(KEYINPUT80), .A3(new_n218), .A4(new_n270), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT12), .ZN(new_n358));
  INV_X1    g0158(.A(new_n352), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(new_n218), .ZN(new_n360));
  AND4_X1   g0160(.A1(new_n358), .A2(new_n274), .A3(G20), .A4(new_n218), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n356), .A2(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n265), .A2(G77), .ZN(new_n363));
  INV_X1    g0163(.A(new_n267), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n363), .B1(new_n207), .B2(G68), .C1(new_n202), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n254), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n366), .A2(KEYINPUT11), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(KEYINPUT11), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n362), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n346), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(G200), .B1(new_n339), .B2(new_n340), .ZN(new_n372));
  INV_X1    g0172(.A(new_n340), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n373), .A2(G190), .A3(new_n338), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n369), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n261), .A2(new_n275), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n271), .B2(new_n261), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n259), .A2(new_n218), .ZN(new_n379));
  OAI21_X1  g0179(.A(G20), .B1(new_n379), .B2(new_n201), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n267), .A2(G159), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n290), .A2(KEYINPUT81), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT81), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G33), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n387), .A3(KEYINPUT3), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n292), .A2(KEYINPUT82), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT82), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n391), .A3(G33), .ZN(new_n392));
  AOI21_X1  g0192(.A(G20), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  OAI21_X1  g0194(.A(G68), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(KEYINPUT83), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT83), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT7), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI211_X1 g0199(.A(G20), .B(new_n399), .C1(new_n388), .C2(new_n392), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n384), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n254), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n394), .A2(G20), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n389), .A2(new_n391), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n290), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n385), .A2(new_n387), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n292), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n399), .B1(new_n207), .B2(new_n334), .ZN(new_n410));
  OAI21_X1  g0210(.A(G68), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n382), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT16), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n378), .B1(new_n402), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  NOR2_X1   g0215(.A1(G223), .A2(G1698), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n335), .B2(G1698), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n388), .A2(new_n417), .A3(new_n392), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n289), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n288), .A2(G232), .A3(new_n311), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n309), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(G179), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n288), .B1(new_n418), .B2(new_n419), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n309), .A2(new_n422), .ZN(new_n426));
  OAI21_X1  g0226(.A(G169), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n414), .A2(new_n415), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n415), .B1(new_n414), .B2(new_n428), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(G190), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n421), .A2(new_n432), .A3(new_n423), .ZN(new_n433));
  INV_X1    g0233(.A(G200), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n425), .B2(new_n426), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n436), .B(new_n378), .C1(new_n402), .C2(new_n413), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n438), .A2(KEYINPUT84), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(KEYINPUT84), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n437), .B2(new_n440), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n431), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n312), .B(KEYINPUT69), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n309), .B1(new_n444), .B2(new_n225), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT73), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n298), .A2(new_n219), .B1(new_n226), .B2(new_n294), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n334), .A2(new_n331), .A3(G1698), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n289), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n445), .A2(new_n446), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n447), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n452), .A2(new_n432), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n353), .A2(new_n224), .A3(new_n270), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n454), .B(KEYINPUT75), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G20), .A2(G77), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT15), .B(G87), .ZN(new_n457));
  OAI221_X1 g0257(.A(new_n456), .B1(new_n256), .B2(new_n364), .C1(new_n263), .C2(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n224), .A2(new_n359), .B1(new_n458), .B2(new_n254), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT76), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n452), .A2(new_n319), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n455), .A2(KEYINPUT76), .A3(new_n459), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n453), .A2(new_n462), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n452), .A2(G179), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n452), .A2(new_n325), .B1(new_n455), .B2(new_n459), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NOR4_X1   g0269(.A1(new_n328), .A2(new_n376), .A3(new_n443), .A4(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n388), .A2(new_n392), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(new_n207), .A3(G68), .ZN(new_n472));
  NOR3_X1   g0272(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT87), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n207), .B1(new_n290), .B2(new_n332), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(KEYINPUT19), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n263), .A2(new_n332), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n472), .B(new_n476), .C1(KEYINPUT19), .C2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(new_n254), .B1(new_n359), .B2(new_n457), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n255), .B(new_n275), .C1(G1), .C2(new_n290), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT88), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n388), .A2(new_n392), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n225), .A2(G1698), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(G238), .B2(G1698), .ZN(new_n488));
  INV_X1    g0288(.A(G116), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT81), .B(G33), .ZN(new_n490));
  OAI22_X1  g0290(.A1(new_n486), .A2(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n289), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n206), .A2(G45), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n221), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n494), .B(new_n288), .C1(G274), .C2(new_n493), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n318), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n484), .A2(new_n485), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(G190), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT88), .B1(new_n483), .B2(new_n498), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n294), .A2(KEYINPUT4), .A3(G244), .A4(new_n295), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n294), .A2(G250), .A3(G1698), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n295), .A2(G244), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n486), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n288), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT5), .B1(new_n305), .B2(new_n307), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT5), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n206), .B(G45), .C1(new_n513), .C2(G41), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n288), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n511), .B1(G257), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n512), .A2(new_n514), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n303), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n275), .A2(G97), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n481), .B2(G97), .ZN(new_n523));
  XNOR2_X1  g0323(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n524));
  OAI22_X1  g0324(.A1(KEYINPUT3), .A2(new_n490), .B1(new_n524), .B2(G33), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n403), .ZN(new_n526));
  INV_X1    g0326(.A(new_n410), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n226), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT6), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n529), .A2(new_n332), .A3(G107), .ZN(new_n530));
  XNOR2_X1  g0330(.A(G97), .B(G107), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(new_n529), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n532), .A2(new_n207), .B1(new_n224), .B2(new_n364), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n254), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n523), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT85), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n523), .A2(new_n534), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT85), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n517), .A2(G190), .A3(new_n519), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n521), .A2(new_n536), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n517), .A2(G179), .A3(new_n519), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n325), .B1(new_n517), .B2(new_n519), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n535), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n496), .A2(new_n325), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n479), .B1(new_n457), .B2(new_n480), .ZN(new_n546));
  INV_X1    g0346(.A(G179), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n497), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n548), .A2(KEYINPUT86), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(KEYINPUT86), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n545), .B(new_n546), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n503), .A2(new_n541), .A3(new_n544), .A4(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT89), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n227), .A2(G1698), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n471), .B(new_n557), .C1(G257), .C2(G1698), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n334), .A2(G303), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n288), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G270), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n519), .B1(new_n561), .B2(new_n515), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(new_n325), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n505), .B(new_n207), .C1(G33), .C2(new_n332), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n254), .B(new_n565), .C1(new_n207), .C2(G116), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT20), .ZN(new_n567));
  OR3_X1    g0367(.A1(new_n566), .A2(KEYINPUT90), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT90), .B1(new_n566), .B2(new_n567), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n567), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n489), .B1(new_n206), .B2(G33), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n354), .A2(new_n572), .B1(new_n489), .B2(new_n359), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n564), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT91), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT21), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT21), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n560), .A2(new_n562), .A3(new_n547), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n221), .A2(new_n295), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n471), .B(new_n584), .C1(G257), .C2(new_n295), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n407), .A2(G294), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n288), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n519), .B1(new_n227), .B2(new_n515), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(new_n434), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(G190), .B2(new_n589), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT22), .ZN(new_n592));
  NOR4_X1   g0392(.A1(new_n486), .A2(new_n592), .A3(G20), .A4(new_n220), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n207), .A2(G87), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n592), .B1(new_n334), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n407), .A2(new_n207), .A3(G116), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT92), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n597), .A2(KEYINPUT23), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(KEYINPUT23), .ZN(new_n599));
  OAI211_X1 g0399(.A(G20), .B(new_n226), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n597), .A2(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n595), .A2(new_n596), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  OR3_X1    g0402(.A1(new_n593), .A2(KEYINPUT24), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT24), .B1(new_n593), .B2(new_n602), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n255), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n480), .A2(new_n226), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n349), .A2(new_n226), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n607), .B(KEYINPUT25), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n591), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n563), .A2(new_n434), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(G190), .B2(new_n563), .ZN(new_n612));
  INV_X1    g0412(.A(new_n574), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n589), .A2(new_n547), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(G169), .B2(new_n589), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  NOR4_X1   g0417(.A1(new_n583), .A2(new_n610), .A3(new_n614), .A4(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n556), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n470), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g0421(.A(new_n621), .B(KEYINPUT93), .Z(G372));
  INV_X1    g0422(.A(new_n442), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n375), .A2(new_n466), .A3(new_n467), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n371), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n431), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n322), .B(new_n324), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n627), .A2(new_n327), .ZN(new_n628));
  INV_X1    g0428(.A(new_n470), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n591), .A2(new_n609), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n484), .A2(new_n499), .A3(new_n501), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n544), .A2(new_n541), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n577), .A2(KEYINPUT21), .B1(new_n574), .B2(new_n581), .ZN(new_n633));
  INV_X1    g0433(.A(new_n617), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n580), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n546), .A2(new_n545), .A3(new_n548), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n520), .A2(G169), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n517), .A2(G179), .A3(new_n519), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n537), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n503), .A2(new_n641), .A3(new_n551), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT26), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n631), .A2(new_n637), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n639), .A2(new_n640), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n539), .A2(new_n536), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n644), .A2(new_n645), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n638), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n628), .B1(new_n629), .B2(new_n650), .ZN(G369));
  NAND2_X1  g0451(.A1(new_n274), .A2(new_n207), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT94), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT27), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n653), .B1(new_n652), .B2(KEYINPUT27), .ZN(new_n655));
  OAI221_X1 g0455(.A(G213), .B1(KEYINPUT27), .B2(new_n652), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n617), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n609), .A2(new_n659), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n610), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n660), .B1(new_n662), .B2(new_n617), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n574), .A2(new_n658), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n583), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n633), .A2(new_n580), .A3(new_n665), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n614), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(KEYINPUT95), .A3(G330), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT95), .B1(new_n669), .B2(G330), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n664), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n662), .A2(new_n583), .A3(new_n634), .A4(new_n659), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n660), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT96), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT96), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n677), .A3(new_n660), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n673), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n210), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n308), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n474), .A2(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n216), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT97), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n643), .A2(new_n648), .ZN(new_n689));
  INV_X1    g0489(.A(new_n637), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n632), .B2(new_n635), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n658), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n688), .B1(new_n692), .B2(KEYINPUT29), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n659), .B1(new_n638), .B2(new_n649), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT29), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(KEYINPUT97), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n642), .A2(KEYINPUT26), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(KEYINPUT26), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n658), .B1(new_n699), .B2(new_n691), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n693), .A2(new_n696), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G330), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n618), .B(new_n659), .C1(new_n554), .C2(new_n555), .ZN(new_n704));
  NOR4_X1   g0504(.A1(new_n563), .A2(new_n589), .A3(G179), .A4(new_n497), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n520), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n517), .A2(new_n497), .A3(new_n581), .A4(new_n589), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n707), .A2(new_n708), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n658), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT31), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n703), .B1(new_n704), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n702), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n687), .B1(new_n716), .B2(G1), .ZN(G364));
  NOR2_X1   g0517(.A1(new_n671), .A2(new_n672), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n273), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n206), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n682), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n718), .B(new_n723), .C1(G330), .C2(new_n669), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n253), .B1(G20), .B2(new_n325), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n207), .A2(new_n547), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G200), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G190), .ZN(new_n728));
  INV_X1    g0528(.A(G317), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT33), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n729), .A2(KEYINPUT33), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n727), .A2(new_n432), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G326), .ZN(new_n734));
  INV_X1    g0534(.A(G294), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n432), .A2(G179), .A3(G200), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n207), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n732), .B(new_n734), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n726), .A2(G190), .A3(new_n434), .ZN(new_n739));
  INV_X1    g0539(.A(G322), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n207), .A2(G179), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G190), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n741), .B1(G329), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n726), .A2(new_n743), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n294), .B1(new_n748), .B2(G311), .ZN(new_n749));
  INV_X1    g0549(.A(G303), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n319), .A2(G190), .A3(new_n742), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n746), .B(new_n749), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n319), .A2(new_n432), .A3(new_n742), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n738), .B(new_n752), .C1(G283), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n737), .A2(new_n332), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n745), .A2(G159), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(KEYINPUT32), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n334), .B1(new_n748), .B2(G77), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n758), .B(new_n759), .C1(new_n259), .C2(new_n739), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G50), .A2(new_n733), .B1(new_n728), .B2(G68), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(KEYINPUT32), .B2(new_n757), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n751), .A2(new_n220), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n753), .A2(new_n226), .ZN(new_n764));
  NOR4_X1   g0564(.A1(new_n760), .A2(new_n762), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n725), .B1(new_n755), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n210), .A2(new_n294), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT98), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n768), .A2(G355), .B1(new_n489), .B2(new_n681), .ZN(new_n769));
  INV_X1    g0569(.A(G45), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n250), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n681), .A2(new_n471), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G45), .B2(new_n216), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n769), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n725), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n723), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n777), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n766), .B(new_n779), .C1(new_n669), .C2(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n724), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  NOR2_X1   g0583(.A1(new_n468), .A2(new_n658), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n460), .A2(new_n658), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n465), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(new_n786), .B2(new_n468), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n692), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n692), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n722), .B1(new_n790), .B2(new_n715), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n715), .B2(new_n790), .ZN(new_n792));
  INV_X1    g0592(.A(new_n725), .ZN(new_n793));
  INV_X1    g0593(.A(new_n739), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G143), .B1(new_n748), .B2(G159), .ZN(new_n795));
  INV_X1    g0595(.A(new_n728), .ZN(new_n796));
  INV_X1    g0596(.A(G150), .ZN(new_n797));
  INV_X1    g0597(.A(G137), .ZN(new_n798));
  INV_X1    g0598(.A(new_n733), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n795), .B1(new_n796), .B2(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT34), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n486), .B1(G132), .B2(new_n745), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n259), .B2(new_n737), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n754), .A2(G68), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n202), .B2(new_n751), .ZN(new_n807));
  OR4_X1    g0607(.A1(new_n802), .A2(new_n803), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G283), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n796), .A2(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n756), .B(new_n810), .C1(G303), .C2(new_n733), .ZN(new_n811));
  INV_X1    g0611(.A(new_n751), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G107), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n754), .A2(G87), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n739), .A2(new_n735), .B1(new_n747), .B2(new_n489), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n294), .B(new_n815), .C1(G311), .C2(new_n745), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n811), .A2(new_n813), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n793), .B1(new_n808), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n725), .A2(new_n775), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n723), .B(new_n818), .C1(new_n224), .C2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n787), .B2(new_n776), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n792), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G384));
  INV_X1    g0623(.A(KEYINPUT104), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT102), .ZN(new_n825));
  INV_X1    g0625(.A(new_n378), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n412), .B1(new_n395), .B2(new_n400), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n383), .ZN(new_n828));
  INV_X1    g0628(.A(new_n399), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n486), .A2(new_n207), .A3(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n830), .B(G68), .C1(new_n394), .C2(new_n393), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n255), .B1(new_n831), .B2(new_n384), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n826), .B1(new_n828), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n656), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n428), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n437), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT101), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n414), .A2(new_n428), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n414), .A2(new_n834), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n437), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n837), .B1(new_n836), .B2(KEYINPUT37), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n825), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n836), .A2(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT101), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n847), .A2(KEYINPUT102), .A3(new_n842), .A4(new_n838), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n833), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n834), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n431), .B2(new_n442), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT38), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n855), .B(new_n852), .C1(new_n845), .C2(new_n848), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT103), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n852), .B1(new_n845), .B2(new_n848), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n859), .A2(KEYINPUT103), .A3(KEYINPUT38), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n824), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n784), .B(KEYINPUT99), .Z(new_n862));
  NAND2_X1  g0662(.A1(new_n789), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT100), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n375), .A2(new_n342), .A3(new_n343), .A4(new_n345), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n369), .A2(new_n659), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n376), .B2(new_n866), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n865), .A2(new_n864), .A3(new_n866), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n849), .A2(new_n853), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n855), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n859), .A2(KEYINPUT38), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(KEYINPUT103), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n860), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(KEYINPUT104), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n861), .A2(new_n873), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT39), .B1(new_n858), .B2(new_n860), .ZN(new_n881));
  INV_X1    g0681(.A(new_n371), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n659), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n856), .A2(KEYINPUT105), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT105), .ZN(new_n887));
  INV_X1    g0687(.A(new_n840), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n839), .A2(new_n840), .A3(new_n437), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n443), .A2(new_n888), .B1(new_n890), .B2(new_n842), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n887), .B1(new_n891), .B2(KEYINPUT38), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n885), .B(new_n886), .C1(new_n856), .C2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n881), .A2(new_n884), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n626), .A2(new_n656), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n880), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n693), .A2(new_n696), .A3(new_n701), .A4(new_n470), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n897), .A2(new_n628), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n896), .B(new_n898), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n868), .A2(new_n787), .A3(new_n869), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n704), .A2(new_n713), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n861), .A2(new_n879), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n885), .B1(new_n856), .B2(new_n892), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT40), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n903), .A2(new_n904), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n470), .A2(new_n901), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n911), .A2(new_n912), .A3(new_n703), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n899), .A2(new_n913), .B1(new_n206), .B2(new_n719), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n899), .B2(new_n913), .ZN(new_n915));
  INV_X1    g0715(.A(new_n532), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n489), .B(new_n215), .C1(new_n916), .C2(KEYINPUT35), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(KEYINPUT35), .B2(new_n916), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT36), .Z(new_n919));
  OR3_X1    g0719(.A1(new_n379), .A2(new_n216), .A3(new_n224), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n206), .B(G13), .C1(new_n920), .C2(new_n246), .ZN(new_n921));
  OR3_X1    g0721(.A1(new_n915), .A2(new_n919), .A3(new_n921), .ZN(G367));
  AOI21_X1  g0722(.A(new_n659), .B1(new_n539), .B2(new_n536), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n645), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(KEYINPUT106), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(KEYINPUT106), .ZN(new_n926));
  INV_X1    g0726(.A(new_n923), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n544), .A3(new_n541), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n583), .A2(new_n659), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n664), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT42), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n929), .A2(new_n617), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n658), .B1(new_n934), .B2(new_n544), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT43), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n484), .A2(new_n659), .ZN(new_n937));
  MUX2_X1   g0737(.A(new_n644), .B(new_n690), .S(new_n937), .Z(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n933), .A2(new_n935), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n936), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n929), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n673), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n682), .B(KEYINPUT41), .Z(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n667), .A2(new_n668), .ZN(new_n948));
  INV_X1    g0748(.A(new_n614), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(G330), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT95), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n952), .A2(new_n670), .A3(new_n663), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n663), .B1(new_n952), .B2(new_n670), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n931), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n670), .A3(new_n663), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n673), .A2(new_n930), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT108), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n716), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n943), .B1(new_n676), .B2(new_n678), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT45), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n676), .A2(new_n678), .A3(new_n943), .ZN(new_n965));
  XOR2_X1   g0765(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n965), .B(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n954), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n962), .B(KEYINPUT45), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n965), .B(new_n966), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n673), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n959), .B1(new_n716), .B2(new_n958), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n961), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n702), .A2(new_n715), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n947), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n945), .B1(new_n977), .B2(new_n720), .ZN(new_n978));
  INV_X1    g0778(.A(new_n772), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n241), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n778), .B1(new_n210), .B2(new_n457), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n722), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n754), .A2(G97), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n983), .B(new_n486), .C1(new_n729), .C2(new_n744), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT109), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n812), .A2(KEYINPUT46), .A3(G116), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT46), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n751), .B2(new_n489), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n739), .A2(new_n750), .B1(new_n747), .B2(new_n809), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G294), .B2(new_n728), .ZN(new_n990));
  INV_X1    g0790(.A(new_n737), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G107), .A2(new_n991), .B1(new_n733), .B2(G311), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n986), .A2(new_n988), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n737), .A2(new_n218), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(G143), .B2(new_n733), .ZN(new_n995));
  INV_X1    g0795(.A(G159), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n995), .B1(new_n996), .B2(new_n796), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n739), .A2(new_n797), .B1(new_n747), .B2(new_n202), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n334), .B(new_n998), .C1(G137), .C2(new_n745), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n754), .A2(G77), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n812), .A2(G58), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n985), .A2(new_n993), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT110), .Z(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT47), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n982), .B1(new_n1006), .B2(new_n725), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n939), .A2(new_n777), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n978), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(G387));
  NAND2_X1  g0811(.A1(new_n716), .A2(new_n958), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n976), .A2(new_n957), .A3(new_n955), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n682), .A3(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n737), .A2(new_n457), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n471), .B1(new_n202), .B2(new_n739), .C1(new_n797), .C2(new_n744), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(G159), .C2(new_n733), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n796), .A2(new_n261), .B1(new_n218), .B2(new_n747), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT111), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n812), .A2(G77), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1017), .A2(new_n983), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n471), .B1(G326), .B2(new_n745), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n751), .A2(new_n735), .B1(new_n737), .B2(new_n809), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n794), .A2(G317), .B1(new_n748), .B2(G303), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n728), .A2(G311), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(new_n740), .C2(new_n799), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT48), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n1027), .B2(new_n1026), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT49), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1022), .B1(new_n489), .B2(new_n753), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1021), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n723), .B1(new_n1033), .B2(new_n725), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n772), .B1(new_n237), .B2(new_n770), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n768), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1035), .B1(new_n684), .B2(new_n1036), .ZN(new_n1037));
  OR3_X1    g0837(.A1(new_n256), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1038));
  OAI21_X1  g0838(.A(KEYINPUT50), .B1(new_n256), .B2(G50), .ZN(new_n1039));
  AOI21_X1  g0839(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n684), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1037), .A2(new_n1041), .B1(new_n226), .B2(new_n681), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n778), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1034), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n663), .B2(new_n777), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n958), .B2(new_n721), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1014), .A2(new_n1046), .ZN(G393));
  NAND3_X1  g0847(.A1(new_n969), .A2(new_n972), .A3(new_n721), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n778), .B1(new_n332), .B2(new_n210), .C1(new_n979), .C2(new_n245), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n722), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G317), .A2(new_n733), .B1(new_n794), .B2(G311), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1051), .B(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n334), .B1(new_n747), .B2(new_n735), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G322), .B2(new_n745), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G116), .A2(new_n991), .B1(new_n728), .B2(G303), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n764), .B1(G283), .B2(new_n812), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G150), .A2(new_n733), .B1(new_n794), .B2(G159), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT51), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n747), .A2(new_n256), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n486), .B(new_n1061), .C1(G143), .C2(new_n745), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n812), .A2(G68), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n737), .A2(new_n224), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G50), .B2(new_n728), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1062), .A2(new_n814), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1058), .B1(new_n1060), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1050), .B1(new_n1067), .B2(new_n725), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n929), .B2(new_n780), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1048), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1012), .A2(KEYINPUT108), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1071), .A2(new_n960), .A3(new_n972), .A4(new_n969), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n683), .B1(new_n973), .B2(new_n1012), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1070), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(G390));
  NAND3_X1  g0875(.A1(new_n714), .A2(new_n787), .A3(new_n871), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n870), .B(KEYINPUT113), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n786), .A2(new_n468), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n784), .B1(new_n700), .B2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n883), .B(new_n906), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n872), .A2(new_n883), .B1(new_n881), .B2(new_n893), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1077), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1083), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n1076), .A3(new_n1081), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1084), .A2(new_n721), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n819), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1088), .A2(new_n262), .ZN(new_n1089));
  INV_X1    g0889(.A(G128), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n799), .A2(new_n1090), .B1(new_n996), .B2(new_n737), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G137), .B2(new_n728), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n745), .A2(G125), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n334), .B(new_n1093), .C1(G132), .C2(new_n794), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n754), .A2(G50), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT54), .B(G143), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT116), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n748), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1092), .A2(new_n1094), .A3(new_n1095), .A4(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n812), .A2(G150), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT53), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1064), .B1(G283), .B2(new_n733), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n226), .B2(new_n796), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n739), .A2(new_n489), .B1(new_n744), .B2(new_n735), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n294), .B(new_n1104), .C1(G97), .C2(new_n748), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n763), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n1106), .A3(new_n806), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1099), .A2(new_n1101), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n723), .B(new_n1089), .C1(new_n1108), .C2(new_n725), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n881), .A2(new_n893), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n776), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT114), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n714), .A2(new_n1112), .A3(new_n470), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n714), .B2(new_n470), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n897), .B(new_n628), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n714), .A2(new_n787), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1078), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n871), .B1(new_n714), .B2(new_n787), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n863), .B1(new_n1077), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1086), .A2(new_n1084), .A3(new_n1116), .A4(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(KEYINPUT115), .A3(new_n682), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1116), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1086), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1084), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT115), .B1(new_n1123), .B2(new_n682), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1087), .B(new_n1111), .C1(new_n1129), .C2(new_n1130), .ZN(G378));
  NOR2_X1   g0931(.A1(new_n277), .A2(new_n656), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT55), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n328), .B(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(G330), .B1(new_n907), .B2(new_n905), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n903), .B2(new_n904), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1136), .B1(new_n1138), .B2(KEYINPUT120), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT120), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1140), .B(new_n1137), .C1(new_n903), .C2(new_n904), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n903), .A2(new_n904), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1137), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1145), .A2(new_n1140), .A3(new_n1136), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n896), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1140), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1138), .A2(KEYINPUT120), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n1149), .A3(new_n1136), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n896), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1123), .A2(new_n1116), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1147), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT57), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1147), .A2(new_n1153), .A3(KEYINPUT57), .A4(new_n1154), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n682), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1147), .A2(new_n1153), .A3(new_n721), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n722), .B1(G50), .B2(new_n1088), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n728), .A2(G132), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n1090), .B2(new_n739), .C1(new_n798), .C2(new_n747), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G150), .A2(new_n991), .B1(new_n733), .B2(G125), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT117), .Z(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(new_n812), .C2(new_n1097), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT59), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G33), .B(G41), .C1(new_n745), .C2(G124), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n996), .B2(new_n753), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT118), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1169), .A2(new_n1170), .A3(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n471), .A2(new_n308), .ZN(new_n1175));
  AOI211_X1 g0975(.A(G50), .B(new_n1175), .C1(new_n290), .C2(new_n304), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n796), .A2(new_n332), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n994), .B(new_n1177), .C1(G116), .C2(new_n733), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n744), .A2(new_n809), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n739), .A2(new_n226), .B1(new_n747), .B2(new_n457), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(new_n812), .C2(G77), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n754), .A2(G58), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1178), .A2(new_n1181), .A3(new_n1175), .A4(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT58), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1176), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1174), .B(new_n1185), .C1(new_n1184), .C2(new_n1183), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1162), .B1(new_n1186), .B2(new_n725), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1136), .B2(new_n776), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1161), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1160), .A2(new_n1189), .ZN(G375));
  NAND3_X1  g0990(.A1(new_n1115), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1125), .A2(new_n947), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n751), .A2(new_n996), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G50), .A2(new_n991), .B1(new_n733), .B2(G132), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G150), .A2(new_n748), .B1(new_n745), .B2(G128), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(new_n798), .C2(new_n739), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1193), .B(new_n1196), .C1(new_n728), .C2(new_n1097), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1182), .A2(new_n471), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT121), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n799), .A2(new_n735), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1015), .B(new_n1200), .C1(G116), .C2(new_n728), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n294), .B1(new_n794), .B2(G283), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G107), .A2(new_n748), .B1(new_n745), .B2(G303), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1000), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G97), .B2(new_n812), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1197), .A2(new_n1199), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n722), .B1(G68), .B2(new_n1088), .C1(new_n1206), .C2(new_n793), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1078), .B2(new_n775), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1122), .B2(new_n721), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1192), .A2(new_n1209), .ZN(G381));
  INV_X1    g1010(.A(G375), .ZN(new_n1211));
  INV_X1    g1011(.A(G378), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1014), .A2(new_n782), .A3(new_n1046), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1074), .A2(new_n822), .A3(new_n1213), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(G387), .A2(G381), .A3(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1211), .A2(new_n1212), .A3(new_n1215), .ZN(G407));
  NAND2_X1  g1016(.A1(new_n657), .A2(G213), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1211), .A2(new_n1212), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(G407), .A2(new_n1219), .A3(G213), .ZN(G409));
  NOR3_X1   g1020(.A1(new_n978), .A2(KEYINPUT123), .A3(new_n1009), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT123), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n945), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n946), .B1(new_n1072), .B2(new_n716), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1223), .B1(new_n1224), .B2(new_n721), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1009), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1222), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n782), .B1(new_n1014), .B2(new_n1046), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1213), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(G390), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1074), .B1(new_n1213), .B2(new_n1228), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1221), .A2(new_n1227), .A3(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1229), .B(new_n1074), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT123), .B1(new_n978), .B2(new_n1009), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1225), .A2(new_n1222), .A3(new_n1226), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1234), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT125), .ZN(new_n1239));
  OAI211_X1 g1039(.A(G378), .B(new_n1189), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1161), .B(new_n1188), .C1(new_n1155), .C2(new_n946), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1212), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1217), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT60), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1191), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1125), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT122), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1246), .A2(KEYINPUT122), .A3(new_n1125), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1191), .A2(new_n1245), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1249), .A2(new_n682), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(G384), .A3(new_n1209), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G384), .B1(new_n1252), .B2(new_n1209), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G2897), .B(new_n1218), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1252), .A2(new_n1209), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n822), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1218), .A2(G2897), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1253), .A3(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1244), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1258), .A2(new_n1253), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1243), .A2(new_n1217), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT62), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1265), .A2(KEYINPUT62), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1239), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT124), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT63), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1263), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1243), .A2(new_n1217), .A3(new_n1272), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1218), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1265), .A2(new_n1271), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1270), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1238), .B1(new_n1277), .B2(new_n1272), .ZN(new_n1283));
  AND4_X1   g1083(.A1(new_n1270), .A2(new_n1262), .A3(new_n1283), .A4(new_n1281), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1269), .B1(new_n1282), .B2(new_n1284), .ZN(G405));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1240), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1263), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1264), .A2(new_n1240), .A3(new_n1286), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n1212), .A3(G375), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1288), .B(new_n1289), .C1(new_n1211), .C2(G378), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1291), .A2(new_n1238), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1238), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(G402));
endmodule


