//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G227), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G953), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G107), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT3), .A3(G104), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(G107), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT4), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G101), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT77), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n199), .A2(new_n203), .A3(new_n200), .A4(G101), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n195), .A2(G104), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n205), .B1(new_n194), .B2(new_n196), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT76), .B(G101), .Z(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n200), .B1(new_n199), .B2(G101), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n202), .A2(new_n204), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AND3_X1   g024(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NOR3_X1   g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT65), .B1(new_n215), .B2(G146), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n218), .B2(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n223), .A2(new_n218), .A3(G143), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT71), .B1(new_n222), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n222), .A2(KEYINPUT71), .A3(new_n229), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n210), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT66), .B1(new_n215), .B2(G146), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n215), .A2(G146), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n228), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n239));
  OAI21_X1  g053(.A(G128), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G128), .ZN(new_n242));
  OR2_X1    g056(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(new_n226), .A3(new_n228), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G101), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n195), .A2(G104), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n198), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(new_n206), .B2(new_n207), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n247), .A2(KEYINPUT78), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT78), .B1(new_n247), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n235), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  INV_X1    g071(.A(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT11), .A3(G134), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(G137), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n259), .A3(new_n263), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n251), .B(KEYINPUT79), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n268));
  OAI21_X1  g082(.A(G128), .B1(new_n268), .B2(new_n237), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n221), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n235), .B1(new_n270), .B2(new_n246), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n234), .A2(new_n254), .A3(new_n266), .A4(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n210), .A2(new_n233), .B1(new_n267), .B2(new_n271), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n266), .B1(new_n275), .B2(new_n254), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n191), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT12), .ZN(new_n278));
  INV_X1    g092(.A(new_n244), .ZN(new_n279));
  NOR2_X1   g093(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n242), .B1(new_n281), .B2(new_n225), .ZN(new_n282));
  INV_X1    g096(.A(new_n221), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n246), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(new_n251), .ZN(new_n285));
  OAI21_X1  g099(.A(G128), .B1(new_n279), .B2(new_n280), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n238), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n226), .A2(new_n228), .B1(new_n288), .B2(G128), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n251), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT78), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n247), .A2(KEYINPUT78), .A3(new_n251), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n285), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n265), .A2(KEYINPUT80), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n278), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n251), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(new_n270), .A3(new_n246), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n298), .B1(new_n252), .B2(new_n253), .ZN(new_n299));
  INV_X1    g113(.A(new_n295), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(KEYINPUT12), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n190), .A3(new_n273), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT82), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n277), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G469), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n302), .A2(KEYINPUT82), .A3(new_n190), .A4(new_n273), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n305), .A2(new_n306), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(G469), .A2(G902), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n190), .B1(new_n274), .B2(new_n276), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n294), .A2(new_n278), .A3(new_n295), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT12), .B1(new_n299), .B2(new_n300), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n273), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT81), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n317), .B(new_n273), .C1(new_n313), .C2(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n312), .B1(new_n319), .B2(new_n191), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n309), .B(new_n310), .C1(new_n320), .C2(new_n306), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT75), .B(G125), .Z(new_n322));
  INV_X1    g136(.A(KEYINPUT16), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(G125), .A2(G140), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n326), .B1(new_n322), .B2(G140), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(new_n327), .B2(new_n323), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n218), .ZN(new_n329));
  INV_X1    g143(.A(G237), .ZN(new_n330));
  INV_X1    g144(.A(G953), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(G214), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT88), .A3(G143), .ZN(new_n333));
  OR2_X1    g147(.A1(KEYINPUT88), .A2(G143), .ZN(new_n334));
  NOR2_X1   g148(.A1(G237), .A2(G953), .ZN(new_n335));
  NAND2_X1  g149(.A1(KEYINPUT88), .A2(G143), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n334), .A2(G214), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(G131), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT17), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n333), .A2(new_n337), .A3(G131), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(G146), .B(new_n325), .C1(new_n327), .C2(new_n323), .ZN(new_n343));
  INV_X1    g157(.A(new_n341), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT17), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n329), .A2(new_n342), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G125), .B(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n218), .ZN(new_n348));
  INV_X1    g162(.A(new_n327), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n348), .B1(new_n349), .B2(new_n218), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n344), .A2(KEYINPUT18), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n333), .A2(new_n337), .B1(KEYINPUT18), .B2(G131), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT89), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n352), .A2(new_n353), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n350), .B(new_n351), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G113), .B(G122), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT91), .B(G104), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n346), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n346), .B2(new_n356), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n307), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G475), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT20), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n346), .A2(new_n356), .A3(new_n360), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n347), .A2(KEYINPUT19), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT19), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n327), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n218), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n339), .A2(KEYINPUT90), .A3(new_n341), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT90), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n344), .B2(new_n338), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n370), .A2(new_n371), .A3(new_n373), .A4(new_n343), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n374), .A2(new_n356), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n366), .B1(new_n375), .B2(new_n360), .ZN(new_n376));
  NOR2_X1   g190(.A1(G475), .A2(G902), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(KEYINPUT92), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n365), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n360), .B1(new_n374), .B2(new_n356), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n365), .B(new_n378), .C1(new_n361), .C2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n364), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT13), .B1(new_n242), .B2(G143), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(new_n256), .ZN(new_n386));
  XNOR2_X1  g200(.A(G128), .B(G143), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G116), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G122), .ZN(new_n390));
  INV_X1    g204(.A(G122), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G116), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT93), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n393), .B1(new_n390), .B2(new_n392), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n195), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n395), .A2(new_n195), .A3(new_n396), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n388), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n387), .B(new_n256), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n390), .A2(KEYINPUT14), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n392), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n390), .A2(KEYINPUT14), .ZN(new_n404));
  OAI21_X1  g218(.A(G107), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n397), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT9), .B(G234), .Z(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G217), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n408), .A2(new_n409), .A3(G953), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n400), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n400), .B2(new_n406), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n307), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT15), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(G478), .ZN(new_n415));
  INV_X1    g229(.A(G478), .ZN(new_n416));
  OAI221_X1 g230(.A(new_n307), .B1(KEYINPUT15), .B2(new_n416), .C1(new_n411), .C2(new_n412), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n384), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G221), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n407), .B2(new_n307), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n321), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n335), .A2(G210), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(G101), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT28), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n222), .A2(KEYINPUT71), .A3(new_n229), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n265), .B1(new_n432), .B2(new_n230), .ZN(new_n433));
  INV_X1    g247(.A(new_n260), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n256), .A2(G137), .ZN(new_n435));
  OAI21_X1  g249(.A(G131), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n284), .A2(new_n264), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(KEYINPUT2), .A2(G113), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT68), .ZN(new_n440));
  NAND2_X1  g254(.A1(KEYINPUT2), .A2(G113), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n441), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT68), .B1(new_n443), .B2(new_n438), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  OR2_X1    g259(.A1(KEYINPUT69), .A2(G119), .ZN(new_n446));
  NAND2_X1  g260(.A1(KEYINPUT69), .A2(G119), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n389), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G119), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(G116), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT70), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  AND2_X1   g265(.A1(KEYINPUT69), .A2(G119), .ZN(new_n452));
  NOR2_X1   g266(.A1(KEYINPUT69), .A2(G119), .ZN(new_n453));
  OAI21_X1  g267(.A(G116), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT70), .ZN(new_n455));
  INV_X1    g269(.A(new_n450), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n445), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT72), .ZN(new_n459));
  NOR4_X1   g273(.A1(new_n448), .A2(new_n450), .A3(new_n438), .A4(new_n443), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n442), .A2(new_n444), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n455), .B1(new_n454), .B2(new_n456), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n460), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT72), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n433), .B(new_n437), .C1(new_n461), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n466), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n222), .A2(new_n229), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n266), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n436), .A2(new_n264), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n270), .B2(new_n246), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n469), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n431), .B1(new_n468), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n467), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT72), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n473), .B1(new_n233), .B2(new_n265), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT28), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n430), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n433), .A2(KEYINPUT30), .A3(new_n437), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n471), .B2(new_n473), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n469), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n468), .A3(new_n429), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT31), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT31), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n485), .A2(new_n488), .A3(new_n468), .A4(new_n429), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n481), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(G472), .A2(G902), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT73), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT32), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT32), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n433), .A2(new_n437), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n476), .A3(new_n477), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n468), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n480), .B1(new_n501), .B2(KEYINPUT28), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n429), .A2(KEYINPUT29), .ZN(new_n503));
  AOI21_X1  g317(.A(G902), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OR3_X1    g318(.A1(new_n475), .A2(new_n480), .A3(new_n430), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n505), .A2(KEYINPUT74), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n485), .A2(new_n468), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT29), .B1(new_n507), .B2(new_n430), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n505), .B2(KEYINPUT74), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n504), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G472), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n498), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT25), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n449), .A2(G128), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n452), .A2(new_n453), .ZN(new_n516));
  OAI211_X1 g330(.A(KEYINPUT23), .B(new_n515), .C1(new_n516), .C2(new_n242), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT23), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n518), .A3(new_n242), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(G110), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n446), .A2(new_n447), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n514), .B1(new_n521), .B2(G128), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT24), .B(G110), .Z(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n329), .B2(new_n343), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(G110), .B1(new_n517), .B2(new_n519), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n522), .A2(new_n523), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n343), .B(new_n348), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT22), .B(G137), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n331), .A2(G221), .A3(G234), .ZN(new_n532));
  XOR2_X1   g346(.A(new_n531), .B(new_n532), .Z(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n533), .ZN(new_n535));
  INV_X1    g349(.A(new_n530), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(new_n526), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n513), .B1(new_n538), .B2(G902), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT25), .A4(new_n307), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n409), .B1(G234), .B2(new_n307), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n538), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n542), .A2(G902), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n331), .A2(G952), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(G234), .B2(G237), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AOI211_X1 g365(.A(new_n307), .B(new_n331), .C1(G234), .C2(G237), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT21), .B(G898), .Z(new_n554));
  OAI21_X1  g368(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G214), .B1(G237), .B2(G902), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT85), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n470), .A2(new_n322), .ZN(new_n558));
  INV_X1    g372(.A(new_n322), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n270), .A2(new_n246), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n557), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n560), .A2(new_n557), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n331), .A2(G224), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n451), .A2(KEYINPUT5), .A3(new_n457), .ZN(new_n566));
  OAI21_X1  g380(.A(G113), .B1(new_n454), .B2(KEYINPUT5), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT83), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT83), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n566), .A2(new_n571), .A3(new_n568), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n570), .A2(new_n466), .A3(new_n267), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n210), .A2(new_n469), .ZN(new_n574));
  XNOR2_X1  g388(.A(G110), .B(G122), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(KEYINPUT84), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n573), .B2(new_n574), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n576), .B1(new_n579), .B2(KEYINPUT6), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT6), .ZN(new_n581));
  AOI211_X1 g395(.A(new_n581), .B(new_n578), .C1(new_n573), .C2(new_n574), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n565), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n575), .B(KEYINPUT8), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n454), .A2(KEYINPUT5), .A3(new_n456), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT86), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n567), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n460), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n584), .B1(new_n589), .B2(new_n297), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n566), .A2(new_n571), .A3(new_n568), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n571), .B1(new_n566), .B2(new_n568), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n591), .A2(new_n592), .A3(new_n460), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n590), .B1(new_n593), .B2(new_n297), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n560), .A2(new_n557), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT87), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT7), .B1(new_n564), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n596), .B2(new_n564), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n558), .A2(new_n560), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n595), .B(new_n598), .C1(new_n599), .C2(new_n557), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT7), .ZN(new_n601));
  INV_X1    g415(.A(new_n564), .ZN(new_n602));
  OAI22_X1  g416(.A1(new_n561), .A2(new_n562), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n594), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n605), .B2(new_n576), .ZN(new_n606));
  OAI21_X1  g420(.A(G210), .B1(G237), .B2(G902), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n583), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n607), .B1(new_n583), .B2(new_n606), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n555), .B(new_n556), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n425), .A2(new_n512), .A3(new_n548), .A4(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n613), .B(new_n207), .Z(G3));
  NAND2_X1  g428(.A1(new_n413), .A2(new_n416), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT95), .B1(new_n411), .B2(new_n412), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n307), .A2(G478), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n383), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n611), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n321), .A2(new_n424), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n490), .A2(new_n307), .ZN(new_n625));
  AOI22_X1  g439(.A1(KEYINPUT94), .A2(new_n492), .B1(new_n625), .B2(G472), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n625), .A2(KEYINPUT94), .A3(G472), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n623), .A2(new_n624), .A3(new_n548), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  INV_X1    g445(.A(new_n556), .ZN(new_n632));
  INV_X1    g446(.A(new_n610), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(new_n608), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n634), .A2(new_n321), .A3(new_n424), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n418), .B(new_n364), .C1(new_n379), .C2(new_n382), .ZN(new_n636));
  INV_X1    g450(.A(new_n555), .ZN(new_n637));
  OR3_X1    g451(.A1(new_n636), .A2(KEYINPUT96), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT96), .B1(new_n636), .B2(new_n637), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n547), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n635), .A2(new_n628), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NOR4_X1   g457(.A1(new_n526), .A2(new_n536), .A3(KEYINPUT36), .A4(new_n535), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n535), .A2(KEYINPUT36), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n527), .B2(new_n530), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n545), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n543), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n425), .A2(new_n612), .A3(new_n628), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  INV_X1    g466(.A(new_n649), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n498), .B2(new_n511), .ZN(new_n654));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n550), .B1(new_n552), .B2(new_n655), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n636), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT97), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n654), .A2(new_n635), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  XNOR2_X1  g474(.A(new_n656), .B(KEYINPUT39), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n321), .A2(new_n424), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n321), .A2(KEYINPUT99), .A3(new_n424), .A4(new_n662), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n666), .B1(new_n665), .B2(new_n667), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n307), .B1(new_n501), .B2(new_n429), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n430), .B1(new_n485), .B2(new_n468), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n498), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n609), .A2(new_n610), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n633), .A2(new_n608), .ZN(new_n678));
  INV_X1    g492(.A(new_n676), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR4_X1   g494(.A1(new_n649), .A2(new_n384), .A3(new_n632), .A4(new_n419), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n674), .A2(new_n677), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n669), .A2(new_n670), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n215), .ZN(G45));
  INV_X1    g498(.A(new_n656), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n621), .A2(new_n383), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n654), .A2(new_n635), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  AOI21_X1  g503(.A(new_n547), .B1(new_n498), .B2(new_n511), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT100), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n309), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n691), .A2(KEYINPUT100), .A3(G469), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n423), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n690), .A2(new_n623), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND4_X1  g513(.A1(new_n696), .A2(new_n512), .A3(new_n634), .A4(new_n640), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  NOR3_X1   g515(.A1(new_n653), .A2(new_n420), .A3(new_n637), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n696), .A2(new_n512), .A3(new_n634), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  NOR2_X1   g518(.A1(new_n384), .A2(new_n419), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n634), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n487), .B(new_n489), .C1(new_n502), .C2(new_n429), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n491), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT101), .B(G472), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n625), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n548), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n707), .A2(new_n696), .A3(new_n555), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  NAND3_X1  g529(.A1(new_n649), .A2(new_n711), .A3(new_n709), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT102), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n649), .A2(new_n711), .A3(KEYINPUT102), .A4(new_n709), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n686), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n621), .A2(KEYINPUT103), .A3(new_n383), .A4(new_n685), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n720), .A2(new_n696), .A3(new_n634), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  NAND2_X1  g540(.A1(new_n321), .A2(new_n424), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n321), .A2(KEYINPUT104), .A3(new_n424), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n675), .A2(new_n556), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT32), .B1(new_n490), .B2(new_n491), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT105), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n734), .A2(KEYINPUT105), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n490), .A2(KEYINPUT32), .A3(new_n491), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n511), .A2(new_n735), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n548), .A3(new_n724), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT42), .B1(new_n733), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n731), .B1(new_n727), .B2(new_n728), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT42), .B1(new_n722), .B2(new_n723), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n690), .A3(new_n730), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n263), .ZN(G33));
  NAND4_X1  g559(.A1(new_n741), .A2(new_n690), .A3(new_n658), .A4(new_n730), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT106), .B(G134), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G36));
  NAND2_X1  g562(.A1(new_n621), .A2(new_n384), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n621), .A2(new_n384), .A3(KEYINPUT43), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n653), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n626), .B2(new_n627), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n731), .B1(new_n754), .B2(new_n755), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n318), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n317), .B1(new_n302), .B2(new_n273), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n191), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n311), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n762), .B1(new_n761), .B2(new_n311), .ZN(new_n764));
  OAI211_X1 g578(.A(G469), .B(new_n763), .C1(new_n764), .C2(KEYINPUT107), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n320), .A2(new_n766), .A3(new_n762), .ZN(new_n767));
  OAI211_X1 g581(.A(KEYINPUT46), .B(new_n310), .C1(new_n765), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n309), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n764), .A2(KEYINPUT107), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n766), .B1(new_n320), .B2(new_n762), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n306), .B1(new_n320), .B2(new_n762), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT46), .B1(new_n773), .B2(new_n310), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n424), .B(new_n662), .C1(new_n769), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT108), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n310), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n309), .A3(new_n768), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n424), .A4(new_n662), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n758), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n258), .ZN(G39));
  OAI21_X1  g598(.A(new_n424), .B1(new_n769), .B2(new_n774), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT47), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n780), .A2(new_n787), .A3(new_n424), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n731), .A2(new_n656), .ZN(new_n789));
  INV_X1    g603(.A(new_n622), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n498), .A2(new_n511), .A3(new_n547), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n786), .A2(new_n788), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  NAND2_X1  g608(.A1(new_n694), .A2(new_n695), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT49), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n680), .A2(new_n677), .ZN(new_n797));
  INV_X1    g611(.A(new_n674), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n749), .A2(new_n547), .A3(new_n632), .A4(new_n423), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n740), .A2(new_n743), .A3(new_n746), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT109), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n636), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n611), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n624), .A3(new_n548), .A4(new_n628), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n613), .A2(new_n629), .A3(new_n650), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n714), .A2(new_n697), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n700), .A2(new_n703), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n720), .A2(new_n724), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n733), .A2(new_n810), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n512), .A2(new_n624), .A3(new_n421), .A4(new_n649), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n811), .B1(new_n789), .B2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n801), .A2(new_n808), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n654), .B(new_n635), .C1(new_n658), .C2(new_n687), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n649), .A2(new_n656), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n707), .A2(new_n674), .A3(new_n624), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n725), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT52), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n814), .A2(new_n815), .A3(new_n820), .ZN(new_n821));
  XOR2_X1   g635(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n816), .A2(new_n725), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT110), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT52), .A4(new_n818), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n819), .A2(KEYINPUT112), .A3(new_n822), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT110), .B1(new_n819), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n825), .A2(new_n828), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n714), .A2(new_n697), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n613), .A2(new_n629), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n650), .A2(new_n805), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n833), .A2(new_n809), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n740), .A2(new_n743), .A3(new_n746), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n812), .A2(new_n789), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n838), .B1(new_n810), .B2(new_n733), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT53), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n821), .B1(new_n841), .B2(KEYINPUT113), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n843), .B(KEYINPUT53), .C1(new_n832), .C2(new_n840), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT54), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n551), .B1(new_n751), .B2(new_n752), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n696), .A2(new_n846), .A3(new_n713), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n556), .B1(new_n680), .B2(new_n677), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(KEYINPUT50), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n851));
  INV_X1    g665(.A(new_n849), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n851), .B1(new_n852), .B2(new_n847), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n696), .A2(new_n732), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n498), .A2(new_n548), .A3(new_n550), .A4(new_n673), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT115), .B1(new_n855), .B2(new_n858), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n621), .A2(new_n383), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n856), .A2(new_n720), .A3(new_n846), .ZN(new_n864));
  AND4_X1   g678(.A1(KEYINPUT51), .A2(new_n854), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n786), .A2(new_n788), .B1(new_n423), .B2(new_n795), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n846), .A2(new_n732), .A3(new_n713), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n865), .B(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n786), .A2(new_n788), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n795), .A2(new_n423), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n854), .A2(new_n863), .A3(KEYINPUT51), .A4(new_n864), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT117), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n871), .B(KEYINPUT114), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n868), .B1(new_n870), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n854), .A2(new_n863), .A3(new_n864), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT116), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT116), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n882), .B(new_n876), .C1(new_n878), .C2(new_n879), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n860), .A2(new_n861), .A3(new_n790), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n549), .B1(new_n848), .B2(new_n634), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n856), .A2(new_n548), .A3(new_n738), .A4(new_n846), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT48), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT48), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND4_X1   g707(.A1(new_n875), .A2(new_n881), .A3(new_n883), .A4(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n832), .A2(new_n840), .A3(KEYINPUT53), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n815), .B1(new_n814), .B2(new_n820), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n845), .A2(new_n894), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(G952), .A2(G953), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n800), .B1(new_n900), .B2(new_n901), .ZN(G75));
  NOR2_X1   g716(.A1(new_n580), .A2(new_n582), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n565), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n897), .A2(G210), .A3(G902), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT119), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n897), .A2(KEYINPUT119), .A3(G210), .A4(G902), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n331), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n905), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(G51));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n895), .B2(new_n896), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n898), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n310), .B(KEYINPUT57), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n305), .B(new_n308), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n897), .A2(G902), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(new_n773), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n913), .B1(new_n921), .B2(new_n923), .ZN(G54));
  INV_X1    g738(.A(new_n913), .ZN(new_n925));
  AND4_X1   g739(.A1(KEYINPUT58), .A2(new_n897), .A3(G475), .A4(G902), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n376), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n376), .B2(new_n926), .ZN(G60));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT59), .Z(new_n930));
  NOR2_X1   g744(.A1(new_n619), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n898), .B2(new_n918), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n925), .ZN(new_n933));
  INV_X1    g747(.A(new_n930), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n814), .A2(new_n820), .A3(new_n815), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n832), .A2(new_n840), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n815), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n937), .B2(new_n843), .ZN(new_n938));
  INV_X1    g752(.A(new_n844), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n917), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n934), .B1(new_n940), .B2(new_n898), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n933), .B1(new_n941), .B2(new_n619), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT60), .Z(new_n944));
  NAND2_X1  g758(.A1(new_n897), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n647), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n925), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n945), .A2(new_n538), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n948), .A2(KEYINPUT61), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  INV_X1    g765(.A(new_n949), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(new_n947), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n950), .A2(new_n953), .ZN(G66));
  AOI21_X1  g768(.A(new_n331), .B1(new_n554), .B2(G224), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT121), .B1(new_n808), .B2(new_n809), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n700), .A2(new_n703), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT121), .ZN(new_n958));
  NOR4_X1   g772(.A1(new_n806), .A2(new_n807), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n955), .B1(new_n960), .B2(new_n331), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n903), .B1(G898), .B2(new_n331), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT122), .Z(new_n963));
  XNOR2_X1  g777(.A(new_n961), .B(new_n963), .ZN(G69));
  OAI21_X1  g778(.A(G953), .B1(new_n188), .B2(new_n655), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n482), .A2(new_n484), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n369), .B(KEYINPUT123), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n331), .A2(G900), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(KEYINPUT125), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n776), .A2(new_n782), .ZN(new_n973));
  INV_X1    g787(.A(new_n758), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n738), .A2(new_n707), .A3(new_n548), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n816), .A2(new_n725), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n837), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n975), .A2(new_n977), .A3(new_n793), .A4(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n972), .B1(new_n980), .B2(new_n331), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n971), .B1(new_n981), .B2(new_n970), .ZN(new_n982));
  AND4_X1   g796(.A1(new_n786), .A2(new_n788), .A3(new_n789), .A4(new_n792), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n983), .A2(new_n783), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n731), .B1(new_n622), .B2(new_n803), .ZN(new_n985));
  AND4_X1   g799(.A1(new_n690), .A2(new_n985), .A3(new_n665), .A4(new_n667), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT62), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n683), .B2(new_n978), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n670), .A2(new_n682), .ZN(new_n989));
  OAI211_X1 g803(.A(KEYINPUT62), .B(new_n826), .C1(new_n989), .C2(new_n669), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n986), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n984), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(new_n331), .A3(new_n969), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n982), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT124), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n966), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI211_X1 g810(.A(KEYINPUT124), .B(new_n965), .C1(new_n982), .C2(new_n993), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n996), .A2(new_n997), .ZN(G72));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n507), .A2(new_n429), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n956), .A2(new_n959), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n984), .A2(new_n1002), .A3(new_n977), .A4(new_n979), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  AOI21_X1  g819(.A(new_n1001), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n999), .B1(new_n1006), .B2(new_n913), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1005), .B1(new_n980), .B2(new_n960), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n1000), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1009), .A2(KEYINPUT127), .A3(new_n925), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n984), .A2(new_n1002), .A3(new_n991), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n1005), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n672), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(KEYINPUT126), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT126), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1013), .A2(new_n1016), .A3(new_n672), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n507), .A2(new_n430), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n486), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1005), .B(new_n1020), .C1(new_n842), .C2(new_n844), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n1011), .A2(new_n1018), .A3(new_n1021), .ZN(G57));
endmodule


