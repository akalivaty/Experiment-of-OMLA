//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1236, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT64), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n212), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n202), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n214), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n229), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n257));
  INV_X1    g0057(.A(G58), .ZN(new_n258));
  OR3_X1    g0058(.A1(new_n258), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n207), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n255), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n254), .B1(new_n206), .B2(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G50), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n269), .B1(G50), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT9), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT69), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT10), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n279), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n282), .A2(G226), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(G222), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n286), .B1(new_n220), .B2(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  AOI211_X1 g0089(.A(new_n280), .B(new_n283), .C1(new_n289), .C2(new_n277), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G190), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(KEYINPUT9), .B2(new_n272), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n275), .A2(new_n276), .A3(new_n295), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n292), .A2(new_n294), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT10), .B1(new_n297), .B2(new_n274), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n272), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(G169), .B2(new_n290), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n290), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT14), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n284), .A2(G226), .A3(new_n285), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n284), .A2(G232), .A3(G1698), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G97), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n277), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n280), .B1(G238), .B2(new_n282), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT13), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n314), .B1(new_n312), .B2(new_n313), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n307), .B(G169), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n312), .A2(new_n313), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT13), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n323), .A2(KEYINPUT70), .A3(new_n307), .A4(G169), .ZN(new_n324));
  OAI21_X1  g0124(.A(G169), .B1(new_n315), .B2(new_n316), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT14), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n315), .A2(new_n316), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G179), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n319), .A2(new_n324), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n265), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n330), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n262), .A2(new_n220), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n254), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT11), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n334), .ZN(new_n336));
  OR3_X1    g0136(.A1(new_n270), .A2(KEYINPUT12), .A3(G68), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT12), .B1(new_n270), .B2(G68), .ZN(new_n338));
  AOI22_X1  g0138(.A1(G68), .A2(new_n268), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n335), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n327), .B2(G190), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n293), .B2(new_n327), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G20), .A2(G77), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT15), .B(G87), .ZN(new_n346));
  OAI221_X1 g0146(.A(new_n345), .B1(new_n256), .B2(new_n330), .C1(new_n262), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n254), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n270), .A2(G77), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n268), .B2(G77), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n284), .A2(G232), .A3(new_n285), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n352), .B1(new_n222), .B2(new_n284), .C1(new_n287), .C2(new_n215), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n277), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n280), .B1(G244), .B2(new_n282), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n351), .B1(new_n357), .B2(G169), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n356), .A2(G179), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n356), .A2(G200), .ZN(new_n362));
  AOI22_X1  g0162(.A1(KEYINPUT68), .A2(new_n362), .B1(new_n357), .B2(G190), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n357), .A2(KEYINPUT68), .A3(G190), .ZN(new_n364));
  INV_X1    g0164(.A(new_n351), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n361), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n306), .A2(new_n344), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n260), .A2(new_n268), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(new_n270), .B2(new_n260), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT74), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G33), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT3), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT3), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G33), .ZN(new_n377));
  AOI21_X1  g0177(.A(G20), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT73), .B1(new_n378), .B2(KEYINPUT7), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT73), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n381), .C1(new_n284), .C2(G20), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT71), .B(KEYINPUT3), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n377), .B1(new_n384), .B2(G33), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G68), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n258), .A2(new_n214), .ZN(new_n389));
  OAI21_X1  g0189(.A(G20), .B1(new_n389), .B2(new_n201), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n265), .A2(G159), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n373), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n376), .A2(KEYINPUT71), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT71), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT3), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n397), .A3(G33), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n375), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(new_n381), .A3(new_n207), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G68), .ZN(new_n401));
  AOI21_X1  g0201(.A(G20), .B1(new_n398), .B2(new_n375), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n381), .ZN(new_n403));
  OAI211_X1 g0203(.A(KEYINPUT16), .B(new_n393), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n254), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n371), .B1(new_n394), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n214), .B1(new_n402), .B2(new_n381), .ZN(new_n407));
  INV_X1    g0207(.A(new_n375), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n384), .B2(G33), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT7), .B1(new_n409), .B2(G20), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n392), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n255), .B1(new_n411), .B2(KEYINPUT16), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n214), .B1(new_n383), .B2(new_n386), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n372), .B1(new_n413), .B2(new_n392), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(KEYINPUT74), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n370), .B1(new_n406), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G87), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n288), .A2(new_n285), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G226), .B2(new_n285), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n417), .B1(new_n399), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n277), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT75), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n280), .B1(G232), .B2(new_n282), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n420), .A2(KEYINPUT75), .A3(new_n277), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n423), .A2(new_n302), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n421), .A2(new_n424), .ZN(new_n427));
  INV_X1    g0227(.A(G169), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT76), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT76), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n426), .A2(new_n432), .A3(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT18), .B1(new_n416), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n370), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n412), .A2(KEYINPUT74), .A3(new_n414), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT74), .B1(new_n412), .B2(new_n414), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n426), .A2(new_n432), .A3(new_n429), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n432), .B1(new_n426), .B2(new_n429), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G190), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n423), .A2(new_n445), .A3(new_n424), .A4(new_n425), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n427), .A2(new_n293), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n436), .B(new_n448), .C1(new_n437), .C2(new_n438), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT17), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n406), .A2(new_n415), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(KEYINPUT17), .A3(new_n436), .A4(new_n448), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n435), .A2(new_n444), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n368), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n277), .ZN(new_n457));
  INV_X1    g0257(.A(G45), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G1), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n278), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n217), .B1(new_n458), .B2(G1), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(G238), .A2(G1698), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n221), .B2(G1698), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(new_n398), .A3(new_n375), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G116), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(G190), .B(new_n462), .C1(new_n467), .C2(new_n457), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n457), .B1(new_n465), .B2(new_n466), .ZN(new_n469));
  INV_X1    g0269(.A(new_n462), .ZN(new_n470));
  OAI21_X1  g0270(.A(G200), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n206), .A2(G33), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n270), .A2(new_n473), .A3(new_n229), .A4(new_n253), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n216), .ZN(new_n475));
  INV_X1    g0275(.A(new_n346), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(new_n270), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT19), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n207), .B1(new_n310), .B2(new_n478), .ZN(new_n479));
  NOR4_X1   g0279(.A1(KEYINPUT81), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  NOR2_X1   g0281(.A1(G87), .A2(G97), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(new_n222), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n479), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n398), .A2(new_n207), .A3(G68), .A4(new_n375), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n478), .B1(new_n262), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT82), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT82), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n489), .B(new_n478), .C1(new_n262), .C2(new_n486), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n484), .A2(new_n485), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  AOI211_X1 g0291(.A(new_n475), .B(new_n477), .C1(new_n491), .C2(new_n254), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n472), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n477), .B1(new_n491), .B2(new_n254), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT83), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n474), .A2(new_n346), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT80), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n462), .B1(new_n467), .B2(new_n457), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n428), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(G179), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI211_X1 g0303(.A(new_n477), .B(new_n496), .C1(new_n491), .C2(new_n254), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n469), .A2(new_n470), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n302), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n504), .A2(new_n495), .B1(new_n506), .B2(new_n499), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n493), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT84), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(KEYINPUT84), .B(new_n493), .C1(new_n503), .C2(new_n507), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(G41), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n459), .B(KEYINPUT78), .C1(KEYINPUT5), .C2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n206), .B(G45), .C1(new_n513), .C2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT78), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(G257), .A3(new_n457), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n515), .A2(new_n516), .B1(KEYINPUT5), .B2(new_n513), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n521), .A2(G274), .A3(new_n457), .A4(new_n514), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n221), .A2(G1698), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT4), .B1(new_n409), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT4), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(new_n221), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n284), .A2(new_n285), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G283), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n375), .A2(new_n377), .A3(G250), .A4(G1698), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n277), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n523), .A2(new_n302), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT79), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n536));
  INV_X1    g0336(.A(new_n524), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n526), .B1(new_n399), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n457), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n520), .A2(new_n522), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(KEYINPUT79), .A3(new_n302), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n222), .B1(new_n383), .B2(new_n386), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT6), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n545), .A2(new_n486), .A3(G107), .ZN(new_n546));
  XNOR2_X1  g0346(.A(G97), .B(G107), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n548), .A2(new_n207), .B1(new_n220), .B2(new_n330), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n254), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n474), .ZN(new_n551));
  INV_X1    g0351(.A(new_n270), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(KEYINPUT77), .A3(new_n486), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT77), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n270), .B2(G97), .ZN(new_n555));
  AOI22_X1  g0355(.A1(G97), .A2(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n523), .A2(new_n532), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n550), .A2(new_n556), .B1(new_n557), .B2(new_n428), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n523), .A2(G190), .A3(new_n532), .ZN(new_n559));
  OAI21_X1  g0359(.A(G200), .B1(new_n539), .B2(new_n540), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n550), .A2(new_n556), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n543), .A2(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  MUX2_X1   g0363(.A(G250), .B(G257), .S(G1698), .Z(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(new_n398), .A3(new_n375), .ZN(new_n565));
  XOR2_X1   g0365(.A(KEYINPUT87), .B(G294), .Z(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G33), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n277), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n519), .A2(G264), .A3(new_n457), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n522), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n293), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n569), .A2(new_n445), .A3(new_n522), .A4(new_n570), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT25), .B1(new_n552), .B2(new_n222), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT25), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n270), .A2(new_n576), .A3(G107), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n575), .A2(new_n577), .B1(new_n222), .B2(new_n474), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n375), .A2(new_n377), .A3(new_n207), .A4(G87), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT22), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n579), .A2(new_n580), .B1(G116), .B2(new_n263), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n216), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n398), .A2(new_n207), .A3(new_n375), .A4(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT86), .B1(new_n207), .B2(G107), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n584), .B(KEYINPUT23), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n581), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT24), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT24), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n581), .A2(new_n585), .A3(new_n588), .A4(new_n583), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n578), .B1(new_n590), .B2(new_n254), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n574), .A2(new_n591), .ZN(new_n592));
  AOI211_X1 g0392(.A(new_n223), .B(new_n277), .C1(new_n521), .C2(new_n514), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n457), .B1(new_n565), .B2(new_n567), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n302), .A3(new_n522), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n571), .A2(new_n428), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n255), .B1(new_n587), .B2(new_n589), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(new_n578), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n592), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G116), .ZN(new_n601));
  OR3_X1    g0401(.A1(new_n474), .A2(KEYINPUT85), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT85), .B1(new_n474), .B2(new_n601), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n529), .B(new_n207), .C1(G33), .C2(new_n486), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n601), .A2(G20), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n254), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n552), .A2(new_n601), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n604), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(G257), .A2(G1698), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n223), .B2(G1698), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(new_n398), .A3(new_n375), .ZN(new_n614));
  INV_X1    g0414(.A(new_n284), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G303), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n277), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n519), .A2(G270), .A3(new_n457), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n619), .A3(new_n522), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n611), .A2(new_n620), .A3(G169), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT21), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n620), .A2(G200), .ZN(new_n624));
  INV_X1    g0424(.A(new_n611), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n618), .A2(G190), .A3(new_n619), .A4(new_n522), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n618), .A2(G179), .A3(new_n619), .A4(new_n522), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n611), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n611), .A2(new_n620), .A3(KEYINPUT21), .A4(G169), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n623), .A2(new_n627), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n563), .A2(new_n600), .A3(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n456), .A2(new_n512), .A3(new_n633), .ZN(G372));
  NAND2_X1  g0434(.A1(new_n435), .A2(new_n444), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n329), .A2(new_n340), .B1(new_n343), .B2(new_n360), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n451), .A2(new_n453), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n304), .B1(new_n639), .B2(new_n299), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n543), .A2(new_n558), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n510), .A2(new_n642), .A3(new_n511), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n643), .A2(KEYINPUT26), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n599), .A2(new_n623), .A3(new_n630), .A4(new_n631), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n561), .A2(new_n562), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n574), .A2(new_n591), .B1(new_n472), .B2(new_n492), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n645), .A2(new_n641), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n505), .A2(G169), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n502), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n504), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n650), .A2(new_n651), .B1(new_n492), .B2(new_n472), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(new_n543), .A4(new_n558), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n648), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n644), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n640), .B1(new_n456), .B2(new_n657), .ZN(G369));
  NAND3_X1  g0458(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G343), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT88), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n600), .B1(new_n591), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n599), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n664), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT89), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n664), .A2(new_n611), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n632), .A2(new_n671), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n623), .A2(new_n630), .A3(new_n631), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n672), .B1(new_n673), .B2(new_n671), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n673), .A2(new_n664), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n669), .A2(KEYINPUT89), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT89), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n666), .B2(new_n668), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n678), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n599), .A2(new_n664), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n677), .A2(new_n682), .A3(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n210), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OR3_X1    g0488(.A1(new_n480), .A2(new_n483), .A3(G116), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n688), .A2(G1), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n228), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n688), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n643), .A2(KEYINPUT26), .ZN(new_n695));
  INV_X1    g0495(.A(new_n653), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT26), .B1(new_n696), .B2(new_n641), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(new_n648), .A3(new_n652), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n664), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n665), .B1(new_n644), .B2(new_n656), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT91), .ZN(new_n703));
  INV_X1    g0503(.A(new_n656), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n643), .A2(KEYINPUT26), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n664), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT91), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT92), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT92), .ZN(new_n712));
  AOI211_X1 g0512(.A(new_n712), .B(KEYINPUT29), .C1(new_n703), .C2(new_n708), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n701), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n563), .A2(new_n632), .A3(new_n600), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(new_n510), .A3(new_n511), .A4(new_n665), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n571), .A2(new_n302), .A3(new_n500), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT90), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n718), .A3(new_n620), .A4(new_n557), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n523), .A2(new_n595), .A3(new_n505), .A4(new_n532), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n628), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n620), .B1(new_n539), .B2(new_n540), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n571), .A2(new_n500), .A3(new_n302), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT90), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR4_X1   g0525(.A1(new_n593), .A2(new_n469), .A3(new_n594), .A4(new_n470), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(new_n629), .A3(KEYINPUT30), .A4(new_n541), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n719), .A2(new_n722), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n664), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n722), .A2(new_n727), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n723), .A2(new_n724), .ZN(new_n733));
  OAI211_X1 g0533(.A(KEYINPUT31), .B(new_n664), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n716), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G330), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n714), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n694), .B1(new_n737), .B2(G1), .ZN(G364));
  AND2_X1   g0538(.A1(new_n207), .A2(G13), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n206), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n687), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n676), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G330), .B2(new_n674), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n210), .A2(new_n284), .ZN(new_n745));
  INV_X1    g0545(.A(G355), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n746), .B1(G116), .B2(new_n210), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n686), .A2(new_n409), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n458), .B2(new_n228), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n251), .A2(new_n458), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n747), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(G1), .B(G13), .C1(new_n207), .C2(G169), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n753), .A2(KEYINPUT93), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(KEYINPUT93), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n742), .B1(new_n752), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n207), .A2(G179), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n445), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n222), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G190), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G159), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT32), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n207), .A2(new_n302), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n445), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n765), .B(new_n770), .C1(G50), .C2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n445), .A2(G179), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n207), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n486), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n771), .A2(new_n766), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n771), .A2(G190), .A3(new_n293), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n284), .B1(new_n778), .B2(new_n220), .C1(new_n258), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n772), .A2(G190), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n777), .B(new_n780), .C1(G68), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT94), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n774), .B(new_n782), .C1(new_n216), .C2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G303), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n615), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT95), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  INV_X1    g0592(.A(G329), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n764), .A2(new_n792), .B1(new_n767), .B2(new_n793), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT96), .Z(new_n795));
  INV_X1    g0595(.A(new_n776), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n566), .ZN(new_n797));
  INV_X1    g0597(.A(new_n779), .ZN(new_n798));
  INV_X1    g0598(.A(new_n778), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n798), .A2(G322), .B1(new_n799), .B2(G311), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT33), .B(G317), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G326), .A2(new_n773), .B1(new_n781), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n795), .A2(new_n797), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n788), .B1(new_n791), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n762), .B1(new_n804), .B2(new_n756), .ZN(new_n805));
  INV_X1    g0605(.A(new_n759), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n674), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n744), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  INV_X1    g0609(.A(G294), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n615), .B1(new_n778), .B2(new_n601), .C1(new_n810), .C2(new_n779), .ZN(new_n811));
  INV_X1    g0611(.A(new_n781), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n812), .A2(new_n792), .B1(new_n486), .B2(new_n776), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n811), .B(new_n813), .C1(G303), .C2(new_n773), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n222), .B2(new_n787), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n764), .A2(new_n216), .B1(new_n767), .B2(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT98), .Z(new_n818));
  AOI22_X1  g0618(.A1(new_n798), .A2(G143), .B1(new_n799), .B2(G159), .ZN(new_n819));
  INV_X1    g0619(.A(new_n773), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n819), .B1(new_n820), .B2(new_n821), .C1(new_n822), .C2(new_n812), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT34), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n764), .A2(new_n214), .ZN(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n409), .B1(new_n827), .B2(new_n767), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n826), .B(new_n828), .C1(G58), .C2(new_n796), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n825), .B(new_n829), .C1(new_n202), .C2(new_n787), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n823), .A2(new_n824), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n815), .A2(new_n818), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n756), .ZN(new_n833));
  INV_X1    g0633(.A(new_n742), .ZN(new_n834));
  INV_X1    g0634(.A(new_n756), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n758), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT97), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n834), .B1(new_n838), .B2(new_n220), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n361), .A2(new_n664), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n366), .A2(new_n363), .B1(new_n365), .B2(new_n665), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(new_n361), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n833), .B(new_n839), .C1(new_n842), .C2(new_n758), .ZN(new_n843));
  INV_X1    g0643(.A(new_n842), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n709), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n367), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n846), .B(new_n665), .C1(new_n644), .C2(new_n656), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(KEYINPUT99), .A3(new_n736), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n849), .B(new_n834), .C1(new_n736), .C2(new_n848), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT99), .B1(new_n848), .B2(new_n736), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n843), .B1(new_n850), .B2(new_n851), .ZN(G384));
  INV_X1    g0652(.A(new_n548), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n230), .A4(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(KEYINPUT100), .B(KEYINPUT36), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n856), .B(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n228), .B(G77), .C1(new_n258), .C2(new_n214), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n206), .B(G13), .C1(new_n859), .C2(new_n247), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n456), .B1(KEYINPUT29), .B2(new_n700), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n711), .B2(new_n713), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n640), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT103), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT39), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT102), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n411), .A2(new_n373), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n370), .B1(new_n868), .B2(new_n412), .ZN(new_n869));
  INV_X1    g0669(.A(new_n662), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n411), .A2(new_n373), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n436), .B1(new_n405), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(KEYINPUT102), .A3(new_n662), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n635), .B2(new_n638), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n431), .A2(new_n873), .A3(new_n433), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n449), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n878), .B2(new_n875), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n439), .A2(new_n443), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n439), .A2(new_n662), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .A4(new_n449), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n876), .A2(KEYINPUT38), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n449), .B1(new_n416), .B2(new_n434), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n416), .A2(new_n870), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n883), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n635), .B2(new_n638), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n866), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n876), .A2(new_n884), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n876), .A2(new_n884), .A3(KEYINPUT38), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n341), .A2(new_n664), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n892), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n636), .A2(new_n662), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n895), .A2(new_n896), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n664), .A2(new_n340), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n902), .B(KEYINPUT101), .Z(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n344), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n341), .A2(new_n903), .A3(new_n343), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n840), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n847), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n900), .B1(new_n901), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n899), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n865), .B(new_n911), .Z(new_n912));
  INV_X1    g0712(.A(KEYINPUT105), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n512), .A2(new_n633), .A3(new_n664), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n731), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n913), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT31), .B1(new_n728), .B2(new_n664), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n716), .A2(KEYINPUT105), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n905), .A2(new_n842), .A3(new_n906), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT38), .B1(new_n876), .B2(new_n884), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n922), .B(new_n924), .C1(new_n885), .C2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n928), .B(new_n923), .C1(new_n917), .C2(new_n921), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n883), .A2(new_n888), .B1(new_n454), .B2(new_n887), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n896), .B1(new_n930), .B2(KEYINPUT38), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n926), .A2(new_n927), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n368), .A2(new_n922), .A3(new_n455), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(G330), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n912), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n206), .B2(new_n739), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n912), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n861), .B1(new_n939), .B2(new_n940), .ZN(G367));
  NOR2_X1   g0741(.A1(new_n665), .A2(new_n492), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n652), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n653), .B2(new_n942), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT106), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n759), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n761), .B1(new_n686), .B2(new_n476), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n748), .A2(new_n240), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n834), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n779), .A2(new_n822), .B1(new_n778), .B2(new_n202), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n615), .B(new_n950), .C1(G137), .C2(new_n768), .ZN(new_n951));
  INV_X1    g0751(.A(new_n787), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(G58), .ZN(new_n953));
  INV_X1    g0753(.A(new_n764), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n773), .A2(G143), .B1(new_n954), .B2(G77), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n776), .A2(new_n214), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(G159), .B2(new_n781), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n951), .A2(new_n953), .A3(new_n955), .A4(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n798), .A2(G303), .B1(new_n768), .B2(G317), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n792), .B2(new_n778), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n409), .B(new_n960), .C1(new_n566), .C2(new_n781), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n952), .A2(KEYINPUT46), .A3(G116), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n820), .A2(new_n816), .B1(new_n222), .B2(new_n776), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(G97), .B2(new_n954), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT46), .B1(new_n952), .B2(G116), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n958), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT47), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n756), .B1(new_n967), .B2(new_n968), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n946), .B(new_n949), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n670), .B(new_n678), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(new_n676), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(new_n714), .A3(new_n736), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT108), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n563), .B1(new_n562), .B2(new_n665), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n642), .A2(new_n664), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n682), .A2(new_n684), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT45), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n682), .A2(new_n684), .ZN(new_n984));
  INV_X1    g0784(.A(new_n979), .ZN(new_n985));
  AND3_X1   g0785(.A1(new_n984), .A2(KEYINPUT44), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT44), .B1(new_n984), .B2(new_n985), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n982), .A2(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(new_n677), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n973), .A2(new_n714), .A3(KEYINPUT108), .A4(new_n736), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n976), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n737), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n687), .B(KEYINPUT41), .Z(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n741), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT43), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n945), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n670), .A2(new_n678), .A3(new_n979), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT42), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n646), .A2(new_n667), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n664), .B1(new_n1000), .B2(new_n641), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n998), .B2(KEYINPUT42), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n997), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n945), .A2(new_n996), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT107), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n670), .A2(new_n676), .A3(new_n979), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1005), .A2(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1007), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n971), .B1(new_n995), .B2(new_n1012), .ZN(G387));
  NAND2_X1  g0813(.A1(new_n973), .A2(new_n741), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n670), .A2(new_n806), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n409), .B1(G326), .B2(new_n768), .ZN(new_n1016));
  INV_X1    g0816(.A(G317), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n779), .A2(new_n1017), .B1(new_n778), .B2(new_n789), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT112), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(KEYINPUT112), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G311), .A2(new_n781), .B1(new_n773), .B2(G322), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n952), .A2(new_n566), .B1(G283), .B2(new_n796), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1016), .B1(new_n601), .B2(new_n764), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1030));
  INV_X1    g0830(.A(G159), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n820), .A2(new_n1031), .B1(new_n346), .B2(new_n776), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n399), .B(new_n1032), .C1(G97), .C2(new_n954), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n798), .A2(G50), .B1(new_n768), .B2(G150), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n214), .B2(new_n778), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n261), .B2(new_n781), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1033), .B(new_n1036), .C1(new_n220), .C2(new_n787), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT111), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n756), .B1(new_n1030), .B2(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n690), .A2(new_n745), .B1(G107), .B2(new_n210), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n237), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n749), .B1(new_n1041), .B2(G45), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n690), .A2(KEYINPUT109), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n690), .A2(KEYINPUT109), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n256), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1040), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1049), .A2(KEYINPUT110), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(KEYINPUT110), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n760), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1039), .B(new_n742), .C1(new_n1050), .C2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n737), .A2(new_n973), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n974), .A2(new_n687), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1014), .B1(new_n1015), .B2(new_n1053), .C1(new_n1054), .C2(new_n1055), .ZN(G393));
  INV_X1    g0856(.A(new_n989), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n688), .B1(new_n1057), .B2(new_n974), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1058), .A2(new_n991), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n245), .A2(new_n749), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n760), .B1(new_n486), .B2(new_n210), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n742), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G317), .A2(new_n773), .B1(new_n798), .B2(G311), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n952), .A2(G283), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n776), .A2(new_n601), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n765), .B(new_n1067), .C1(G303), .C2(new_n781), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n615), .B1(new_n778), .B2(new_n810), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G322), .B2(new_n768), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n820), .A2(new_n822), .B1(new_n1031), .B2(new_n779), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT51), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n764), .A2(new_n216), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n399), .B(new_n1074), .C1(G143), .C2(new_n768), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1073), .B(new_n1075), .C1(new_n214), .C2(new_n787), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n776), .A2(new_n220), .B1(new_n778), .B2(new_n256), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G50), .B2(new_n781), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT113), .Z(new_n1079));
  OAI21_X1  g0879(.A(new_n1071), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1062), .B1(new_n1080), .B2(new_n756), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n979), .B2(new_n806), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n1057), .B2(new_n740), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1059), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(G390));
  XNOR2_X1  g0885(.A(KEYINPUT54), .B(G143), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n781), .A2(G137), .B1(new_n799), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1089), .A2(KEYINPUT116), .B1(G159), .B2(new_n796), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(KEYINPUT116), .B2(new_n1089), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT117), .Z(new_n1092));
  NAND2_X1  g0892(.A1(new_n952), .A2(G150), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT53), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n615), .B1(new_n768), .B2(G125), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n827), .B2(new_n779), .ZN(new_n1096));
  INV_X1    g0896(.A(G128), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n820), .A2(new_n1097), .B1(new_n764), .B2(new_n202), .ZN(new_n1098));
  NOR4_X1   g0898(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n812), .A2(new_n222), .B1(new_n820), .B2(new_n792), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n826), .B(new_n1100), .C1(G77), .C2(new_n796), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n778), .A2(new_n486), .B1(new_n767), .B2(new_n810), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n284), .B(new_n1102), .C1(G116), .C2(new_n798), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(new_n216), .C2(new_n787), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT118), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n756), .B1(new_n1099), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1106), .B(new_n742), .C1(new_n261), .C2(new_n837), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n892), .A2(new_n897), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1107), .B1(new_n1108), .B2(new_n757), .ZN(new_n1109));
  INV_X1    g0909(.A(G330), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n917), .B2(new_n921), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1111), .A2(new_n924), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n907), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n664), .B(new_n367), .C1(new_n704), .C2(new_n705), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n840), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n898), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n892), .A2(new_n897), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n841), .A2(new_n361), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n665), .B(new_n1118), .C1(new_n695), .C2(new_n698), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n908), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n1113), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1121), .A2(new_n1116), .A3(new_n931), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1112), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n840), .B1(new_n706), .B2(new_n846), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1116), .B1(new_n1124), .B2(new_n907), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n889), .A2(new_n890), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n894), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT39), .B1(new_n1127), .B2(new_n896), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n885), .A2(new_n925), .A3(new_n866), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1125), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1121), .A2(new_n1116), .A3(new_n931), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1113), .A2(new_n735), .A3(G330), .A4(new_n842), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1123), .A2(new_n1133), .A3(KEYINPUT115), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT115), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1135), .B(new_n1112), .C1(new_n1117), .C2(new_n1122), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1109), .B1(new_n1137), .B2(new_n741), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n735), .A2(G330), .A3(new_n842), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1111), .A2(new_n924), .B1(new_n1139), .B2(new_n907), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1113), .B1(new_n1111), .B2(new_n842), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1132), .A2(new_n908), .A3(new_n1119), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1140), .A2(new_n1124), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1111), .A2(new_n455), .A3(new_n368), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n863), .A2(new_n1143), .A3(new_n640), .A4(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1134), .A2(new_n1145), .A3(new_n1136), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n687), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1138), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT119), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1138), .B(KEYINPUT119), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(G378));
  INV_X1    g0954(.A(KEYINPUT57), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n863), .A2(new_n640), .A3(new_n1144), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n1137), .B2(new_n1143), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n885), .A2(new_n925), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n914), .A2(new_n916), .A3(new_n913), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT105), .B1(new_n716), .B2(new_n920), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n924), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n927), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n931), .A2(KEYINPUT40), .A3(new_n922), .A4(new_n924), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(G330), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1164), .A2(new_n899), .A3(new_n910), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n911), .A2(new_n932), .A3(G330), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n300), .A2(new_n662), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT55), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n306), .B(new_n1169), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1171));
  XOR2_X1   g0971(.A(new_n1170), .B(new_n1171), .Z(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1167), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1165), .A2(new_n1166), .A3(new_n1172), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1155), .B1(new_n1157), .B2(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1165), .A2(new_n1166), .A3(new_n1172), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1172), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(KEYINPUT57), .C1(new_n1156), .C2(new_n1148), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1177), .A2(new_n1181), .A3(new_n687), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1178), .A2(new_n1179), .A3(new_n740), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n742), .B1(new_n836), .B2(G50), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n812), .A2(new_n486), .B1(new_n346), .B2(new_n778), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(KEYINPUT120), .A2(new_n1185), .B1(new_n952), .B2(G77), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(KEYINPUT120), .B2(new_n1185), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n513), .B1(new_n767), .B2(new_n792), .C1(new_n779), .C2(new_n222), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n956), .A2(new_n409), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n258), .B2(new_n764), .C1(new_n601), .C2(new_n820), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n513), .B1(new_n384), .B2(new_n374), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1191), .A2(KEYINPUT58), .B1(new_n202), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n952), .A2(new_n1087), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT121), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT121), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n779), .A2(new_n1097), .B1(new_n778), .B2(new_n821), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G125), .B2(new_n773), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G150), .A2(new_n796), .B1(new_n781), .B2(G132), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1195), .A2(new_n1196), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n954), .A2(G159), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G33), .B(G41), .C1(new_n768), .C2(G124), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1193), .B1(KEYINPUT58), .B2(new_n1191), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1184), .B1(new_n1206), .B2(new_n756), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1172), .B2(new_n758), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1183), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1182), .A2(new_n1210), .ZN(G375));
  INV_X1    g1011(.A(new_n1143), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1156), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(new_n994), .A3(new_n1145), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n907), .A2(new_n757), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n820), .A2(new_n827), .B1(new_n202), .B2(new_n776), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n781), .B2(new_n1087), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n952), .A2(G159), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n778), .A2(new_n822), .B1(new_n767), .B2(new_n1097), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G137), .B2(new_n798), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n399), .B1(G58), .B2(new_n954), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1217), .A2(new_n1218), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n779), .A2(new_n792), .B1(new_n767), .B2(new_n789), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n284), .B(new_n1223), .C1(G107), .C2(new_n799), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n952), .A2(G97), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n796), .A2(new_n476), .B1(new_n954), .B2(G77), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G116), .A2(new_n781), .B1(new_n773), .B2(G294), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n835), .B1(new_n1222), .B2(new_n1228), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n834), .B(new_n1229), .C1(new_n214), .C2(new_n838), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1143), .A2(new_n741), .B1(new_n1215), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1214), .A2(new_n1231), .ZN(G381));
  OR2_X1    g1032(.A1(G381), .A2(G384), .ZN(new_n1233));
  OR4_X1    g1033(.A1(G396), .A2(G390), .A3(G393), .A4(new_n1233), .ZN(new_n1234));
  OR4_X1    g1034(.A1(G387), .A2(new_n1234), .A3(new_n1149), .A4(G375), .ZN(G407));
  INV_X1    g1035(.A(new_n1149), .ZN(new_n1236));
  INV_X1    g1036(.A(G343), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G407), .B(G213), .C1(G375), .C2(new_n1238), .ZN(G409));
  XNOR2_X1  g1039(.A(G387), .B(new_n1084), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(G393), .B(new_n808), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1240), .B(new_n1241), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1182), .A2(new_n1151), .A3(new_n1152), .A4(new_n1210), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT123), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1183), .B2(new_n1209), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1180), .B(new_n994), .C1(new_n1156), .C2(new_n1148), .ZN(new_n1246));
  OAI211_X1 g1046(.A(KEYINPUT123), .B(new_n1208), .C1(new_n1176), .C2(new_n740), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1236), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1243), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1237), .A2(G213), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1237), .A2(G213), .A3(G2897), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT124), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G384), .A2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(KEYINPUT124), .B(new_n843), .C1(new_n850), .C2(new_n851), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1257), .A2(new_n1231), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT60), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1213), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1156), .A2(new_n1212), .A3(KEYINPUT60), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1260), .A2(new_n687), .A3(new_n1145), .A4(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1256), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1258), .A2(new_n1262), .A3(new_n1256), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1254), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1265), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1267), .A2(new_n1263), .A3(new_n1253), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT61), .B1(new_n1252), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1250), .A2(new_n1251), .A3(new_n1271), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1272), .A2(KEYINPUT125), .A3(KEYINPUT63), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT63), .B1(new_n1272), .B2(KEYINPUT125), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1242), .B(new_n1270), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1275));
  AND4_X1   g1075(.A1(KEYINPUT62), .A2(new_n1250), .A3(new_n1251), .A4(new_n1271), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1243), .A2(new_n1249), .B1(G213), .B2(new_n1237), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT62), .B1(new_n1277), .B2(new_n1271), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1270), .B(KEYINPUT126), .C1(new_n1276), .C2(new_n1278), .ZN(new_n1279));
  XOR2_X1   g1079(.A(new_n1240), .B(new_n1241), .Z(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT62), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1272), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1277), .A2(KEYINPUT62), .A3(new_n1271), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT126), .B1(new_n1285), .B2(new_n1270), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1275), .B1(new_n1281), .B2(new_n1286), .ZN(G405));
  NAND2_X1  g1087(.A1(G375), .A2(new_n1236), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1243), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1271), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1288), .A2(new_n1243), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1290), .A2(KEYINPUT127), .A3(new_n1291), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1280), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1242), .A2(KEYINPUT127), .A3(new_n1290), .A4(new_n1291), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(G402));
endmodule


