

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  XOR2_X1 U322 ( .A(n307), .B(n417), .Z(n534) );
  XNOR2_X1 U323 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U324 ( .A(n407), .B(KEYINPUT47), .ZN(n408) );
  XNOR2_X1 U325 ( .A(n339), .B(n338), .ZN(n343) );
  XNOR2_X1 U326 ( .A(n409), .B(n408), .ZN(n415) );
  NOR2_X1 U327 ( .A1(n534), .A2(n454), .ZN(n568) );
  XNOR2_X1 U328 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U329 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n292) );
  XOR2_X1 U331 ( .A(G190GAT), .B(G134GAT), .Z(n394) );
  XNOR2_X1 U332 ( .A(G127GAT), .B(KEYINPUT85), .ZN(n290) );
  XNOR2_X1 U333 ( .A(n290), .B(KEYINPUT0), .ZN(n444) );
  XNOR2_X1 U334 ( .A(n394), .B(n444), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n302) );
  XOR2_X1 U336 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n294) );
  NAND2_X1 U337 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U339 ( .A(n295), .B(KEYINPUT87), .Z(n300) );
  XOR2_X1 U340 ( .A(G15GAT), .B(G113GAT), .Z(n297) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(G43GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n351) );
  XNOR2_X1 U343 ( .A(G99GAT), .B(G71GAT), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n298), .B(G120GAT), .ZN(n341) );
  XNOR2_X1 U345 ( .A(n351), .B(n341), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n307) );
  XOR2_X1 U348 ( .A(G176GAT), .B(KEYINPUT18), .Z(n304) );
  XNOR2_X1 U349 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n306) );
  XOR2_X1 U351 ( .A(KEYINPUT17), .B(KEYINPUT88), .Z(n305) );
  XOR2_X1 U352 ( .A(n306), .B(n305), .Z(n417) );
  XOR2_X1 U353 ( .A(KEYINPUT21), .B(KEYINPUT94), .Z(n309) );
  XNOR2_X1 U354 ( .A(G218GAT), .B(KEYINPUT93), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U356 ( .A(n310), .B(G211GAT), .Z(n312) );
  XNOR2_X1 U357 ( .A(G197GAT), .B(G204GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n424) );
  XOR2_X1 U359 ( .A(KEYINPUT92), .B(KEYINPUT24), .Z(n314) );
  XNOR2_X1 U360 ( .A(G50GAT), .B(KEYINPUT23), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n424), .B(n315), .ZN(n325) );
  XOR2_X1 U363 ( .A(G155GAT), .B(KEYINPUT3), .Z(n317) );
  XNOR2_X1 U364 ( .A(KEYINPUT95), .B(KEYINPUT2), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n431) );
  XOR2_X1 U366 ( .A(KEYINPUT76), .B(G162GAT), .Z(n399) );
  XOR2_X1 U367 ( .A(n431), .B(n399), .Z(n323) );
  XOR2_X1 U368 ( .A(G141GAT), .B(G22GAT), .Z(n347) );
  XNOR2_X1 U369 ( .A(G106GAT), .B(G78GAT), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n318), .B(G148GAT), .ZN(n340) );
  XOR2_X1 U371 ( .A(n340), .B(KEYINPUT22), .Z(n320) );
  NAND2_X1 U372 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n347), .B(n321), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n475) );
  XOR2_X1 U377 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n365) );
  XOR2_X1 U378 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n327) );
  XNOR2_X1 U379 ( .A(G176GAT), .B(G204GAT), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n345) );
  INV_X1 U381 ( .A(KEYINPUT13), .ZN(n328) );
  NAND2_X1 U382 ( .A1(n328), .A2(KEYINPUT72), .ZN(n331) );
  INV_X1 U383 ( .A(KEYINPUT72), .ZN(n329) );
  NAND2_X1 U384 ( .A1(n329), .A2(KEYINPUT13), .ZN(n330) );
  NAND2_X1 U385 ( .A1(n331), .A2(n330), .ZN(n333) );
  XNOR2_X1 U386 ( .A(G57GAT), .B(G64GAT), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n382) );
  XOR2_X1 U388 ( .A(G85GAT), .B(G92GAT), .Z(n398) );
  XNOR2_X1 U389 ( .A(n382), .B(n398), .ZN(n339) );
  XOR2_X1 U390 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n335) );
  XNOR2_X1 U391 ( .A(KEYINPUT32), .B(KEYINPUT74), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n337) );
  AND2_X1 U393 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  XOR2_X1 U394 ( .A(n341), .B(n340), .Z(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n410) );
  XOR2_X1 U397 ( .A(n410), .B(KEYINPUT41), .Z(n555) );
  XNOR2_X1 U398 ( .A(G1GAT), .B(G8GAT), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n346), .B(KEYINPUT69), .ZN(n383) );
  XOR2_X1 U400 ( .A(n347), .B(n383), .Z(n349) );
  NAND2_X1 U401 ( .A1(G229GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U403 ( .A(n350), .B(KEYINPUT65), .Z(n353) );
  XNOR2_X1 U404 ( .A(n351), .B(KEYINPUT70), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n363) );
  XOR2_X1 U406 ( .A(G50GAT), .B(G29GAT), .Z(n355) );
  XNOR2_X1 U407 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U409 ( .A(n356), .B(KEYINPUT7), .Z(n358) );
  XNOR2_X1 U410 ( .A(G36GAT), .B(KEYINPUT68), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n358), .B(n357), .ZN(n395) );
  XOR2_X1 U412 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n360) );
  XNOR2_X1 U413 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U415 ( .A(n395), .B(n361), .Z(n362) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n574) );
  NAND2_X1 U417 ( .A1(n555), .A2(n574), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n366), .B(KEYINPUT113), .ZN(n386) );
  XOR2_X1 U420 ( .A(G127GAT), .B(G71GAT), .Z(n368) );
  XNOR2_X1 U421 ( .A(G15GAT), .B(G183GAT), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U423 ( .A(G155GAT), .B(G78GAT), .Z(n370) );
  XNOR2_X1 U424 ( .A(G22GAT), .B(G211GAT), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U426 ( .A(n372), .B(n371), .Z(n377) );
  XOR2_X1 U427 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n374) );
  NAND2_X1 U428 ( .A1(G231GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U430 ( .A(KEYINPUT12), .B(n375), .ZN(n376) );
  XNOR2_X1 U431 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U432 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n379) );
  XNOR2_X1 U433 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U435 ( .A(n381), .B(n380), .Z(n385) );
  XNOR2_X1 U436 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U437 ( .A(n385), .B(n384), .Z(n580) );
  INV_X1 U438 ( .A(n580), .ZN(n542) );
  NAND2_X1 U439 ( .A1(n386), .A2(n542), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n387), .B(KEYINPUT115), .ZN(n406) );
  XOR2_X1 U441 ( .A(G106GAT), .B(KEYINPUT78), .Z(n389) );
  NAND2_X1 U442 ( .A1(G232GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U443 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U444 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n391) );
  XNOR2_X1 U445 ( .A(G43GAT), .B(KEYINPUT79), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U447 ( .A(n393), .B(n392), .Z(n397) );
  XNOR2_X1 U448 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U449 ( .A(n397), .B(n396), .ZN(n403) );
  XOR2_X1 U450 ( .A(KEYINPUT77), .B(n398), .Z(n401) );
  XNOR2_X1 U451 ( .A(G218GAT), .B(n399), .ZN(n400) );
  XNOR2_X1 U452 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U453 ( .A(n403), .B(n402), .ZN(n405) );
  XNOR2_X1 U454 ( .A(G99GAT), .B(KEYINPUT11), .ZN(n404) );
  XNOR2_X1 U455 ( .A(n405), .B(n404), .ZN(n567) );
  INV_X1 U456 ( .A(n567), .ZN(n547) );
  NAND2_X1 U457 ( .A1(n406), .A2(n547), .ZN(n409) );
  XNOR2_X1 U458 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n407) );
  XOR2_X1 U459 ( .A(KEYINPUT36), .B(n567), .Z(n496) );
  NOR2_X1 U460 ( .A1(n542), .A2(n496), .ZN(n411) );
  XOR2_X1 U461 ( .A(KEYINPUT45), .B(n411), .Z(n412) );
  NOR2_X1 U462 ( .A1(n410), .A2(n412), .ZN(n413) );
  XOR2_X1 U463 ( .A(KEYINPUT71), .B(n574), .Z(n564) );
  INV_X1 U464 ( .A(n564), .ZN(n536) );
  NAND2_X1 U465 ( .A1(n413), .A2(n536), .ZN(n414) );
  NAND2_X1 U466 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X1 U467 ( .A(n416), .B(KEYINPUT48), .ZN(n551) );
  INV_X1 U468 ( .A(n417), .ZN(n428) );
  XOR2_X1 U469 ( .A(KEYINPUT97), .B(G64GAT), .Z(n419) );
  NAND2_X1 U470 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U472 ( .A(G92GAT), .B(G190GAT), .Z(n421) );
  XNOR2_X1 U473 ( .A(G169GAT), .B(G36GAT), .ZN(n420) );
  XNOR2_X1 U474 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U475 ( .A(n423), .B(n422), .Z(n426) );
  XNOR2_X1 U476 ( .A(G8GAT), .B(n424), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U478 ( .A(n428), .B(n427), .Z(n470) );
  NAND2_X1 U479 ( .A1(n551), .A2(n470), .ZN(n430) );
  XOR2_X1 U480 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n429) );
  XNOR2_X1 U481 ( .A(n430), .B(n429), .ZN(n451) );
  XOR2_X1 U482 ( .A(n431), .B(G134GAT), .Z(n433) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U484 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U485 ( .A(G29GAT), .B(n434), .ZN(n450) );
  XOR2_X1 U486 ( .A(G57GAT), .B(G148GAT), .Z(n436) );
  XNOR2_X1 U487 ( .A(G141GAT), .B(G120GAT), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U489 ( .A(KEYINPUT79), .B(G85GAT), .Z(n438) );
  XNOR2_X1 U490 ( .A(G113GAT), .B(G162GAT), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n448) );
  XOR2_X1 U493 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n442) );
  XNOR2_X1 U494 ( .A(KEYINPUT1), .B(KEYINPUT96), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U496 ( .A(KEYINPUT5), .B(n443), .Z(n446) );
  XNOR2_X1 U497 ( .A(G1GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U500 ( .A(n450), .B(n449), .ZN(n522) );
  NAND2_X1 U501 ( .A1(n451), .A2(n522), .ZN(n452) );
  XNOR2_X1 U502 ( .A(n452), .B(KEYINPUT64), .ZN(n461) );
  NOR2_X1 U503 ( .A1(n475), .A2(n461), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n453), .B(KEYINPUT55), .ZN(n454) );
  NAND2_X1 U505 ( .A1(n568), .A2(n555), .ZN(n458) );
  XOR2_X1 U506 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n456) );
  XOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT56), .Z(n455) );
  INV_X1 U508 ( .A(G218GAT), .ZN(n465) );
  XOR2_X1 U509 ( .A(KEYINPUT99), .B(KEYINPUT26), .Z(n460) );
  NAND2_X1 U510 ( .A1(n475), .A2(n534), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n460), .B(n459), .ZN(n553) );
  NOR2_X1 U512 ( .A1(n461), .A2(n553), .ZN(n581) );
  INV_X1 U513 ( .A(n581), .ZN(n462) );
  NOR2_X1 U514 ( .A1(n496), .A2(n462), .ZN(n463) );
  XNOR2_X1 U515 ( .A(KEYINPUT62), .B(n463), .ZN(n464) );
  XNOR2_X1 U516 ( .A(n465), .B(n464), .ZN(G1355GAT) );
  XOR2_X1 U517 ( .A(KEYINPUT34), .B(KEYINPUT104), .Z(n467) );
  XNOR2_X1 U518 ( .A(G1GAT), .B(KEYINPUT103), .ZN(n466) );
  XNOR2_X1 U519 ( .A(n467), .B(n466), .ZN(n487) );
  NOR2_X1 U520 ( .A1(n536), .A2(n410), .ZN(n499) );
  XOR2_X1 U521 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n469) );
  NAND2_X1 U522 ( .A1(n547), .A2(n580), .ZN(n468) );
  XNOR2_X1 U523 ( .A(n469), .B(n468), .ZN(n485) );
  INV_X1 U524 ( .A(n470), .ZN(n524) );
  XNOR2_X1 U525 ( .A(KEYINPUT27), .B(n524), .ZN(n478) );
  NOR2_X1 U526 ( .A1(n522), .A2(n478), .ZN(n550) );
  XOR2_X1 U527 ( .A(n475), .B(KEYINPUT28), .Z(n530) );
  NAND2_X1 U528 ( .A1(n550), .A2(n530), .ZN(n533) );
  XNOR2_X1 U529 ( .A(KEYINPUT91), .B(n534), .ZN(n471) );
  NOR2_X1 U530 ( .A1(n533), .A2(n471), .ZN(n472) );
  XOR2_X1 U531 ( .A(KEYINPUT98), .B(n472), .Z(n484) );
  XNOR2_X1 U532 ( .A(KEYINPUT100), .B(KEYINPUT25), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n473), .B(KEYINPUT101), .ZN(n477) );
  NOR2_X1 U534 ( .A1(n524), .A2(n534), .ZN(n474) );
  NOR2_X1 U535 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n480) );
  NOR2_X1 U537 ( .A1(n478), .A2(n553), .ZN(n479) );
  NOR2_X1 U538 ( .A1(n480), .A2(n479), .ZN(n481) );
  XOR2_X1 U539 ( .A(KEYINPUT102), .B(n481), .Z(n482) );
  NAND2_X1 U540 ( .A1(n522), .A2(n482), .ZN(n483) );
  NAND2_X1 U541 ( .A1(n484), .A2(n483), .ZN(n494) );
  AND2_X1 U542 ( .A1(n485), .A2(n494), .ZN(n510) );
  NAND2_X1 U543 ( .A1(n499), .A2(n510), .ZN(n491) );
  NOR2_X1 U544 ( .A1(n522), .A2(n491), .ZN(n486) );
  XOR2_X1 U545 ( .A(n487), .B(n486), .Z(G1324GAT) );
  NOR2_X1 U546 ( .A1(n524), .A2(n491), .ZN(n488) );
  XOR2_X1 U547 ( .A(G8GAT), .B(n488), .Z(G1325GAT) );
  NOR2_X1 U548 ( .A1(n534), .A2(n491), .ZN(n490) );
  XNOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NOR2_X1 U551 ( .A1(n530), .A2(n491), .ZN(n493) );
  XNOR2_X1 U552 ( .A(G22GAT), .B(KEYINPUT105), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1327GAT) );
  NAND2_X1 U554 ( .A1(n542), .A2(n494), .ZN(n495) );
  NOR2_X1 U555 ( .A1(n496), .A2(n495), .ZN(n498) );
  XNOR2_X1 U556 ( .A(KEYINPUT107), .B(KEYINPUT37), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(n521) );
  NAND2_X1 U558 ( .A1(n499), .A2(n521), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n500), .B(KEYINPUT108), .ZN(n501) );
  XNOR2_X1 U560 ( .A(KEYINPUT38), .B(n501), .ZN(n508) );
  NOR2_X1 U561 ( .A1(n522), .A2(n508), .ZN(n503) );
  XNOR2_X1 U562 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(n504), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n524), .A2(n508), .ZN(n505) );
  XOR2_X1 U566 ( .A(G36GAT), .B(n505), .Z(G1329GAT) );
  NOR2_X1 U567 ( .A1(n534), .A2(n508), .ZN(n506) );
  XOR2_X1 U568 ( .A(KEYINPUT40), .B(n506), .Z(n507) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NOR2_X1 U570 ( .A1(n530), .A2(n508), .ZN(n509) );
  XOR2_X1 U571 ( .A(G50GAT), .B(n509), .Z(G1331GAT) );
  INV_X1 U572 ( .A(n555), .ZN(n539) );
  NOR2_X1 U573 ( .A1(n539), .A2(n574), .ZN(n520) );
  NAND2_X1 U574 ( .A1(n520), .A2(n510), .ZN(n516) );
  NOR2_X1 U575 ( .A1(n522), .A2(n516), .ZN(n511) );
  XOR2_X1 U576 ( .A(G57GAT), .B(n511), .Z(n512) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U578 ( .A1(n524), .A2(n516), .ZN(n513) );
  XOR2_X1 U579 ( .A(G64GAT), .B(n513), .Z(G1333GAT) );
  NOR2_X1 U580 ( .A1(n534), .A2(n516), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1334GAT) );
  NOR2_X1 U583 ( .A1(n530), .A2(n516), .ZN(n518) );
  XNOR2_X1 U584 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n529) );
  NOR2_X1 U588 ( .A1(n522), .A2(n529), .ZN(n523) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n529), .ZN(n525) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U592 ( .A1(n534), .A2(n529), .ZN(n526) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n528) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(KEYINPUT112), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(n532) );
  NOR2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U598 ( .A(n532), .B(n531), .Z(G1339GAT) );
  NOR2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n551), .A2(n535), .ZN(n546) );
  NOR2_X1 U601 ( .A1(n536), .A2(n546), .ZN(n537) );
  XOR2_X1 U602 ( .A(KEYINPUT118), .B(n537), .Z(n538) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  NOR2_X1 U604 ( .A1(n539), .A2(n546), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NOR2_X1 U607 ( .A1(n542), .A2(n546), .ZN(n544) );
  XNOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT119), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  NOR2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n549) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n574), .A2(n561), .ZN(n554) );
  XNOR2_X1 U617 ( .A(n554), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n559) );
  XOR2_X1 U619 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U620 ( .A1(n561), .A2(n555), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n580), .A2(n561), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U625 ( .A(G162GAT), .B(KEYINPUT121), .Z(n563) );
  NAND2_X1 U626 ( .A1(n561), .A2(n567), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n568), .A2(n564), .ZN(n565) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n580), .A2(n568), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n570), .B(n569), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(n573), .Z(n576) );
  NAND2_X1 U639 ( .A1(n581), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U642 ( .A1(n581), .A2(n410), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(n579), .ZN(G1353GAT) );
  XOR2_X1 U645 ( .A(G211GAT), .B(KEYINPUT127), .Z(n583) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1354GAT) );
endmodule

