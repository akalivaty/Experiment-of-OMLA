//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1195,
    new_n1196, new_n1197, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT64), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n209), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n214), .A2(new_n225), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT65), .B(G50), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  AOI21_X1  g0048(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n251));
  NOR3_X1   g0051(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G45), .ZN(new_n254));
  AOI21_X1  g0054(.A(G1), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G226), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n249), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G222), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n259), .B1(new_n260), .B2(new_n258), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  AOI211_X1 g0064(.A(new_n252), .B(new_n257), .C1(new_n264), .C2(new_n249), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT66), .B1(new_n265), .B2(G169), .ZN(new_n266));
  INV_X1    g0066(.A(G179), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT8), .B(G58), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n209), .A2(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G150), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n270), .A2(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(G20), .B2(new_n203), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n228), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(new_n228), .A3(new_n277), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n208), .A2(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G50), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n282), .A2(new_n284), .B1(G50), .B2(new_n281), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT66), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n287), .B1(new_n268), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n269), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n286), .A2(KEYINPUT9), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT70), .ZN(new_n292));
  INV_X1    g0092(.A(new_n265), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n293), .A2(G200), .B1(KEYINPUT9), .B2(new_n286), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n292), .B(new_n294), .C1(new_n295), .C2(new_n293), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT71), .B1(new_n265), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(new_n299), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n290), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n258), .A2(G232), .A3(G1698), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G97), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT72), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT72), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G33), .A3(G97), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n303), .B(new_n308), .C1(new_n262), .C2(new_n256), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n249), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT13), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n249), .A2(new_n255), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n252), .B1(G238), .B2(new_n312), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n311), .B1(new_n310), .B2(new_n313), .ZN(new_n315));
  OAI21_X1  g0115(.A(G200), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n310), .A2(new_n313), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT13), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(G190), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n281), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n216), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT12), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n273), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n260), .B2(new_n271), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(KEYINPUT11), .A3(new_n278), .ZN(new_n326));
  INV_X1    g0126(.A(new_n282), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(G68), .A3(new_n283), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n323), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT11), .B1(new_n325), .B2(new_n278), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n316), .A2(new_n320), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n314), .A2(new_n315), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT14), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(G169), .C1(new_n314), .C2(new_n315), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT73), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n334), .B2(G179), .ZN(new_n340));
  NOR4_X1   g0140(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT73), .A4(new_n267), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n336), .B(new_n338), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n331), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n333), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n283), .A2(G77), .ZN(new_n345));
  OR3_X1    g0145(.A1(new_n282), .A2(KEYINPUT68), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT68), .B1(new_n282), .B2(new_n345), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n321), .A2(new_n260), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n270), .A2(new_n274), .B1(new_n209), .B2(new_n260), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n271), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n278), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n348), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n249), .A2(new_n250), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n255), .ZN(new_n356));
  INV_X1    g0156(.A(new_n249), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(G244), .A3(new_n251), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT67), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n258), .A2(G232), .A3(new_n261), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n258), .A2(G238), .A3(G1698), .ZN(new_n363));
  INV_X1    g0163(.A(G107), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n362), .B(new_n363), .C1(new_n364), .C2(new_n258), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n249), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT67), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n361), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n354), .B1(new_n368), .B2(G200), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT69), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n370), .ZN(new_n372));
  INV_X1    g0172(.A(new_n368), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G190), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n368), .A2(new_n335), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n376), .B(new_n354), .C1(G179), .C2(new_n368), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n302), .A2(new_n344), .A3(new_n375), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT16), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n258), .B2(G20), .ZN(new_n381));
  INV_X1    g0181(.A(G33), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT3), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT3), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G33), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n216), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G58), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(new_n216), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n390), .B2(new_n201), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n273), .A2(G159), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n379), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n381), .A2(new_n387), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n393), .B1(new_n396), .B2(G68), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n279), .B1(new_n397), .B2(KEYINPUT16), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT74), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n399), .B(new_n379), .C1(new_n388), .C2(new_n393), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n395), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n270), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n283), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n403), .A2(new_n282), .B1(new_n281), .B2(new_n402), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n258), .A2(G226), .A3(G1698), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n258), .A2(G223), .A3(new_n261), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n249), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n252), .B1(G232), .B2(new_n312), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n411), .A2(new_n412), .A3(G179), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n335), .B1(new_n411), .B2(new_n412), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n406), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT18), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n415), .B1(new_n401), .B2(new_n405), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n411), .A2(new_n412), .A3(new_n295), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n312), .A2(G232), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n356), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n249), .B2(new_n410), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n422), .B1(new_n425), .B2(G200), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n401), .A2(new_n426), .A3(new_n405), .ZN(new_n427));
  NOR2_X1   g0227(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XOR2_X1   g0229(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n430));
  NAND4_X1  g0230(.A1(new_n401), .A2(new_n426), .A3(new_n405), .A4(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n418), .A2(new_n421), .A3(new_n429), .A4(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n378), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n217), .A2(new_n261), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n258), .B(new_n434), .C1(G244), .C2(new_n261), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G116), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n357), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n254), .A2(G1), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n250), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n219), .B1(new_n254), .B2(G1), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n357), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n335), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT78), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n437), .A2(new_n441), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n267), .ZN(new_n446));
  NOR4_X1   g0246(.A1(new_n437), .A2(new_n441), .A3(KEYINPUT78), .A4(G179), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n386), .A2(G20), .A3(new_n216), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT19), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT76), .B(G97), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n271), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT80), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT80), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n454), .B(new_n450), .C1(new_n451), .C2(new_n271), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n449), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n209), .B1(new_n308), .B2(new_n450), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n451), .A2(new_n218), .A3(new_n364), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT79), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT79), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(new_n461), .A3(new_n458), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n456), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n278), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n351), .A2(new_n321), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n282), .B1(new_n208), .B2(G33), .ZN(new_n466));
  INV_X1    g0266(.A(new_n351), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n448), .B1(new_n469), .B2(KEYINPUT81), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n463), .A2(new_n278), .B1(new_n321), .B2(new_n351), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT81), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n472), .A3(new_n468), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n442), .A2(G200), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n466), .A2(G87), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n464), .A2(new_n474), .A3(new_n465), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n445), .A2(G190), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n470), .A2(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n258), .A2(new_n209), .A3(G87), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT22), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT22), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n258), .A2(new_n482), .A3(new_n209), .A4(G87), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT24), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n436), .A2(G20), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT23), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(new_n209), .B2(G107), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n364), .A2(KEYINPUT23), .A3(G20), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n484), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n485), .B1(new_n484), .B2(new_n490), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n278), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT25), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n281), .B2(G107), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n321), .A2(KEYINPUT25), .A3(new_n364), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n466), .A2(G107), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n383), .A2(new_n385), .A3(G257), .A4(G1698), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n383), .A2(new_n385), .A3(G250), .A4(new_n261), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G294), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT85), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT85), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n499), .A2(new_n500), .A3(new_n504), .A4(new_n501), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n249), .A3(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n208), .B(G45), .C1(new_n253), .C2(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT77), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n507), .B2(KEYINPUT77), .ZN(new_n511));
  OAI211_X1 g0311(.A(G264), .B(new_n357), .C1(new_n509), .C2(new_n511), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n507), .A2(KEYINPUT77), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n513), .A2(new_n355), .A3(new_n508), .A4(new_n510), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n506), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n515), .A2(G179), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n335), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n498), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G283), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n209), .B(new_n520), .C1(new_n451), .C2(G33), .ZN(new_n521));
  INV_X1    g0321(.A(G116), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n277), .A2(new_n228), .B1(G20), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT20), .ZN(new_n525));
  OR2_X1    g0325(.A1(new_n525), .A2(KEYINPUT84), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(KEYINPUT84), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT83), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n281), .B2(G116), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n321), .A2(KEYINPUT83), .A3(new_n522), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n466), .A2(G116), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n521), .A2(KEYINPUT84), .A3(new_n525), .A4(new_n523), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G169), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n258), .A2(G264), .A3(G1698), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT82), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n258), .A2(KEYINPUT82), .A3(G264), .A4(G1698), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n258), .A2(G257), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(new_n261), .B1(G303), .B2(new_n386), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n357), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G270), .B(new_n357), .C1(new_n509), .C2(new_n511), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n514), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n519), .B1(new_n535), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n540), .A2(new_n542), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n249), .ZN(new_n549));
  INV_X1    g0349(.A(new_n545), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n551), .A2(KEYINPUT21), .A3(G169), .A4(new_n534), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n546), .A2(G179), .A3(new_n534), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n547), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n518), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G97), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n364), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n205), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n364), .A2(KEYINPUT6), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n558), .A2(KEYINPUT6), .B1(new_n451), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(G20), .B1(G77), .B2(new_n273), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n396), .A2(G107), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n279), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n281), .A2(G97), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n466), .B2(G97), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT4), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n383), .A2(new_n385), .A3(G244), .A4(new_n261), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n568), .B(new_n520), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n570), .A2(new_n569), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n249), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G257), .B(new_n357), .C1(new_n509), .C2(new_n511), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n573), .A2(new_n267), .A3(new_n514), .A4(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n514), .A3(new_n574), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n335), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n567), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n515), .A2(G200), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n506), .A2(new_n512), .A3(G190), .A4(new_n514), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n493), .A2(new_n579), .A3(new_n497), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(G200), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n573), .A2(G190), .A3(new_n514), .A4(new_n574), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n582), .A2(new_n564), .A3(new_n566), .A4(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n534), .ZN(new_n585));
  OAI21_X1  g0385(.A(G200), .B1(new_n543), .B2(new_n545), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n585), .B(new_n586), .C1(new_n551), .C2(new_n295), .ZN(new_n587));
  AND4_X1   g0387(.A1(new_n578), .A2(new_n581), .A3(new_n584), .A4(new_n587), .ZN(new_n588));
  AND4_X1   g0388(.A1(new_n433), .A2(new_n479), .A3(new_n555), .A4(new_n588), .ZN(G372));
  INV_X1    g0389(.A(new_n290), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n300), .A2(new_n301), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n419), .B(KEYINPUT18), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n342), .A2(new_n343), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n333), .B2(new_n377), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n429), .A2(new_n431), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n594), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n590), .B1(new_n592), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n433), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n470), .A2(new_n473), .ZN(new_n603));
  INV_X1    g0403(.A(new_n578), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n477), .A2(new_n478), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .A4(KEYINPUT26), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT87), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT86), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n476), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n471), .A2(KEYINPUT86), .A3(new_n474), .A4(new_n475), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n478), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n445), .A2(G169), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n267), .B2(new_n445), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n469), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n604), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT26), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n479), .A2(KEYINPUT87), .A3(KEYINPUT26), .A4(new_n604), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n608), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n578), .A2(new_n581), .A3(new_n584), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n555), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n622), .A2(new_n612), .B1(new_n469), .B2(new_n614), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n601), .B1(new_n602), .B2(new_n625), .ZN(G369));
  NAND3_X1  g0426(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n627), .A2(KEYINPUT27), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(KEYINPUT27), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(G213), .ZN(new_n630));
  INV_X1    g0430(.A(G343), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n585), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n554), .B(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n635), .A2(new_n587), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G330), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n518), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(new_n632), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n498), .A2(new_n632), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n518), .B1(new_n581), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n640), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n554), .A3(new_n633), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(G399));
  INV_X1    g0447(.A(new_n212), .ZN(new_n648));
  OR3_X1    g0448(.A1(new_n648), .A2(KEYINPUT88), .A3(G41), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT88), .B1(new_n648), .B2(G41), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n458), .A2(G116), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G1), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n227), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(new_n651), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT89), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT28), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n632), .B1(new_n620), .B2(new_n623), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT29), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n603), .A2(new_n604), .A3(new_n605), .A4(new_n617), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n578), .A2(new_n584), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n662), .B(new_n581), .C1(new_n554), .C2(new_n518), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n612), .A2(new_n615), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n615), .B(new_n661), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n616), .A2(KEYINPUT26), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n633), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT29), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n660), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n479), .A2(new_n555), .A3(new_n588), .A4(new_n633), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n445), .A2(G179), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n551), .A2(new_n515), .A3(new_n576), .A4(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n549), .A2(G179), .A3(new_n550), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n573), .A2(new_n445), .A3(new_n514), .A4(new_n574), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n506), .A2(new_n512), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n673), .B1(new_n677), .B2(KEYINPUT30), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  NOR4_X1   g0479(.A1(new_n674), .A2(new_n675), .A3(new_n679), .A4(new_n676), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n632), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT31), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g0483(.A(KEYINPUT31), .B(new_n632), .C1(new_n678), .C2(new_n680), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n671), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n670), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n657), .B1(new_n689), .B2(G1), .ZN(G364));
  INV_X1    g0490(.A(new_n651), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n209), .A2(G13), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n208), .B1(new_n692), .B2(G45), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n638), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n636), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(G13), .A2(G33), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT90), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n209), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT91), .Z(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(G1), .B(G13), .C1(new_n209), .C2(G169), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT92), .Z(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n648), .A2(new_n258), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n654), .B2(G45), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n244), .B2(G45), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n212), .A2(new_n258), .ZN(new_n712));
  INV_X1    g0512(.A(G355), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n712), .A2(new_n713), .B1(G116), .B2(new_n212), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n708), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n209), .A2(G179), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(G190), .A3(G200), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n218), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n209), .A2(new_n267), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G200), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n295), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G190), .A2(G200), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G159), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n722), .A2(new_n202), .B1(new_n726), .B2(KEYINPUT32), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n720), .A2(G190), .ZN(new_n728));
  AOI211_X1 g0528(.A(new_n718), .B(new_n727), .C1(G68), .C2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n716), .A2(new_n295), .A3(G200), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT93), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G107), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n719), .A2(G190), .A3(new_n297), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n258), .B1(new_n737), .B2(new_n389), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n719), .A2(new_n723), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n738), .B1(G77), .B2(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n209), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n726), .A2(KEYINPUT32), .B1(new_n744), .B2(G97), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n729), .A2(new_n736), .A3(new_n741), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n735), .A2(G283), .ZN(new_n747));
  INV_X1    g0547(.A(G322), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n737), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G311), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n386), .B1(new_n739), .B2(new_n750), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n749), .B(new_n751), .C1(G329), .C2(new_n725), .ZN(new_n752));
  XNOR2_X1  g0552(.A(KEYINPUT33), .B(G317), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G294), .A2(new_n744), .B1(new_n728), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n717), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n721), .A2(G326), .B1(new_n755), .B2(G303), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n747), .A2(new_n752), .A3(new_n754), .A4(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n746), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n715), .B(new_n695), .C1(new_n758), .C2(new_n706), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT94), .Z(new_n760));
  OR2_X1    g0560(.A1(new_n636), .A2(new_n703), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n696), .A2(new_n698), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(G396));
  NAND2_X1  g0563(.A1(new_n354), .A2(new_n632), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n374), .B1(new_n369), .B2(new_n370), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n369), .A2(new_n370), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n377), .B(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT96), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n375), .A2(KEYINPUT96), .A3(new_n377), .A4(new_n764), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n632), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n624), .A2(new_n771), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n377), .A2(new_n633), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n769), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n772), .B1(new_n658), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n695), .B1(new_n775), .B2(new_n687), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n687), .B2(new_n775), .ZN(new_n777));
  INV_X1    g0577(.A(new_n695), .ZN(new_n778));
  INV_X1    g0578(.A(new_n737), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n779), .A2(G143), .B1(new_n740), .B2(G159), .ZN(new_n780));
  INV_X1    g0580(.A(new_n728), .ZN(new_n781));
  INV_X1    g0581(.A(G137), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n780), .B1(new_n781), .B2(new_n272), .C1(new_n782), .C2(new_n722), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT34), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n735), .A2(G68), .ZN(new_n787));
  INV_X1    g0587(.A(G132), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n258), .B1(new_n724), .B2(new_n788), .C1(new_n743), .C2(new_n389), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(G50), .B2(new_n755), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n785), .A2(new_n786), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G294), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n737), .A2(new_n792), .B1(new_n724), .B2(new_n750), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n258), .B(new_n793), .C1(G116), .C2(new_n740), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n735), .A2(G87), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n744), .A2(G97), .B1(new_n755), .B2(G107), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G283), .A2(new_n728), .B1(new_n721), .B2(G303), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n706), .B1(new_n791), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n699), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n706), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT95), .Z(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n778), .B(new_n799), .C1(new_n260), .C2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n774), .B2(new_n700), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n777), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G384));
  OR2_X1    g0607(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n808), .A2(G116), .A3(new_n229), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(KEYINPUT97), .B(KEYINPUT36), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n227), .B(G77), .C1(new_n389), .C2(new_n216), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n202), .A2(G68), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n208), .B(G13), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n331), .A2(new_n633), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n595), .A2(new_n332), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT98), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n334), .A2(new_n339), .A3(G179), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n318), .A2(G179), .A3(new_n319), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(KEYINPUT73), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n824), .A2(new_n336), .A3(new_n338), .A4(new_n332), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n820), .B1(new_n825), .B2(new_n817), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n819), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n825), .A2(new_n820), .A3(new_n817), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n377), .A2(new_n632), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n829), .B1(new_n772), .B2(new_n831), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n401), .A2(new_n405), .A3(new_n426), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n419), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  INV_X1    g0635(.A(new_n630), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT100), .B1(new_n406), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT100), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n838), .B(new_n630), .C1(new_n401), .C2(new_n405), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n834), .B(new_n835), .C1(new_n837), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n398), .A2(new_n394), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n405), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT99), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(new_n843), .A3(new_n836), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n404), .B1(new_n398), .B2(new_n394), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT99), .B1(new_n845), .B2(new_n630), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n427), .B1(new_n415), .B2(new_n845), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT37), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n840), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n432), .A2(new_n847), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n850), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n832), .A2(new_n855), .B1(new_n594), .B2(new_n630), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT39), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n597), .A2(KEYINPUT101), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT101), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n429), .A2(new_n859), .A3(new_n431), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n858), .A2(new_n593), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n837), .A2(new_n839), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n417), .A2(new_n427), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT37), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n861), .A2(new_n862), .B1(new_n864), .B2(new_n840), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n857), .B(new_n854), .C1(new_n865), .C2(KEYINPUT38), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n850), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT39), .B1(new_n867), .B2(new_n852), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT102), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n595), .A2(new_n632), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n861), .A2(new_n862), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n864), .A2(new_n840), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n875), .A2(KEYINPUT102), .A3(new_n857), .A4(new_n854), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n870), .A2(new_n871), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n856), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n600), .B1(new_n669), .B2(new_n433), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n878), .B(new_n879), .Z(new_n880));
  OAI21_X1  g0680(.A(new_n854), .B1(new_n865), .B2(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n685), .A2(KEYINPUT103), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT103), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n671), .A2(new_n683), .A3(new_n883), .A4(new_n684), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n827), .A2(new_n774), .A3(new_n828), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n881), .A2(new_n882), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n828), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n819), .B2(new_n826), .ZN(new_n888));
  AND4_X1   g0688(.A1(new_n774), .A2(new_n882), .A3(new_n888), .A4(new_n884), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT40), .B1(new_n853), .B2(new_n854), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n886), .A2(KEYINPUT40), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n882), .A2(new_n884), .ZN(new_n892));
  OR3_X1    g0692(.A1(new_n891), .A2(new_n602), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n891), .B1(new_n602), .B2(new_n892), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(G330), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n880), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n208), .B2(new_n692), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n880), .A2(new_n895), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n816), .B1(new_n897), .B2(new_n898), .ZN(G367));
  AOI21_X1  g0699(.A(new_n633), .B1(new_n471), .B2(new_n475), .ZN(new_n900));
  MUX2_X1   g0700(.A(new_n664), .B(new_n615), .S(new_n900), .Z(new_n901));
  AND2_X1   g0701(.A1(new_n901), .A2(new_n704), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n709), .A2(new_n239), .B1(new_n648), .B2(new_n467), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n778), .B1(new_n708), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n743), .A2(new_n216), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(G58), .B2(new_n755), .ZN(new_n906));
  INV_X1    g0706(.A(G143), .ZN(new_n907));
  INV_X1    g0707(.A(G159), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n906), .B1(new_n907), .B2(new_n722), .C1(new_n908), .C2(new_n781), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n734), .A2(new_n260), .ZN(new_n910));
  XOR2_X1   g0710(.A(KEYINPUT106), .B(G137), .Z(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n725), .A2(new_n912), .B1(new_n740), .B2(G50), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n913), .B(new_n258), .C1(new_n272), .C2(new_n737), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n909), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n792), .A2(new_n781), .B1(new_n722), .B2(new_n750), .ZN(new_n916));
  AOI22_X1  g0716(.A1(G283), .A2(new_n740), .B1(new_n725), .B2(G317), .ZN(new_n917));
  INV_X1    g0717(.A(G303), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n917), .B(new_n386), .C1(new_n918), .C2(new_n737), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n916), .B(new_n919), .C1(G107), .C2(new_n744), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT105), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n717), .B2(new_n522), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n922), .A2(KEYINPUT46), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n922), .A2(KEYINPUT46), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n451), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n923), .B(new_n925), .C1(new_n926), .C2(new_n735), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n915), .B1(new_n920), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT47), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n707), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n928), .A2(KEYINPUT47), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n904), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n902), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n646), .A2(new_n645), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n567), .A2(new_n632), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n662), .A2(new_n935), .B1(new_n604), .B2(new_n632), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT104), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT44), .Z(new_n939));
  NOR2_X1   g0739(.A1(new_n934), .A2(new_n937), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT45), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n644), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n939), .A2(new_n644), .A3(new_n941), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n554), .A2(new_n633), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n643), .B(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(new_n638), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n688), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n651), .B(KEYINPUT41), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n693), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n937), .A2(new_n646), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n578), .B1(new_n937), .B2(new_n639), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n953), .A2(KEYINPUT42), .B1(new_n954), .B2(new_n633), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(KEYINPUT42), .B2(new_n953), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT43), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n901), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n901), .A2(new_n957), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n959), .B(new_n960), .Z(new_n961));
  NOR2_X1   g0761(.A1(new_n644), .A2(new_n937), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n933), .B1(new_n952), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(G387));
  NOR2_X1   g0765(.A1(new_n688), .A2(new_n948), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(new_n651), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n689), .B2(new_n949), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n709), .B1(new_n236), .B2(new_n254), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n652), .B2(new_n712), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n270), .A2(G50), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT50), .ZN(new_n972));
  AOI21_X1  g0772(.A(G45), .B1(G68), .B2(G77), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n652), .A3(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n970), .A2(new_n974), .B1(new_n364), .B2(new_n648), .ZN(new_n975));
  INV_X1    g0775(.A(new_n708), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n695), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n258), .B1(new_n724), .B2(new_n272), .C1(new_n216), .C2(new_n739), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n722), .A2(new_n908), .B1(new_n717), .B2(new_n260), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n402), .C2(new_n728), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n744), .A2(new_n467), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n202), .B2(new_n737), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT108), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n980), .B(new_n983), .C1(new_n556), .C2(new_n734), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n779), .A2(G317), .B1(new_n740), .B2(G303), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n781), .B2(new_n750), .C1(new_n748), .C2(new_n722), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT48), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(G283), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n988), .B1(new_n989), .B2(new_n743), .C1(new_n792), .C2(new_n717), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n986), .A2(new_n987), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT49), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n735), .A2(G116), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n258), .B1(new_n725), .B2(G326), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n992), .A2(KEYINPUT49), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n984), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n977), .B1(new_n998), .B2(new_n707), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n643), .B2(new_n703), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT109), .Z(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT107), .B1(new_n949), .B2(new_n694), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n949), .A2(KEYINPUT107), .A3(new_n694), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n968), .B(new_n1001), .C1(new_n1002), .C2(new_n1003), .ZN(G393));
  AOI22_X1  g0804(.A1(new_n709), .A2(new_n247), .B1(new_n648), .B2(new_n926), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n778), .B1(new_n708), .B2(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G317), .A2(new_n721), .B1(new_n779), .B2(G311), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT52), .Z(new_n1008));
  OAI21_X1  g0808(.A(new_n386), .B1(new_n739), .B2(new_n792), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G322), .B2(new_n725), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n781), .A2(new_n918), .B1(new_n717), .B2(new_n989), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G116), .B2(new_n744), .ZN(new_n1012));
  AND4_X1   g0812(.A1(new_n736), .A2(new_n1008), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n258), .B1(new_n724), .B2(new_n907), .C1(new_n216), .C2(new_n717), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n744), .A2(G77), .B1(new_n740), .B2(new_n402), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n202), .B2(new_n781), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT113), .Z(new_n1017));
  AOI211_X1 g0817(.A(new_n1014), .B(new_n1017), .C1(G87), .C2(new_n735), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n722), .A2(new_n272), .B1(new_n908), .B2(new_n737), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT112), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT51), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1013), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1006), .B1(new_n1022), .B2(new_n706), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n937), .B2(new_n704), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT110), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n943), .A2(new_n1025), .A3(new_n944), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n944), .A2(new_n1025), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n942), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT111), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n693), .B1(new_n1029), .B2(KEYINPUT111), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1024), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n651), .B1(new_n945), .B2(new_n966), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n966), .B2(new_n1029), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1034), .ZN(G390));
  INV_X1    g0835(.A(KEYINPUT115), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n885), .A2(G330), .A3(new_n882), .A4(new_n884), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n769), .A2(new_n770), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n633), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n620), .B2(new_n623), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n888), .B1(new_n1041), .B2(new_n830), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n871), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n870), .A2(new_n876), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n871), .B(KEYINPUT114), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n881), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n771), .B1(new_n665), .B2(new_n666), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n829), .B1(new_n1047), .B2(new_n831), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1036), .B(new_n1038), .C1(new_n1044), .C2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n870), .A2(new_n876), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(KEYINPUT115), .B1(new_n1053), .B2(new_n1037), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n686), .A2(new_n774), .A3(new_n888), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1044), .A2(new_n1049), .A3(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1050), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1051), .A2(new_n701), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n802), .A2(new_n402), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n737), .A2(new_n522), .B1(new_n739), .B2(new_n451), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n258), .B(new_n1061), .C1(G294), .C2(new_n725), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n718), .B1(G77), .B2(new_n744), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G107), .A2(new_n728), .B1(new_n721), .B2(G283), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1062), .A2(new_n787), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n779), .A2(G132), .B1(new_n725), .B2(G125), .ZN(new_n1066));
  OR3_X1    g0866(.A1(new_n717), .A2(KEYINPUT53), .A3(new_n272), .ZN(new_n1067));
  OAI21_X1  g0867(.A(KEYINPUT53), .B1(new_n717), .B2(new_n272), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(KEYINPUT54), .B(G143), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n386), .B1(new_n740), .B2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G159), .A2(new_n744), .B1(new_n728), .B2(new_n912), .ZN(new_n1073));
  INV_X1    g0873(.A(G128), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1073), .B1(new_n1074), .B2(new_n722), .C1(new_n202), .C2(new_n734), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1065), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n778), .B(new_n1060), .C1(new_n707), .C2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1058), .A2(new_n694), .B1(new_n1059), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT118), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n888), .B1(new_n686), .B2(new_n774), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1038), .A2(new_n1080), .B1(new_n1041), .B2(new_n830), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1047), .A2(new_n831), .ZN(new_n1082));
  INV_X1    g0882(.A(G330), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n774), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n892), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1082), .B(new_n1055), .C1(new_n1085), .C2(new_n888), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n433), .A2(G330), .A3(new_n882), .A4(new_n884), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(new_n879), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(KEYINPUT117), .B1(new_n1058), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1049), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1092), .A2(new_n1093), .A3(new_n1055), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1038), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n1095), .A3(KEYINPUT115), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT117), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1096), .A2(new_n1097), .A3(new_n1050), .A4(new_n1089), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1058), .A2(new_n1090), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(KEYINPUT116), .A3(new_n691), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT116), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1089), .B1(new_n1096), .B2(new_n1050), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n651), .ZN(new_n1103));
  AOI221_X4 g0903(.A(new_n1079), .B1(new_n1091), .B2(new_n1098), .C1(new_n1100), .C2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1091), .A2(new_n1098), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT118), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1078), .B1(new_n1104), .B2(new_n1107), .ZN(G378));
  NAND2_X1  g0908(.A1(new_n886), .A2(KEYINPUT40), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n889), .A2(new_n890), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1083), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n878), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n856), .B(new_n877), .C1(new_n891), .C2(new_n1083), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n287), .A2(new_n836), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT55), .Z(new_n1115));
  AND2_X1   g0915(.A1(new_n302), .A2(KEYINPUT120), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n302), .A2(KEYINPUT120), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n302), .A2(KEYINPUT120), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1115), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n302), .A2(KEYINPUT120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1118), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1112), .A2(new_n1113), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n1127), .A2(new_n1128), .A3(new_n693), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n386), .A2(new_n253), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1130), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT119), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n556), .A2(new_n781), .B1(new_n722), .B2(new_n522), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n905), .B(new_n1133), .C1(G77), .C2(new_n755), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n734), .A2(new_n389), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1130), .B1(G283), .B2(new_n725), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n779), .A2(G107), .B1(new_n740), .B2(new_n467), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1132), .B1(new_n1140), .B2(KEYINPUT58), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n737), .A2(new_n1074), .B1(new_n739), .B2(new_n782), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n721), .A2(G125), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n717), .B2(new_n1069), .C1(new_n781), .C2(new_n788), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(G150), .C2(new_n744), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1146), .A2(KEYINPUT59), .ZN(new_n1147));
  AOI211_X1 g0947(.A(G33), .B(G41), .C1(new_n725), .C2(G124), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT59), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1148), .B1(new_n908), .B2(new_n734), .C1(new_n1145), .C2(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1141), .B1(KEYINPUT58), .B2(new_n1140), .C1(new_n1147), .C2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n707), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n778), .B1(new_n803), .B2(new_n202), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(new_n1126), .C2(new_n700), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1129), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n879), .A2(new_n1088), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(KEYINPUT57), .C1(new_n1158), .C2(new_n1102), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n691), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1158), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1099), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT57), .B1(new_n1162), .B2(new_n1157), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1156), .B1(new_n1160), .B2(new_n1163), .ZN(G375));
  INV_X1    g0964(.A(new_n1087), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n1158), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n951), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n1167), .A3(new_n1089), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n910), .A2(new_n258), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT122), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G107), .A2(new_n740), .B1(new_n725), .B2(G303), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n989), .B2(new_n737), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n981), .B1(new_n781), .B2(new_n522), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n722), .A2(new_n792), .B1(new_n717), .B2(new_n556), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1170), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n728), .A2(new_n1070), .B1(new_n755), .B2(G159), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n202), .B2(new_n743), .C1(new_n788), .C2(new_n722), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n258), .B1(new_n724), .B2(new_n1074), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n737), .A2(new_n911), .B1(new_n739), .B2(new_n272), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1177), .A2(new_n1135), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n707), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n778), .B1(new_n803), .B2(new_n216), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n888), .C2(new_n800), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1165), .B2(new_n693), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1168), .A2(new_n1185), .ZN(G381));
  OR3_X1    g0986(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1187));
  NOR4_X1   g0987(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(G375), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT116), .B1(new_n1099), .B2(new_n691), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1102), .A2(new_n1101), .A3(new_n651), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1106), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1192), .A2(new_n1078), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1188), .A2(new_n1189), .A3(new_n1193), .ZN(G407));
  NAND2_X1  g0994(.A1(new_n631), .A2(G213), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1189), .A2(new_n1193), .A3(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(G407), .A2(G213), .A3(new_n1197), .ZN(G409));
  XNOR2_X1  g0998(.A(G393), .B(new_n762), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(G390), .A2(new_n964), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(G390), .A2(new_n964), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1200), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1203), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1165), .A2(new_n1158), .A3(KEYINPUT60), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n691), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1089), .A2(KEYINPUT60), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n1166), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1184), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  OR3_X1    g1013(.A1(new_n1213), .A2(KEYINPUT125), .A3(G384), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT125), .B1(new_n1213), .B2(G384), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1213), .A2(G384), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(KEYINPUT124), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT124), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1213), .A2(new_n1219), .A3(G384), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1216), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1192), .A2(new_n1079), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1105), .A2(KEYINPUT118), .A3(new_n1106), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G375), .B1(new_n1225), .B2(new_n1078), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT123), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1129), .B2(new_n1155), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1126), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1112), .A2(new_n1113), .A3(new_n1126), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(KEYINPUT123), .B(new_n1154), .C1(new_n1233), .C2(new_n693), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1157), .B(new_n1167), .C1(new_n1158), .C2(new_n1102), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1228), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1236), .A2(new_n1078), .A3(new_n1192), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1195), .B(new_n1222), .C1(new_n1226), .C2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT126), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G378), .A2(new_n1189), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1237), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1243), .A2(KEYINPUT126), .A3(new_n1195), .A4(new_n1222), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT62), .B1(new_n1240), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1196), .A2(G2897), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1216), .A2(new_n1221), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1216), .A2(new_n1221), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1246), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1237), .B1(G378), .B2(new_n1189), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1247), .B(new_n1250), .C1(new_n1251), .C2(new_n1196), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1251), .A2(new_n1196), .A3(new_n1248), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT62), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1252), .B(new_n1253), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1207), .B1(new_n1245), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT63), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1240), .A2(new_n1258), .A3(new_n1244), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1207), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1254), .A2(KEYINPUT63), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1257), .A2(new_n1263), .ZN(G405));
  AOI21_X1  g1064(.A(new_n1226), .B1(G375), .B2(new_n1193), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1207), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1207), .A2(new_n1265), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1248), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1222), .A3(new_n1267), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(G402));
endmodule


