//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G69), .Z(G235));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G236), .A3(G237), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n467), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n471), .A2(new_n473), .A3(G137), .A4(new_n469), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT70), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n467), .A2(new_n476), .A3(G137), .A4(new_n469), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n470), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n471), .A2(new_n473), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n469), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n485));
  OR3_X1    g060(.A1(new_n485), .A2(G100), .A3(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(G100), .B2(G2105), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n469), .A2(G112), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n486), .A2(new_n487), .A3(G2104), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n482), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND4_X1  g066(.A1(new_n471), .A2(new_n473), .A3(G126), .A4(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n471), .A2(new_n473), .A3(G138), .A4(new_n469), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n467), .A2(new_n500), .A3(G138), .A4(new_n469), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT72), .A3(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(new_n507), .B1(KEYINPUT5), .B2(new_n504), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(G543), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(G75), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n506), .A2(KEYINPUT72), .A3(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(KEYINPUT72), .B1(new_n506), .B2(G543), .ZN(new_n520));
  OAI211_X1 g095(.A(G62), .B(new_n518), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n517), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n508), .A2(KEYINPUT73), .A3(G62), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n516), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n515), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI211_X1 g102(.A(KEYINPUT74), .B(new_n516), .C1(new_n523), .C2(new_n524), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(G166));
  INV_X1    g104(.A(new_n513), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT75), .B(G89), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n510), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n516), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n510), .A2(new_n541), .B1(new_n542), .B2(new_n513), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  NAND3_X1  g119(.A1(new_n509), .A2(G43), .A3(G543), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n510), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n508), .A2(G56), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n516), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(G188));
  NAND3_X1  g132(.A1(new_n508), .A2(G91), .A3(new_n509), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(KEYINPUT76), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT6), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n560), .A2(new_n561), .A3(new_n563), .A4(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n509), .A2(new_n566), .A3(G543), .A4(new_n560), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n558), .B(new_n568), .C1(new_n569), .C2(new_n516), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  NAND2_X1  g147(.A1(new_n521), .A2(new_n522), .ZN(new_n573));
  INV_X1    g148(.A(new_n517), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n573), .A2(new_n524), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n514), .B1(new_n576), .B2(KEYINPUT74), .ZN(new_n577));
  INV_X1    g152(.A(new_n528), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT77), .B1(new_n527), .B2(new_n528), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G303));
  NAND2_X1  g157(.A1(new_n530), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n510), .ZN(G288));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  INV_X1    g162(.A(G48), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n510), .A2(new_n587), .B1(new_n588), .B2(new_n513), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n508), .A2(G61), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT78), .Z(new_n592));
  AOI21_X1  g167(.A(new_n516), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n589), .A2(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(G72), .A2(G543), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n505), .A2(new_n507), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(new_n518), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G651), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n510), .ZN(new_n603));
  XOR2_X1   g178(.A(KEYINPUT80), .B(G47), .Z(new_n604));
  AOI22_X1  g179(.A1(new_n603), .A2(G85), .B1(new_n530), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT81), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n596), .A2(G66), .A3(new_n518), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n516), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g186(.A1(new_n509), .A2(G54), .A3(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n612), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n615));
  OAI211_X1 g190(.A(KEYINPUT81), .B(new_n614), .C1(new_n615), .C2(new_n516), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n603), .A2(KEYINPUT10), .A3(G92), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  INV_X1    g194(.A(G92), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n510), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n607), .B1(new_n624), .B2(G868), .ZN(G321));
  XNOR2_X1  g200(.A(G321), .B(KEYINPUT82), .ZN(G284));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(G299), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G168), .B2(new_n627), .ZN(G297));
  OAI21_X1  g204(.A(new_n628), .B1(G168), .B2(new_n627), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(G148));
  AOI22_X1  g207(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n633));
  OAI221_X1 g208(.A(new_n545), .B1(new_n510), .B2(new_n546), .C1(new_n633), .C2(new_n516), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(new_n627), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n623), .A2(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n467), .A2(new_n465), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT13), .Z(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n483), .A2(G123), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n481), .A2(G135), .ZN(new_n644));
  OR2_X1    g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n645), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2096), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n641), .A2(G2100), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n642), .A2(new_n648), .A3(new_n649), .ZN(G156));
  INV_X1    g225(.A(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT83), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2430), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT14), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n654), .A2(new_n655), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n651), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n657), .A2(new_n658), .ZN(new_n663));
  AOI21_X1  g238(.A(KEYINPUT84), .B1(new_n656), .B2(KEYINPUT14), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n651), .B(new_n660), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2451), .B(G2454), .Z(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n666), .B(new_n667), .Z(new_n668));
  NAND3_X1  g243(.A1(new_n662), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n668), .ZN(new_n670));
  INV_X1    g245(.A(new_n665), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n670), .B1(new_n661), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1341), .B(G1348), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n669), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n674), .B1(new_n669), .B2(new_n672), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT85), .ZN(new_n677));
  OAI211_X1 g252(.A(G14), .B(new_n675), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(G401));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2067), .B(G2678), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2072), .B(G2078), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT18), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  AND3_X1   g263(.A1(new_n688), .A2(KEYINPUT17), .A3(new_n685), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n685), .B1(new_n688), .B2(KEYINPUT17), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n689), .A2(new_n690), .A3(new_n684), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G2096), .B(G2100), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G227));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1956), .B(G2474), .Z(new_n699));
  XOR2_X1   g274(.A(G1961), .B(G1966), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1971), .B(G1976), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT19), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n699), .A2(new_n700), .A3(KEYINPUT86), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n703), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(new_n706), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n699), .A2(new_n700), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n712), .A2(new_n713), .A3(new_n701), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n710), .A2(new_n711), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(G1991), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(G1991), .ZN(new_n718));
  AOI21_X1  g293(.A(G1996), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(G1996), .A3(new_n718), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n698), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n721), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n723), .A2(new_n697), .A3(new_n719), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n696), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n697), .B1(new_n723), .B2(new_n719), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n720), .A2(new_n698), .A3(new_n721), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n726), .A2(new_n727), .A3(new_n695), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n725), .A2(new_n728), .ZN(G229));
  NAND2_X1  g304(.A1(G168), .A2(G16), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G16), .B2(G21), .ZN(new_n731));
  INV_X1    g306(.A(G1966), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT98), .Z(new_n734));
  NOR2_X1   g309(.A1(G5), .A2(G16), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G171), .B2(G16), .ZN(new_n736));
  INV_X1    g311(.A(G1961), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G29), .A2(G35), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G162), .B2(G29), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2090), .ZN(new_n744));
  NOR2_X1   g319(.A1(G16), .A2(G19), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n551), .B2(G16), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(G1341), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT31), .B(G11), .Z(new_n749));
  INV_X1    g324(.A(G28), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n750), .A2(KEYINPUT30), .ZN(new_n751));
  AOI21_X1  g326(.A(G29), .B1(new_n750), .B2(KEYINPUT30), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G29), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n465), .A2(G105), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n471), .A2(new_n473), .A3(G129), .A4(G2105), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n471), .A2(new_n473), .A3(G141), .A4(new_n469), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G29), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G29), .B2(G32), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT27), .B(G1996), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n753), .B1(new_n754), .B2(new_n647), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n764), .B2(new_n765), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n754), .A2(G27), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n754), .ZN(new_n769));
  INV_X1    g344(.A(G2084), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT24), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n754), .B1(new_n771), .B2(G34), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT97), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n772), .A2(new_n773), .B1(new_n771), .B2(G34), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n773), .B2(new_n772), .ZN(new_n775));
  INV_X1    g350(.A(G160), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n754), .ZN(new_n777));
  OAI221_X1 g352(.A(new_n767), .B1(G2078), .B2(new_n769), .C1(new_n770), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n731), .A2(new_n732), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n777), .A2(new_n770), .B1(new_n769), .B2(G2078), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n739), .A2(new_n748), .A3(new_n778), .A4(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G299), .ZN(new_n783));
  INV_X1    g358(.A(G16), .ZN(new_n784));
  OAI21_X1  g359(.A(KEYINPUT23), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(G20), .ZN(new_n786));
  MUX2_X1   g361(.A(KEYINPUT23), .B(new_n785), .S(new_n786), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G1956), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n754), .A2(G33), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n481), .A2(G139), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT95), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n465), .A2(G103), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT25), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(G115), .A2(G2104), .ZN(new_n796));
  INV_X1    g371(.A(G127), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n480), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G2105), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n790), .B1(new_n792), .B2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n791), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n803), .A2(KEYINPUT96), .A3(new_n799), .A4(new_n795), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n789), .B1(new_n805), .B2(new_n754), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(G2072), .Z(new_n807));
  OR2_X1    g382(.A1(new_n787), .A2(G1956), .ZN(new_n808));
  INV_X1    g383(.A(G26), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(G29), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n471), .A2(new_n473), .A3(G140), .A4(new_n469), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT94), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n467), .A2(KEYINPUT94), .A3(G140), .A4(new_n469), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n467), .A2(G128), .A3(G2105), .ZN(new_n815));
  OR2_X1    g390(.A1(G104), .A2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n810), .B1(new_n818), .B2(G29), .ZN(new_n819));
  MUX2_X1   g394(.A(new_n810), .B(new_n819), .S(KEYINPUT28), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2067), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n807), .A2(new_n808), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(G4), .A2(G16), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT93), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n623), .B2(new_n784), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1348), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n782), .A2(new_n788), .A3(new_n822), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT32), .B(G1981), .Z(new_n829));
  NAND2_X1  g404(.A1(G305), .A2(G16), .ZN(new_n830));
  INV_X1    g405(.A(G6), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(G16), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n829), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n829), .ZN(new_n835));
  AOI211_X1 g410(.A(new_n832), .B(new_n835), .C1(G305), .C2(G16), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(G16), .A2(G23), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G288), .B2(new_n784), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT33), .B(G1976), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT89), .B(G1971), .ZN(new_n843));
  NAND2_X1  g418(.A1(G166), .A2(G16), .ZN(new_n844));
  OR2_X1    g419(.A1(G16), .A2(G22), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n844), .A2(new_n845), .A3(new_n843), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n842), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT34), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT90), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n844), .A2(new_n845), .A3(new_n843), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n837), .B(new_n841), .C1(new_n852), .C2(new_n846), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT90), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT34), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT92), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n784), .A2(G24), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(G290), .B2(G16), .ZN(new_n859));
  INV_X1    g434(.A(G1986), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n467), .A2(G2105), .ZN(new_n863));
  INV_X1    g438(.A(G119), .ZN(new_n864));
  OR3_X1    g439(.A1(new_n863), .A2(KEYINPUT88), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT88), .B1(new_n863), .B2(new_n864), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n481), .A2(G131), .ZN(new_n867));
  OR2_X1    g442(.A1(G95), .A2(G2105), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  MUX2_X1   g445(.A(G25), .B(new_n870), .S(G29), .Z(new_n871));
  XNOR2_X1  g446(.A(KEYINPUT35), .B(G1991), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n871), .B(new_n872), .Z(new_n873));
  NAND3_X1  g448(.A1(new_n861), .A2(new_n862), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n850), .B2(new_n849), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n856), .A2(new_n857), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n857), .B1(new_n856), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n828), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n849), .A2(KEYINPUT90), .A3(new_n850), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n854), .B1(new_n853), .B2(KEYINPUT34), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT92), .ZN(new_n883));
  INV_X1    g458(.A(new_n828), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n884), .A3(new_n876), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n827), .B1(new_n879), .B2(new_n885), .ZN(G311));
  INV_X1    g461(.A(new_n827), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n883), .A2(new_n884), .A3(new_n876), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n884), .B1(new_n883), .B2(new_n876), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(G150));
  NOR2_X1   g465(.A1(new_n623), .A2(new_n631), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n596), .A2(G93), .A3(new_n518), .A4(new_n509), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n509), .A2(G55), .A3(G543), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n894), .B(KEYINPUT100), .C1(new_n516), .C2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n596), .A2(G67), .A3(new_n518), .ZN(new_n898));
  NAND2_X1  g473(.A1(G80), .A2(G543), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n516), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n892), .A2(new_n893), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n896), .A2(new_n634), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n900), .A2(new_n901), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n551), .A2(KEYINPUT100), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n891), .B(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n908));
  AOI21_X1  g483(.A(G860), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n908), .B2(new_n907), .ZN(new_n910));
  INV_X1    g485(.A(new_n904), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(G860), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(KEYINPUT37), .Z(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT101), .ZN(G145));
  XOR2_X1   g490(.A(new_n870), .B(KEYINPUT107), .Z(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n647), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n647), .A2(new_n918), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(G160), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n776), .A3(new_n920), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(G162), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n490), .A3(new_n923), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n801), .A2(new_n804), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n762), .A2(new_n818), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n815), .A2(new_n817), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(new_n761), .A3(new_n814), .A4(new_n813), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n497), .A2(KEYINPUT103), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n492), .A2(new_n933), .A3(new_n496), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n932), .A2(new_n934), .B1(new_n499), .B2(new_n501), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n929), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n929), .A2(new_n931), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n499), .A2(new_n501), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n492), .A2(new_n933), .A3(new_n496), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n933), .B1(new_n492), .B2(new_n496), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n928), .A2(new_n936), .A3(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n929), .A2(new_n931), .A3(new_n935), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n935), .B1(new_n929), .B2(new_n931), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT104), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(new_n947), .A3(new_n936), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n928), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI211_X1 g526(.A(KEYINPUT105), .B(new_n928), .C1(new_n946), .C2(new_n948), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n927), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n946), .A2(new_n948), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n805), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT105), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n949), .A2(new_n950), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n922), .A2(new_n490), .A3(new_n923), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n490), .B1(new_n922), .B2(new_n923), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n956), .A2(new_n957), .A3(new_n943), .A4(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n640), .B(KEYINPUT106), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n483), .A2(G130), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n481), .A2(G142), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n469), .A2(G118), .ZN(new_n965));
  OAI21_X1  g540(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n963), .B(new_n964), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n962), .B(new_n967), .Z(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n953), .A2(new_n961), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n953), .B2(new_n961), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n917), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n943), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n955), .B2(KEYINPUT105), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n960), .B1(new_n974), .B2(new_n957), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n951), .A2(new_n952), .A3(new_n927), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n968), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n953), .A2(new_n961), .A3(new_n969), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n916), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G37), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n972), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT40), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT40), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n972), .A2(new_n979), .A3(new_n983), .A4(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(G395));
  NAND2_X1  g560(.A1(new_n911), .A2(new_n627), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n988));
  XNOR2_X1  g563(.A(G290), .B(G305), .ZN(new_n989));
  INV_X1    g564(.A(G288), .ZN(new_n990));
  XNOR2_X1  g565(.A(G166), .B(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n589), .A2(new_n593), .ZN(new_n993));
  XNOR2_X1  g568(.A(G290), .B(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(G166), .B(G288), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n988), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n992), .A2(new_n996), .A3(KEYINPUT109), .A4(KEYINPUT42), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n636), .B(new_n906), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n617), .A2(G299), .A3(new_n622), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G299), .B1(new_n617), .B2(new_n622), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT41), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n623), .A2(new_n783), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1003), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1007), .B1(new_n1002), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n987), .B1(new_n1001), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1001), .A2(new_n1015), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n999), .A2(new_n1014), .A3(KEYINPUT110), .A4(new_n1000), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n986), .B1(new_n1019), .B2(new_n627), .ZN(G295));
  OAI21_X1  g595(.A(new_n986), .B1(new_n1019), .B2(new_n627), .ZN(G331));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT43), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n906), .A2(G171), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n903), .A2(new_n905), .A3(G301), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(G168), .A3(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n903), .A2(G301), .A3(new_n905), .ZN(new_n1027));
  AOI21_X1  g602(.A(G301), .B1(new_n903), .B2(new_n905), .ZN(new_n1028));
  OAI21_X1  g603(.A(G286), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1013), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1006), .B1(new_n1029), .B2(new_n1026), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(KEYINPUT111), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n1033));
  AOI211_X1 g608(.A(new_n1033), .B(new_n1006), .C1(new_n1029), .C2(new_n1026), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(G37), .B1(new_n1035), .B2(new_n997), .ZN(new_n1036));
  INV_X1    g611(.A(new_n997), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1023), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1010), .A2(new_n1003), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1027), .A2(new_n1028), .A3(G286), .ZN(new_n1041));
  AOI21_X1  g616(.A(G168), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n1033), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1031), .A2(KEYINPUT111), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1044), .A2(new_n997), .A3(new_n1045), .A4(new_n1030), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1029), .A2(new_n1026), .A3(new_n1011), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1040), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1006), .A2(new_n1049), .A3(KEYINPUT41), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT112), .B1(new_n1040), .B2(new_n1008), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(new_n1026), .A4(new_n1029), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n1037), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1046), .A2(new_n1054), .A3(new_n980), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(KEYINPUT43), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1022), .B1(new_n1039), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1036), .A2(new_n1058), .A3(new_n1023), .A4(new_n1038), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1022), .B1(new_n1055), .B2(KEYINPUT43), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1038), .A2(new_n1046), .A3(new_n1023), .A4(new_n980), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT113), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1057), .A2(new_n1063), .ZN(G397));
  INV_X1    g639(.A(G1384), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT45), .B1(new_n941), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G113), .A2(G2104), .ZN(new_n1068));
  INV_X1    g643(.A(G125), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1068), .B1(new_n480), .B2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1070), .A2(G2105), .B1(G101), .B2(new_n465), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1071), .A2(G40), .A3(new_n475), .A4(new_n477), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n870), .B(new_n872), .ZN(new_n1074));
  INV_X1    g649(.A(G2067), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n818), .B(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1996), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n761), .B(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1073), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(G290), .B(new_n860), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1073), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(new_n1083), .B(KEYINPUT114), .Z(new_n1084));
  INV_X1    g659(.A(G8), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G168), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT45), .ZN(new_n1087));
  NOR3_X1   g662(.A1(G164), .A2(new_n1087), .A3(G1384), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1066), .A2(new_n1088), .A3(new_n1072), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n941), .A2(new_n1090), .A3(new_n1065), .ZN(new_n1091));
  INV_X1    g666(.A(G40), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n470), .A2(new_n1092), .A3(new_n478), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1089), .A2(G1966), .B1(G2084), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1086), .B1(new_n1096), .B2(G8), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT51), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1086), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1100), .B(G8), .C1(new_n1096), .C2(G286), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n497), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n938), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(new_n1090), .A3(new_n1065), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT50), .B1(new_n935), .B2(G1384), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1105), .A2(KEYINPUT116), .A3(new_n1090), .A4(new_n1065), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1093), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G1956), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n941), .A2(KEYINPUT45), .A3(new_n1065), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1087), .B1(G164), .B2(G1384), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1113), .A2(new_n1093), .A3(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1111), .A2(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n596), .A2(G65), .A3(new_n518), .ZN(new_n1118));
  NAND2_X1  g693(.A1(G78), .A2(G543), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n516), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n558), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT120), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1123), .B(new_n558), .C1(new_n569), .C2(new_n516), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1122), .A2(new_n568), .A3(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(KEYINPUT57), .A4(new_n568), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT121), .B1(G299), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1127), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1117), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1117), .A2(new_n1134), .ZN(new_n1136));
  INV_X1    g711(.A(G1348), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1095), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n941), .A2(new_n1065), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1139), .A2(new_n1072), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1075), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n623), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1135), .B1(new_n1136), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1144), .A2(new_n1134), .A3(KEYINPUT123), .A4(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT61), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1113), .A2(new_n1093), .A3(new_n1114), .A4(new_n1077), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT58), .B(G1341), .Z(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1139), .B2(new_n1072), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n551), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(KEYINPUT122), .A3(new_n551), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(KEYINPUT59), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT122), .B1(new_n1151), .B2(new_n551), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1095), .A2(new_n1137), .B1(new_n1140), .B2(new_n1075), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n623), .A2(KEYINPUT60), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1157), .A2(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1138), .A2(new_n623), .A3(new_n1141), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT60), .B1(new_n1162), .B2(new_n1142), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1156), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1143), .B1(new_n1147), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n579), .B1(new_n577), .B2(new_n578), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n527), .A2(KEYINPUT77), .A3(new_n528), .ZN(new_n1167));
  OAI21_X1  g742(.A(G8), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT55), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1072), .B1(new_n1139), .B2(KEYINPUT50), .ZN(new_n1172));
  INV_X1    g747(.A(G2090), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1172), .A2(new_n1173), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1113), .A2(new_n1093), .A3(new_n1114), .ZN(new_n1175));
  INV_X1    g750(.A(G1971), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1174), .A2(KEYINPUT117), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(G8), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT117), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1170), .B(new_n1171), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n1095), .A2(G2090), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1085), .B1(new_n1182), .B2(new_n1177), .ZN(new_n1183));
  AOI21_X1  g758(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1184));
  AOI211_X1 g759(.A(new_n1169), .B(new_n1085), .C1(new_n580), .C2(new_n581), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(G1976), .ZN(new_n1187));
  OAI221_X1 g762(.A(G8), .B1(G288), .B2(new_n1187), .C1(new_n1139), .C2(new_n1072), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(KEYINPUT52), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT52), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1190), .B1(new_n990), .B2(G1976), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1189), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(G305), .A2(G1981), .ZN(new_n1193));
  INV_X1    g768(.A(G1981), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n993), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1193), .A2(KEYINPUT49), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT115), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1193), .A2(KEYINPUT115), .A3(KEYINPUT49), .A4(new_n1195), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(KEYINPUT49), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1201));
  OAI21_X1  g776(.A(G8), .B1(new_n1139), .B2(new_n1072), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1192), .B1(new_n1200), .B2(new_n1203), .ZN(new_n1204));
  AND3_X1   g779(.A1(new_n1181), .A2(new_n1186), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(G2078), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1113), .A2(new_n1093), .A3(new_n1114), .A4(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT53), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1209), .A2(KEYINPUT124), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1207), .A2(new_n1211), .A3(new_n1208), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  AND3_X1   g788(.A1(new_n1095), .A2(KEYINPUT125), .A3(new_n737), .ZN(new_n1214));
  AOI21_X1  g789(.A(KEYINPUT125), .B1(new_n1095), .B2(new_n737), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1067), .A2(new_n1217), .A3(new_n1093), .ZN(new_n1218));
  OAI21_X1  g793(.A(KEYINPUT126), .B1(new_n1066), .B2(new_n1072), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1208), .A2(G2078), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n1218), .A2(new_n1219), .A3(new_n1113), .A4(new_n1220), .ZN(new_n1221));
  NAND4_X1  g796(.A1(new_n1213), .A2(new_n1216), .A3(G301), .A4(new_n1221), .ZN(new_n1222));
  AOI22_X1  g797(.A1(new_n1089), .A2(new_n1220), .B1(new_n737), .B2(new_n1095), .ZN(new_n1223));
  AND3_X1   g798(.A1(new_n1207), .A2(new_n1211), .A3(new_n1208), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1211), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1223), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1226), .A2(G171), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1222), .A2(new_n1227), .A3(KEYINPUT127), .ZN(new_n1228));
  INV_X1    g803(.A(KEYINPUT54), .ZN(new_n1229));
  INV_X1    g804(.A(new_n1215), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1095), .A2(KEYINPUT125), .A3(new_n737), .ZN(new_n1231));
  AND3_X1   g806(.A1(new_n1221), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1233));
  NAND4_X1  g808(.A1(new_n1232), .A2(new_n1233), .A3(G301), .A4(new_n1213), .ZN(new_n1234));
  NAND3_X1  g809(.A1(new_n1228), .A2(new_n1229), .A3(new_n1234), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1213), .A2(G301), .A3(new_n1223), .ZN(new_n1236));
  AND3_X1   g811(.A1(new_n1213), .A2(new_n1221), .A3(new_n1216), .ZN(new_n1237));
  OAI211_X1 g812(.A(new_n1236), .B(KEYINPUT54), .C1(new_n1237), .C2(G301), .ZN(new_n1238));
  NAND4_X1  g813(.A1(new_n1165), .A2(new_n1205), .A3(new_n1235), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g814(.A(new_n1227), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1102), .A2(KEYINPUT62), .ZN(new_n1241));
  NAND3_X1  g816(.A1(new_n1205), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AOI21_X1  g817(.A(new_n1103), .B1(new_n1239), .B2(new_n1242), .ZN(new_n1243));
  AND3_X1   g818(.A1(new_n1096), .A2(G8), .A3(G168), .ZN(new_n1244));
  NAND4_X1  g819(.A1(new_n1181), .A2(new_n1186), .A3(new_n1204), .A4(new_n1244), .ZN(new_n1245));
  INV_X1    g820(.A(KEYINPUT63), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OR2_X1    g822(.A1(new_n1183), .A2(KEYINPUT118), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1183), .A2(KEYINPUT118), .ZN(new_n1249));
  NAND4_X1  g824(.A1(new_n1248), .A2(new_n1249), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1250));
  AND2_X1   g825(.A1(new_n1244), .A2(KEYINPUT63), .ZN(new_n1251));
  NAND4_X1  g826(.A1(new_n1250), .A2(new_n1186), .A3(new_n1204), .A4(new_n1251), .ZN(new_n1252));
  NAND2_X1  g827(.A1(new_n1247), .A2(new_n1252), .ZN(new_n1253));
  NAND4_X1  g828(.A1(new_n1205), .A2(KEYINPUT62), .A3(new_n1103), .A4(new_n1240), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1255));
  NAND3_X1  g830(.A1(new_n1255), .A2(new_n1187), .A3(new_n990), .ZN(new_n1256));
  AOI21_X1  g831(.A(new_n1202), .B1(new_n1256), .B2(new_n1195), .ZN(new_n1257));
  INV_X1    g832(.A(new_n1186), .ZN(new_n1258));
  AOI21_X1  g833(.A(new_n1257), .B1(new_n1258), .B2(new_n1204), .ZN(new_n1259));
  NAND3_X1  g834(.A1(new_n1253), .A2(new_n1254), .A3(new_n1259), .ZN(new_n1260));
  OAI21_X1  g835(.A(new_n1084), .B1(new_n1243), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g836(.A(KEYINPUT48), .ZN(new_n1262));
  NOR2_X1   g837(.A1(G290), .A2(G1986), .ZN(new_n1263));
  INV_X1    g838(.A(new_n1263), .ZN(new_n1264));
  OAI21_X1  g839(.A(new_n1262), .B1(new_n1264), .B2(new_n1082), .ZN(new_n1265));
  NAND3_X1  g840(.A1(new_n1263), .A2(KEYINPUT48), .A3(new_n1073), .ZN(new_n1266));
  AND3_X1   g841(.A1(new_n1265), .A2(new_n1080), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g842(.A(new_n1082), .B1(new_n762), .B2(new_n1076), .ZN(new_n1268));
  AND3_X1   g843(.A1(new_n1073), .A2(KEYINPUT46), .A3(new_n1077), .ZN(new_n1269));
  AOI21_X1  g844(.A(KEYINPUT46), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1270));
  NOR3_X1   g845(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g846(.A(new_n1271), .B(KEYINPUT47), .ZN(new_n1272));
  OR2_X1    g847(.A1(new_n870), .A2(new_n872), .ZN(new_n1273));
  OAI22_X1  g848(.A1(new_n1079), .A2(new_n1273), .B1(G2067), .B2(new_n818), .ZN(new_n1274));
  AOI211_X1 g849(.A(new_n1267), .B(new_n1272), .C1(new_n1073), .C2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g850(.A1(new_n1261), .A2(new_n1275), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g851(.A1(new_n1039), .A2(new_n1056), .ZN(new_n1278));
  NOR2_X1   g852(.A1(G227), .A2(new_n462), .ZN(new_n1279));
  OAI21_X1  g853(.A(new_n1279), .B1(new_n678), .B2(new_n679), .ZN(new_n1280));
  NOR2_X1   g854(.A1(new_n1280), .A2(G229), .ZN(new_n1281));
  NAND2_X1  g855(.A1(new_n981), .A2(new_n1281), .ZN(new_n1282));
  NOR2_X1   g856(.A1(new_n1278), .A2(new_n1282), .ZN(G308));
  OAI211_X1 g857(.A(new_n981), .B(new_n1281), .C1(new_n1039), .C2(new_n1056), .ZN(G225));
endmodule


