//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  AOI22_X1  g039(.A1(G101), .A2(new_n460), .B1(new_n464), .B2(G137), .ZN(new_n465));
  INV_X1    g040(.A(new_n463), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n468), .B(KEYINPUT65), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n458), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(KEYINPUT66), .ZN(new_n471));
  XOR2_X1   g046(.A(new_n468), .B(KEYINPUT65), .Z(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n463), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n465), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT68), .ZN(G160));
  NAND2_X1  g054(.A1(new_n464), .A2(G136), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n463), .A2(new_n458), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND2_X1  g063(.A1(new_n485), .A2(G126), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n458), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n464), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT4), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n464), .A2(new_n497), .A3(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n496), .B2(new_n498), .ZN(G164));
  AND3_X1   g074(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n500));
  AOI21_X1  g075(.A(G543), .B1(KEYINPUT70), .B2(KEYINPUT5), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(KEYINPUT71), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n500), .A2(new_n501), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n512), .A2(G543), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n520), .A2(G651), .B1(new_n521), .B2(G50), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n516), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n515), .A2(G89), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n526));
  AND3_X1   g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(KEYINPUT73), .B1(new_n512), .B2(G543), .ZN(new_n528));
  OAI211_X1 g103(.A(KEYINPUT73), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT74), .B(G51), .Z(new_n532));
  OAI221_X1 g107(.A(new_n525), .B1(new_n526), .B2(new_n527), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n518), .A2(KEYINPUT72), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n511), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n537), .A3(G63), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n526), .A2(G76), .A3(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n534), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n533), .A2(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n535), .A2(new_n537), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G651), .ZN(new_n546));
  INV_X1    g121(.A(new_n531), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G52), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n515), .A2(G90), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n552), .A2(new_n531), .B1(new_n514), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n535), .A2(new_n537), .A3(G56), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n534), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n521), .A2(new_n564), .A3(G53), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n512), .A2(G53), .A3(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n565), .A2(new_n570), .A3(new_n567), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n504), .A2(new_n505), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT71), .B1(new_n511), .B2(new_n512), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT77), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n506), .A2(new_n576), .A3(new_n513), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(G91), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n511), .A2(G65), .ZN(new_n579));
  NAND2_X1  g154(.A1(G78), .A2(G543), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT78), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n572), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G299));
  INV_X1    g159(.A(G168), .ZN(G286));
  AND2_X1   g160(.A1(new_n575), .A2(new_n577), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G87), .ZN(new_n587));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n534), .B1(new_n543), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(G49), .B2(new_n521), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(new_n521), .A2(G48), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n518), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n592), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n597), .B2(new_n596), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n586), .A2(G86), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G60), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n543), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n515), .A2(G85), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT80), .B(G47), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n547), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n518), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n547), .A2(G54), .B1(G651), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n575), .A2(G92), .A3(new_n577), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(KEYINPUT81), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n575), .A2(new_n618), .A3(G92), .A4(new_n577), .ZN(new_n619));
  AND3_X1   g194(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n617), .B1(new_n616), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n610), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n610), .B1(new_n623), .B2(G868), .ZN(G321));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(G299), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n626), .B2(G168), .ZN(G297));
  OAI21_X1  g203(.A(new_n627), .B1(new_n626), .B2(G168), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n623), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n623), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n460), .A2(new_n466), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT13), .Z(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2100), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n464), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n485), .A2(G123), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n458), .A2(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n640), .A2(new_n641), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1341), .B(G1348), .Z(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT84), .ZN(G401));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT85), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2084), .B(G2090), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n671), .B1(new_n667), .B2(new_n670), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n669), .B2(new_n670), .ZN(new_n674));
  INV_X1    g249(.A(new_n670), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n675), .A2(new_n671), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n667), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  OR3_X1    g253(.A1(new_n672), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n688), .A2(new_n689), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(new_n695), .B(new_n694), .S(new_n687), .Z(new_n696));
  NOR2_X1   g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1991), .B(G1996), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n699), .A2(new_n700), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n699), .A2(new_n700), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G229));
  AND2_X1   g284(.A1(new_n599), .A2(new_n600), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G16), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G6), .B2(G16), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT32), .B(G1981), .Z(new_n713));
  AND2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n716), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1971), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n714), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G23), .B(G288), .S(G16), .Z(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT33), .B(G1976), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(KEYINPUT90), .ZN(new_n724));
  INV_X1    g299(.A(new_n722), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n721), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT90), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n720), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G25), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT88), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n464), .A2(G131), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n485), .A2(G119), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n458), .A2(G107), .ZN(new_n737));
  OAI21_X1  g312(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n735), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT89), .Z(new_n740));
  AOI21_X1  g315(.A(new_n734), .B1(new_n740), .B2(G29), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT35), .B(G1991), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n744));
  INV_X1    g319(.A(G290), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(new_n716), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n716), .B2(G24), .ZN(new_n747));
  INV_X1    g322(.A(G1986), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n744), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n743), .B(new_n749), .C1(new_n748), .C2(new_n747), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n731), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G29), .A2(G33), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT93), .Z(new_n755));
  NAND3_X1  g330(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT25), .Z(new_n757));
  INV_X1    g332(.A(G139), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n494), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n466), .A2(G127), .ZN(new_n760));
  NAND2_X1  g335(.A1(G115), .A2(G2104), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n458), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n755), .B1(new_n763), .B2(G29), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G2072), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n732), .A2(G27), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G164), .B2(new_n732), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G2078), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n558), .A2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G16), .B2(G19), .ZN(new_n771));
  INV_X1    g346(.A(G1341), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n767), .A2(G2078), .ZN(new_n775));
  NOR4_X1   g350(.A1(new_n769), .A2(new_n773), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n732), .A2(G26), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT28), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n464), .A2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n485), .A2(G128), .ZN(new_n780));
  OR2_X1    g355(.A1(G104), .A2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n781), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n782));
  AND3_X1   g357(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(KEYINPUT92), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(KEYINPUT92), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n778), .B1(new_n786), .B2(G29), .ZN(new_n787));
  INV_X1    g362(.A(G2067), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n732), .A2(G35), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G162), .B2(new_n732), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT29), .B(G2090), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n716), .A2(G5), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G171), .B2(new_n716), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT97), .ZN(new_n797));
  INV_X1    g372(.A(G1961), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(G160), .A2(G29), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT24), .B(G34), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(new_n732), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT94), .Z(new_n803));
  NAND3_X1  g378(.A1(new_n800), .A2(G2084), .A3(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n776), .A2(new_n794), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(G2084), .B1(new_n800), .B2(new_n803), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n732), .A2(G32), .ZN(new_n807));
  NAND3_X1  g382(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT26), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G129), .B2(new_n485), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n460), .A2(G105), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n464), .A2(G141), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(KEYINPUT95), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(KEYINPUT95), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n807), .B1(new_n817), .B2(new_n732), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT27), .Z(new_n819));
  AOI21_X1  g394(.A(new_n806), .B1(new_n819), .B2(G1996), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n716), .A2(G20), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT23), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n583), .B2(new_n716), .ZN(new_n823));
  INV_X1    g398(.A(G1956), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n820), .B(new_n825), .C1(G1996), .C2(new_n819), .ZN(new_n826));
  INV_X1    g401(.A(G1348), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n623), .A2(G16), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G4), .B2(G16), .ZN(new_n829));
  AOI211_X1 g404(.A(new_n805), .B(new_n826), .C1(new_n827), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n716), .A2(G21), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G168), .B2(new_n716), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(G1966), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT96), .Z(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT30), .B(G28), .ZN(new_n835));
  OR2_X1    g410(.A1(KEYINPUT31), .A2(G11), .ZN(new_n836));
  NAND2_X1  g411(.A1(KEYINPUT31), .A2(G11), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n835), .A2(new_n732), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n646), .B2(new_n732), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n832), .B2(G1966), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n834), .B(new_n840), .C1(new_n798), .C2(new_n797), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT98), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n830), .B(new_n842), .C1(new_n827), .C2(new_n829), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n753), .A2(new_n843), .ZN(G311));
  OR2_X1    g419(.A1(new_n753), .A2(new_n843), .ZN(G150));
  NAND2_X1  g420(.A1(new_n623), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  OAI21_X1  g422(.A(G55), .B1(new_n528), .B2(new_n530), .ZN(new_n848));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n514), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n535), .A2(new_n537), .A3(G67), .ZN(new_n851));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n534), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n558), .A2(new_n854), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n554), .A2(new_n557), .B1(new_n850), .B2(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n847), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n859));
  AOI21_X1  g434(.A(G860), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n859), .B2(new_n858), .ZN(new_n861));
  INV_X1    g436(.A(new_n854), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n865), .ZN(G145));
  NAND2_X1  g441(.A1(new_n485), .A2(G130), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n458), .A2(G118), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(G142), .B2(new_n464), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n739), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n638), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n786), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n784), .A2(new_n785), .A3(KEYINPUT101), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n496), .A2(new_n498), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n493), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n490), .A2(new_n491), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n485), .B2(G126), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT100), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n878), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n817), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n814), .B2(new_n815), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n877), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n878), .A2(new_n880), .A3(new_n883), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n816), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n875), .B(new_n876), .C1(new_n890), .C2(new_n886), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n759), .A2(new_n762), .A3(KEYINPUT102), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n888), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n763), .B(KEYINPUT102), .Z(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(new_n888), .B2(new_n891), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n873), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n888), .A2(new_n891), .ZN(new_n897));
  INV_X1    g472(.A(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n888), .A2(new_n891), .A3(new_n892), .ZN(new_n900));
  INV_X1    g475(.A(new_n873), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G160), .B(new_n646), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(G162), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n904), .B(new_n487), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n908));
  OAI22_X1  g483(.A1(new_n893), .A2(new_n895), .B1(new_n908), .B2(new_n873), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n907), .B(new_n909), .C1(new_n902), .C2(new_n908), .ZN(new_n910));
  INV_X1    g485(.A(G37), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g488(.A1(new_n862), .A2(new_n626), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n632), .B(new_n857), .Z(new_n915));
  NAND2_X1  g490(.A1(new_n622), .A2(G299), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n583), .B(new_n614), .C1(new_n620), .C2(new_n621), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n916), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n916), .A2(new_n918), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n916), .A2(KEYINPUT104), .A3(new_n918), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n921), .B1(new_n915), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G305), .A2(new_n745), .ZN(new_n928));
  NAND3_X1  g503(.A1(G290), .A2(new_n599), .A3(new_n600), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G288), .A2(G166), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n587), .A2(G303), .A3(new_n590), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n928), .A2(new_n931), .A3(new_n932), .A4(new_n929), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT42), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n934), .A2(KEYINPUT105), .A3(new_n935), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT105), .B1(new_n934), .B2(new_n935), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n936), .B2(KEYINPUT106), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n938), .B1(new_n943), .B2(KEYINPUT42), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n927), .B(new_n944), .Z(new_n945));
  OAI21_X1  g520(.A(new_n914), .B1(new_n945), .B2(new_n626), .ZN(G295));
  OAI21_X1  g521(.A(new_n914), .B1(new_n945), .B2(new_n626), .ZN(G331));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n855), .A2(G301), .A3(new_n856), .ZN(new_n949));
  AOI21_X1  g524(.A(G301), .B1(new_n855), .B2(new_n856), .ZN(new_n950));
  OAI21_X1  g525(.A(G286), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n857), .A2(G171), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n855), .A2(G301), .A3(new_n856), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(G168), .A3(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n919), .B2(new_n920), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n936), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n939), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n951), .A2(new_n954), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(new_n916), .A3(new_n918), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n956), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n962), .A2(new_n911), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n616), .A2(new_n619), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT10), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n583), .B1(new_n968), .B2(new_n614), .ZN(new_n969));
  INV_X1    g544(.A(new_n918), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT41), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n960), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n955), .A2(new_n922), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n942), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n964), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n924), .A2(new_n925), .A3(new_n960), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n971), .B2(new_n972), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n955), .B1(new_n920), .B2(KEYINPUT108), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n942), .B(new_n977), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n911), .A3(new_n962), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n948), .B1(new_n976), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n975), .A2(new_n962), .A3(new_n911), .ZN(new_n985));
  INV_X1    g560(.A(new_n963), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n964), .A2(new_n981), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n984), .B1(new_n948), .B2(new_n987), .ZN(G397));
  XNOR2_X1  g563(.A(new_n786), .B(new_n788), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT109), .ZN(new_n990));
  INV_X1    g565(.A(G1996), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n817), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n816), .A2(G1996), .ZN(new_n993));
  OR3_X1    g568(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n742), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n739), .B(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n884), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n470), .A2(KEYINPUT66), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n475), .A2(new_n476), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(G40), .A3(new_n465), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n997), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n748), .A3(new_n745), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT124), .B(KEYINPUT48), .Z(new_n1009));
  XNOR2_X1  g584(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n740), .A2(new_n995), .ZN(new_n1011));
  OAI22_X1  g586(.A1(new_n994), .A2(new_n1011), .B1(G2067), .B2(new_n786), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1007), .A2(new_n1010), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1006), .B1(new_n990), .B2(new_n816), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n1014), .B(KEYINPUT123), .Z(new_n1015));
  NAND2_X1  g590(.A1(new_n1006), .A2(new_n991), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT46), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(KEYINPUT47), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT47), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(G8), .B1(new_n999), .B2(new_n1005), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT113), .B(G1981), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n710), .A2(new_n1023), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n515), .A2(G86), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n596), .A2(new_n592), .ZN(new_n1026));
  OAI21_X1  g601(.A(G1981), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1022), .B1(new_n1029), .B2(KEYINPUT49), .ZN(new_n1030));
  AOI211_X1 g605(.A(KEYINPUT114), .B(KEYINPUT49), .C1(new_n1024), .C2(new_n1027), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1030), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G288), .A2(G1976), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1035), .A2(new_n1036), .B1(new_n710), .B2(new_n1023), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G288), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(new_n1022), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1042), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1035), .A2(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1004), .A2(G40), .A3(new_n465), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n884), .A2(KEYINPUT45), .A3(new_n998), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1000), .B1(G164), .B2(G1384), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT110), .B(G1971), .Z(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n999), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1005), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n878), .A2(new_n882), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n998), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n1058));
  NOR2_X1   g633(.A1(G164), .A2(G1384), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(new_n1053), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1054), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1051), .B1(new_n1062), .B2(G2090), .ZN(new_n1063));
  INV_X1    g638(.A(G8), .ZN(new_n1064));
  NOR2_X1   g639(.A1(G166), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1065), .B1(new_n1068), .B2(KEYINPUT55), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1063), .A2(G8), .A3(new_n1070), .ZN(new_n1071));
  OAI22_X1  g646(.A1(new_n1037), .A2(new_n1022), .B1(new_n1045), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1055), .A2(new_n1053), .A3(new_n998), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1046), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1053), .B1(new_n884), .B2(new_n998), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1075), .A2(G2090), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1067), .B(new_n1069), .C1(new_n1078), .C2(new_n1064), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1035), .A2(new_n1079), .A3(new_n1044), .A4(new_n1071), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1001), .B(new_n1046), .C1(new_n1000), .C2(new_n1056), .ZN(new_n1081));
  INV_X1    g656(.A(G1966), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G2084), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1054), .A2(new_n1061), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1064), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G168), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1073), .B1(new_n1080), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1063), .A2(G8), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1070), .A2(KEYINPUT115), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1087), .A2(new_n1073), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n1035), .A3(new_n1044), .A4(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1072), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1083), .A2(new_n1085), .A3(G168), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G8), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(KEYINPUT122), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT51), .B1(new_n1095), .B2(G8), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1101), .A2(new_n1102), .B1(G286), .B2(new_n1086), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT62), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1100), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1049), .A2(G2078), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1108), .A2(new_n1109), .B1(new_n1062), .B2(new_n798), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(G2078), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1110), .B1(new_n1081), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1080), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1105), .A2(new_n1107), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1094), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n824), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT56), .B(G2072), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n583), .A2(KEYINPUT57), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n565), .A2(new_n1123), .A3(new_n567), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n568), .A2(KEYINPUT117), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n578), .A3(new_n582), .A4(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT118), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1128), .A2(KEYINPUT118), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1122), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1121), .A2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n999), .A2(new_n1005), .A3(G2067), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n1062), .B2(new_n827), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(new_n622), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1121), .A2(new_n1132), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1133), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1135), .A2(KEYINPUT60), .A3(new_n622), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n622), .B1(new_n1135), .B2(KEYINPUT60), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1139), .A2(new_n1140), .B1(KEYINPUT60), .B2(new_n1135), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1131), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1129), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(new_n1122), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1133), .A2(new_n1145), .A3(KEYINPUT61), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1046), .A2(new_n1047), .A3(new_n991), .A4(new_n1048), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT58), .B(G1341), .Z(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n999), .B2(new_n1005), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n558), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT119), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(new_n1154), .A3(new_n558), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1147), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1154), .B1(new_n1151), .B2(new_n558), .ZN(new_n1157));
  INV_X1    g732(.A(new_n558), .ZN(new_n1158));
  AOI211_X1 g733(.A(KEYINPUT119), .B(new_n1158), .C1(new_n1148), .C2(new_n1150), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1157), .A2(new_n1159), .A3(KEYINPUT59), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1146), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1144), .B1(new_n1143), .B2(new_n1122), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1137), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(KEYINPUT120), .B(new_n1162), .C1(new_n1137), .C2(new_n1163), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1161), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1141), .B1(new_n1168), .B2(KEYINPUT121), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n1170));
  AOI211_X1 g745(.A(new_n1170), .B(new_n1161), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1138), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(G301), .B(KEYINPUT54), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1113), .A2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n465), .A2(new_n475), .A3(G40), .A4(new_n1111), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1175), .B1(new_n1052), .B2(KEYINPUT45), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1173), .B1(new_n1176), .B2(new_n1001), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1110), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g754(.A(new_n1080), .B(new_n1179), .C1(new_n1100), .C2(new_n1103), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1117), .B1(new_n1172), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n997), .ZN(new_n1182));
  XNOR2_X1  g757(.A(G290), .B(new_n748), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1005), .B(new_n1001), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1021), .B1(new_n1181), .B2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n1187));
  NAND3_X1  g761(.A1(new_n682), .A2(G319), .A3(new_n683), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1188), .A2(KEYINPUT125), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n1190));
  NAND4_X1  g764(.A1(new_n682), .A2(new_n1190), .A3(G319), .A4(new_n683), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g766(.A1(new_n708), .A2(new_n664), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g767(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n912), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g769(.A(new_n1187), .B1(new_n987), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g770(.A(G37), .B1(new_n903), .B2(new_n905), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1193), .B1(new_n1197), .B2(new_n910), .ZN(new_n1198));
  AND2_X1   g772(.A1(new_n985), .A2(new_n986), .ZN(new_n1199));
  AND4_X1   g773(.A1(new_n911), .A2(new_n981), .A3(new_n962), .A4(new_n963), .ZN(new_n1200));
  OAI211_X1 g774(.A(KEYINPUT126), .B(new_n1198), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  AND3_X1   g775(.A1(new_n1196), .A2(KEYINPUT127), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g776(.A(KEYINPUT127), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1203));
  NOR2_X1   g777(.A1(new_n1202), .A2(new_n1203), .ZN(G308));
  NAND2_X1  g778(.A1(new_n1196), .A2(new_n1201), .ZN(G225));
endmodule


