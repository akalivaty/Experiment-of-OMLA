//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  OR2_X1    g004(.A1(new_n190), .A2(KEYINPUT16), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(G146), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n187), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n199), .B(KEYINPUT72), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT24), .B(G110), .Z(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n203));
  INV_X1    g017(.A(new_n198), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n196), .B(new_n203), .C1(new_n204), .C2(KEYINPUT23), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G110), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n192), .B(new_n194), .C1(new_n202), .C2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n192), .A2(KEYINPUT73), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n188), .A2(new_n191), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n193), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT73), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n188), .A2(new_n211), .A3(new_n191), .A4(G146), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n200), .A2(new_n201), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n205), .A2(G110), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n207), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G137), .ZN(new_n218));
  INV_X1    g032(.A(G953), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n219), .A2(G221), .A3(G234), .ZN(new_n220));
  XOR2_X1   g034(.A(new_n218), .B(new_n220), .Z(new_n221));
  XNOR2_X1  g035(.A(new_n217), .B(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G902), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n224), .B(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G217), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(G234), .B2(new_n223), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n222), .B(KEYINPUT74), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n228), .A2(G902), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(G472), .A2(G902), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G143), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT65), .B1(new_n237), .B2(G146), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n193), .A3(G143), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(G146), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n238), .A2(new_n240), .A3(new_n241), .A4(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n193), .A2(G143), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n242), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT64), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT64), .B1(new_n245), .B2(new_n247), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n243), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(G137), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT11), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n256), .B1(new_n253), .B2(G137), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(G131), .ZN(new_n260));
  OAI211_X1 g074(.A(KEYINPUT66), .B(new_n243), .C1(new_n248), .C2(new_n249), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n252), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  XOR2_X1   g076(.A(G116), .B(G119), .Z(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT2), .B(G113), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n237), .A2(G146), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n268));
  OAI21_X1  g082(.A(G128), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n245), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n238), .A2(new_n240), .A3(new_n242), .A4(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n258), .ZN(new_n274));
  OAI21_X1  g088(.A(G131), .B1(new_n274), .B2(new_n254), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n273), .B(new_n275), .C1(G131), .C2(new_n259), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n262), .A2(new_n266), .A3(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(G237), .A2(G953), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G210), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT27), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT26), .B(G101), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n262), .A2(KEYINPUT30), .A3(new_n276), .ZN(new_n284));
  INV_X1    g098(.A(G131), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n259), .B(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n276), .B1(new_n286), .B2(new_n250), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n284), .A2(new_n265), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT67), .B1(new_n291), .B2(KEYINPUT31), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT67), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT31), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n293), .B(new_n294), .C1(new_n283), .C2(new_n290), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n277), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n287), .A2(new_n265), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n262), .A2(KEYINPUT28), .A3(new_n266), .A4(new_n276), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n282), .B(KEYINPUT68), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n283), .A2(new_n294), .A3(new_n290), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT69), .B1(new_n296), .B2(new_n305), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n284), .A2(new_n265), .A3(new_n289), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n277), .A2(new_n282), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT31), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n293), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n291), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT69), .ZN(new_n313));
  INV_X1    g127(.A(new_n305), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n236), .B1(new_n306), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n298), .ZN(new_n317));
  OR2_X1    g131(.A1(new_n277), .A2(KEYINPUT71), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n277), .A2(KEYINPUT71), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n262), .A2(new_n276), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n318), .B(new_n319), .C1(new_n266), .C2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n317), .B1(new_n321), .B2(KEYINPUT28), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(KEYINPUT29), .A3(new_n282), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n290), .A2(new_n277), .ZN(new_n324));
  INV_X1    g138(.A(new_n282), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(new_n327), .C1(new_n301), .C2(new_n302), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n223), .A3(new_n328), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n316), .A2(KEYINPUT32), .B1(G472), .B2(new_n329), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n296), .A2(KEYINPUT69), .A3(new_n305), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n313), .B1(new_n312), .B2(new_n314), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n235), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n234), .B1(new_n330), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G469), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n238), .A2(new_n240), .A3(new_n242), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n340), .A2(new_n269), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n272), .A2(KEYINPUT75), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G107), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(G104), .ZN(new_n345));
  INV_X1    g159(.A(G104), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G107), .ZN(new_n347));
  OAI21_X1  g161(.A(G101), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT3), .B1(new_n346), .B2(G107), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n344), .A3(G104), .ZN(new_n351));
  INV_X1    g165(.A(G101), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n346), .A2(G107), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n349), .A2(new_n351), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n348), .B(new_n354), .C1(new_n272), .C2(KEYINPUT75), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT76), .B1(new_n343), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n355), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n340), .A2(new_n269), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(KEYINPUT75), .A3(new_n272), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n273), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n354), .A2(new_n348), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n356), .A2(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT12), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n364), .A2(new_n365), .A3(new_n286), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(new_n363), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n343), .A2(KEYINPUT76), .A3(new_n355), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n358), .B1(new_n357), .B2(new_n360), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT12), .B1(new_n370), .B2(new_n260), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n339), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n368), .B2(new_n369), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G101), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT4), .A3(new_n354), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n378), .A3(G101), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n252), .A3(new_n261), .ZN(new_n381));
  INV_X1    g195(.A(new_n363), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n273), .A3(KEYINPUT10), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n374), .A2(new_n286), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(G110), .B(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n219), .A2(G227), .ZN(new_n386));
  XOR2_X1   g200(.A(new_n385), .B(new_n386), .Z(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n365), .B1(new_n364), .B2(new_n286), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n370), .A2(KEYINPUT12), .A3(new_n260), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT79), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n372), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n381), .A2(new_n383), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT10), .B1(new_n356), .B2(new_n361), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT78), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT78), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n374), .A2(new_n397), .A3(new_n381), .A4(new_n383), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n398), .A3(new_n260), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n388), .B1(new_n399), .B2(new_n384), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n393), .B1(new_n400), .B2(KEYINPUT80), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT80), .ZN(new_n402));
  AOI211_X1 g216(.A(new_n402), .B(new_n388), .C1(new_n399), .C2(new_n384), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n338), .B(new_n223), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(G469), .A2(G902), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n390), .A2(new_n391), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT77), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n406), .A2(new_n407), .A3(new_n384), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n406), .B2(new_n384), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n387), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n389), .A2(new_n399), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(G469), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n404), .A2(new_n405), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT9), .B(G234), .ZN(new_n414));
  OAI21_X1  g228(.A(G221), .B1(new_n414), .B2(G902), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G214), .B1(G237), .B2(G902), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G210), .B1(G237), .B2(G902), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT85), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n219), .A2(G224), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT7), .ZN(new_n423));
  INV_X1    g237(.A(G125), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n362), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n425), .B2(KEYINPUT83), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n250), .A2(G125), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n427), .A2(new_n425), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n426), .B1(new_n428), .B2(KEYINPUT83), .ZN(new_n429));
  XNOR2_X1  g243(.A(G110), .B(G122), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT8), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n263), .A2(new_n264), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT5), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n195), .A3(G116), .ZN(new_n434));
  OAI211_X1 g248(.A(G113), .B(new_n434), .C1(new_n263), .C2(new_n433), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n382), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n382), .B1(new_n432), .B2(new_n435), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n431), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT7), .B1(new_n422), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(new_n440), .B2(new_n422), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n427), .A2(new_n425), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n429), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n265), .A2(new_n377), .A3(new_n379), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT81), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT81), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n265), .A2(new_n377), .A3(new_n448), .A4(new_n379), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n447), .A2(new_n430), .A3(new_n436), .A4(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(G902), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n436), .A3(new_n449), .ZN(new_n452));
  INV_X1    g266(.A(new_n430), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT6), .A3(new_n450), .ZN(new_n455));
  XOR2_X1   g269(.A(new_n422), .B(KEYINPUT82), .Z(new_n456));
  XNOR2_X1  g270(.A(new_n428), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n458), .A3(new_n453), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n421), .B1(new_n451), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n451), .A2(new_n460), .A3(new_n421), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n418), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(G143), .B1(new_n278), .B2(G214), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n278), .A2(G143), .A3(G214), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT17), .A3(G131), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT88), .ZN(new_n471));
  INV_X1    g285(.A(new_n468), .ZN(new_n472));
  OAI21_X1  g286(.A(G131), .B1(new_n472), .B2(new_n466), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n467), .A2(new_n285), .A3(new_n468), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n471), .B1(new_n475), .B2(KEYINPUT17), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT17), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT88), .A4(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n213), .A2(new_n470), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G113), .B(G122), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(new_n346), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n469), .A2(KEYINPUT18), .A3(G131), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n424), .A2(G140), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n190), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G146), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n194), .ZN(new_n486));
  NAND2_X1  g300(.A1(KEYINPUT18), .A2(G131), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n467), .A2(new_n468), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n482), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n479), .A2(new_n481), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n481), .B1(new_n479), .B2(new_n489), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n223), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G475), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT87), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n190), .A2(new_n483), .A3(KEYINPUT19), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT19), .B1(new_n190), .B2(new_n483), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n193), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n192), .A3(KEYINPUT86), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n475), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT86), .B1(new_n498), .B2(new_n192), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n495), .B(new_n489), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n481), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n501), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(new_n475), .A3(new_n499), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n495), .B1(new_n506), .B2(new_n489), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n490), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT20), .ZN(new_n509));
  NOR2_X1   g323(.A1(G475), .A2(G902), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n494), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT89), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT89), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n494), .B(new_n515), .C1(new_n511), .C2(new_n512), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n219), .A2(G952), .ZN(new_n518));
  NAND2_X1  g332(.A1(G234), .A2(G237), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT21), .B(G898), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n519), .A2(G902), .A3(G953), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G478), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(KEYINPUT15), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n527));
  INV_X1    g341(.A(G122), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n527), .B1(new_n528), .B2(G116), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n530));
  INV_X1    g344(.A(G116), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT90), .A3(G122), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n528), .A2(G116), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n529), .A2(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT14), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT93), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT93), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n539), .A3(KEYINPUT14), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n535), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT94), .B1(new_n541), .B2(new_n344), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT94), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n539), .B1(new_n536), .B2(KEYINPUT14), .ZN(new_n544));
  AOI211_X1 g358(.A(KEYINPUT93), .B(new_n530), .C1(new_n529), .C2(new_n532), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n543), .B(G107), .C1(new_n546), .C2(new_n535), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n197), .B2(G143), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n237), .A2(KEYINPUT91), .A3(G128), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(G128), .B2(new_n237), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n553), .A2(G134), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(G134), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n536), .A2(new_n534), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n554), .A2(new_n555), .B1(G107), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n548), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n550), .A2(new_n551), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(KEYINPUT13), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n237), .A2(G128), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT92), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT92), .ZN(new_n564));
  OAI221_X1 g378(.A(new_n564), .B1(G128), .B2(new_n237), .C1(new_n560), .C2(KEYINPUT13), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n560), .A2(KEYINPUT13), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G134), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n553), .A2(G134), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n556), .A2(G107), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n344), .B1(new_n536), .B2(new_n534), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n414), .A2(new_n227), .A3(G953), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT95), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n559), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n575), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n557), .B1(new_n542), .B2(new_n547), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n569), .B1(new_n571), .B2(new_n570), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n567), .B2(G134), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n577), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n576), .A2(new_n581), .A3(new_n582), .A4(new_n223), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n526), .B1(new_n583), .B2(KEYINPUT96), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(KEYINPUT96), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n576), .A2(new_n581), .A3(new_n586), .A4(new_n223), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n584), .B1(new_n588), .B2(new_n526), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n517), .A2(new_n524), .A3(new_n589), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n416), .A2(new_n465), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n337), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n306), .B2(new_n315), .ZN(new_n595));
  INV_X1    g409(.A(G472), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n233), .B(new_n333), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n594), .B1(new_n597), .B2(new_n416), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n223), .B1(new_n331), .B2(new_n332), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n316), .B1(new_n599), .B2(G472), .ZN(new_n600));
  INV_X1    g414(.A(new_n415), .ZN(new_n601));
  INV_X1    g415(.A(new_n411), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n384), .B1(new_n366), .B2(new_n371), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT77), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n406), .A2(new_n407), .A3(new_n384), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n602), .B1(new_n606), .B2(new_n387), .ZN(new_n607));
  OAI21_X1  g421(.A(G469), .B1(new_n607), .B2(G902), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n601), .B1(new_n608), .B2(new_n404), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n600), .A2(KEYINPUT98), .A3(new_n233), .A4(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n598), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n517), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n576), .A2(new_n581), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n525), .A2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n576), .A2(new_n581), .A3(new_n223), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n525), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n618), .A2(KEYINPUT99), .A3(new_n525), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n612), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n464), .A2(new_n524), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n611), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NOR3_X1   g444(.A1(new_n626), .A2(new_n513), .A3(new_n589), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n611), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  INV_X1    g448(.A(new_n221), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n217), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n231), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n229), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n333), .B(new_n639), .C1(new_n595), .C2(new_n596), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n591), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  OAI211_X1 g458(.A(KEYINPUT32), .B(new_n235), .C1(new_n331), .C2(new_n332), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n329), .A2(G472), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n306), .A2(new_n315), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n334), .B1(new_n648), .B2(new_n235), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n639), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n523), .A2(G900), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n520), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n494), .B(new_n652), .C1(new_n511), .C2(new_n512), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n589), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n609), .A2(new_n464), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT100), .B1(new_n650), .B2(new_n655), .ZN(new_n656));
  AND4_X1   g470(.A1(new_n415), .A2(new_n413), .A3(new_n464), .A4(new_n654), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n645), .B(new_n646), .C1(new_n316), .C2(new_n334), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n657), .A2(new_n658), .A3(new_n659), .A4(new_n639), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  NOR4_X1   g476(.A1(new_n639), .A2(new_n517), .A3(new_n418), .A4(new_n589), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT101), .ZN(new_n664));
  INV_X1    g478(.A(new_n291), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n321), .B2(new_n302), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n666), .B2(G902), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n336), .A2(new_n645), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n462), .A2(new_n463), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT38), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n652), .B(KEYINPUT39), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n609), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n664), .A2(new_n673), .A3(new_n676), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  AOI22_X1  g493(.A1(new_n330), .A2(new_n336), .B1(new_n229), .B2(new_n638), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n416), .A2(new_n465), .ZN(new_n681));
  INV_X1    g495(.A(new_n652), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n625), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  OAI21_X1  g499(.A(new_n223), .B1(new_n401), .B2(new_n403), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(G469), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n687), .A2(new_n415), .A3(new_n404), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n659), .A2(new_n627), .A3(new_n233), .A4(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n337), .A2(KEYINPUT102), .A3(new_n627), .A4(new_n688), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT41), .B(G113), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT103), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n693), .B(new_n695), .ZN(G15));
  NAND4_X1  g510(.A1(new_n659), .A2(new_n233), .A3(new_n631), .A4(new_n688), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  AND4_X1   g512(.A1(new_n415), .A2(new_n687), .A3(new_n404), .A4(new_n464), .ZN(new_n699));
  INV_X1    g513(.A(new_n590), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n659), .A2(new_n699), .A3(new_n700), .A4(new_n639), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  OAI21_X1  g516(.A(KEYINPUT105), .B1(new_n517), .B2(new_n589), .ZN(new_n703));
  INV_X1    g517(.A(new_n589), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(new_n705), .A3(new_n514), .A4(new_n516), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n626), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n688), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n302), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n322), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n309), .A2(new_n304), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n236), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n595), .B2(new_n596), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n599), .A2(KEYINPUT104), .A3(G472), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n709), .A2(KEYINPUT106), .A3(new_n233), .A4(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n719));
  INV_X1    g533(.A(new_n713), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT104), .B1(new_n599), .B2(G472), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n595), .A2(new_n714), .A3(new_n596), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n233), .B(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n719), .B1(new_n723), .B2(new_n708), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NAND4_X1  g540(.A1(new_n717), .A2(new_n639), .A3(new_n683), .A4(new_n699), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT107), .B(G125), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G27));
  NOR2_X1   g543(.A1(new_n601), .A2(new_n418), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n462), .A2(new_n463), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n413), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n413), .A2(KEYINPUT108), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(new_n316), .B2(KEYINPUT32), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT32), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n333), .A2(KEYINPUT109), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n330), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n737), .A2(new_n233), .A3(new_n683), .A4(new_n742), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n734), .B(new_n731), .C1(new_n608), .C2(new_n404), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT108), .B1(new_n413), .B2(new_n732), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n233), .B1(new_n647), .B2(new_n649), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n683), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(KEYINPUT42), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n743), .A2(KEYINPUT42), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  NAND3_X1  g566(.A1(new_n737), .A2(new_n337), .A3(new_n654), .ZN(new_n753));
  XOR2_X1   g567(.A(KEYINPUT110), .B(G134), .Z(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G36));
  NAND2_X1  g569(.A1(new_n517), .A2(new_n624), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT43), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n333), .B1(new_n595), .B2(new_n596), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n639), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n404), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n410), .A2(new_n411), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n607), .A2(KEYINPUT45), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n767), .A3(G469), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n405), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT46), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n763), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(KEYINPUT46), .A3(new_n405), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n601), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n674), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n451), .A2(new_n460), .A3(new_n421), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n775), .A2(new_n461), .A3(new_n418), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n760), .B2(new_n761), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n762), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  XNOR2_X1  g594(.A(new_n773), .B(KEYINPUT47), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n749), .A2(new_n659), .A3(new_n233), .A4(new_n777), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  NOR2_X1   g598(.A1(new_n757), .A2(new_n520), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n688), .A2(new_n776), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n233), .A3(new_n742), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT48), .ZN(new_n789));
  INV_X1    g603(.A(new_n699), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n785), .A2(new_n233), .A3(new_n717), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n789), .B(new_n518), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n625), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n234), .A2(new_n520), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n669), .A2(new_n786), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT117), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n792), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  OR2_X1    g611(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n672), .A2(new_n688), .A3(new_n418), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n612), .A2(new_n624), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n802), .B1(new_n796), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n791), .A2(new_n777), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n687), .A2(new_n404), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(new_n601), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n805), .B1(new_n781), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n717), .A2(new_n639), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n800), .A2(new_n801), .B1(new_n810), .B2(new_n787), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n804), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n797), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n416), .A2(new_n639), .A3(new_n682), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n703), .A2(new_n706), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n464), .A3(new_n668), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n661), .A2(new_n684), .A3(new_n727), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n727), .A2(new_n684), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n823), .A2(KEYINPUT52), .A3(new_n661), .A4(new_n819), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n737), .A2(new_n717), .A3(new_n639), .A4(new_n683), .ZN(new_n826));
  INV_X1    g640(.A(new_n653), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n776), .A2(new_n827), .A3(new_n589), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n828), .A2(new_n413), .A3(new_n415), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT113), .B1(new_n680), .B2(new_n829), .ZN(new_n830));
  AND4_X1   g644(.A1(KEYINPUT113), .A2(new_n829), .A3(new_n659), .A4(new_n639), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n826), .B(new_n753), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n517), .A2(new_n589), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n517), .B2(new_n624), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n626), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n598), .A2(new_n610), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n591), .B1(new_n337), .B2(new_n641), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n701), .A2(new_n697), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n691), .B2(new_n692), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(new_n725), .A3(new_n751), .A4(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n825), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n841), .A2(new_n751), .A3(new_n725), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n836), .A2(new_n837), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT113), .ZN(new_n847));
  INV_X1    g661(.A(new_n829), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n848), .B2(new_n650), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n680), .A2(KEYINPUT113), .A3(new_n829), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n846), .A2(new_n753), .A3(new_n826), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n822), .A2(new_n824), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT53), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT54), .B1(new_n844), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n843), .B1(new_n825), .B2(new_n842), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  AND4_X1   g672(.A1(KEYINPUT53), .A2(new_n841), .A3(new_n751), .A4(new_n725), .ZN(new_n859));
  OR3_X1    g673(.A1(new_n832), .A2(KEYINPUT115), .A3(new_n838), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT115), .B1(new_n832), .B2(new_n838), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n854), .A2(new_n859), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n857), .A2(new_n858), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  OAI22_X1  g678(.A1(new_n816), .A2(new_n864), .B1(G952), .B2(G953), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT49), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n806), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT112), .Z(new_n868));
  NAND2_X1  g682(.A1(new_n233), .A2(new_n730), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT111), .Z(new_n870));
  NOR3_X1   g684(.A1(new_n870), .A2(new_n671), .A3(new_n756), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n871), .B(new_n669), .C1(new_n866), .C2(new_n806), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n865), .B1(new_n868), .B2(new_n872), .ZN(G75));
  AND4_X1   g687(.A1(new_n854), .A2(new_n859), .A3(new_n860), .A4(new_n861), .ZN(new_n874));
  INV_X1    g688(.A(new_n843), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n853), .B2(new_n854), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n223), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n420), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT56), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n455), .A2(new_n459), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n457), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT55), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n879), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n883), .B1(new_n879), .B2(new_n880), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n219), .A2(G952), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G51));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n877), .A2(new_n223), .A3(new_n768), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n405), .B(KEYINPUT57), .Z(new_n890));
  NOR3_X1   g704(.A1(new_n874), .A2(new_n876), .A3(KEYINPUT54), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n858), .B1(new_n857), .B2(new_n862), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n401), .A2(new_n403), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n889), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n888), .B1(new_n896), .B2(new_n886), .ZN(new_n897));
  INV_X1    g711(.A(new_n886), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT54), .B1(new_n874), .B2(new_n876), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n863), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n894), .B1(new_n900), .B2(new_n890), .ZN(new_n901));
  OAI211_X1 g715(.A(KEYINPUT118), .B(new_n898), .C1(new_n901), .C2(new_n889), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n897), .A2(new_n902), .ZN(G54));
  NAND3_X1  g717(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .ZN(new_n904));
  INV_X1    g718(.A(new_n508), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n886), .ZN(G60));
  INV_X1    g722(.A(new_n615), .ZN(new_n909));
  NAND2_X1  g723(.A1(G478), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT59), .Z(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n900), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n898), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n911), .B1(new_n856), .B2(new_n863), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n615), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT119), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n886), .B1(new_n900), .B2(new_n912), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT119), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n918), .B(new_n919), .C1(new_n615), .C2(new_n915), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n920), .ZN(G63));
  NAND2_X1  g735(.A1(new_n857), .A2(new_n862), .ZN(new_n922));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n230), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT121), .B1(new_n926), .B2(new_n886), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n924), .B1(new_n857), .B2(new_n862), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n928), .B(new_n898), .C1(new_n929), .C2(new_n230), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n637), .B(new_n925), .C1(new_n874), .C2(new_n876), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT120), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n922), .A2(new_n933), .A3(new_n637), .A4(new_n925), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n927), .A2(new_n930), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n926), .A2(KEYINPUT122), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n926), .A2(KEYINPUT122), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n886), .A2(new_n937), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n939), .A2(new_n935), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n938), .A2(new_n942), .ZN(G66));
  NAND3_X1  g757(.A1(new_n841), .A2(new_n725), .A3(new_n846), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n219), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT123), .Z(new_n946));
  INV_X1    g760(.A(G224), .ZN(new_n947));
  OAI21_X1  g761(.A(G953), .B1(new_n521), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT124), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n881), .B1(G898), .B2(new_n219), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G69));
  AND2_X1   g766(.A1(new_n742), .A2(new_n233), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n774), .A2(new_n464), .A3(new_n818), .A4(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n783), .A2(new_n751), .A3(new_n753), .A4(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n779), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n823), .A2(new_n661), .ZN(new_n957));
  OR3_X1    g771(.A1(new_n956), .A2(KEYINPUT125), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(KEYINPUT125), .B1(new_n956), .B2(new_n957), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n219), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n284), .A2(new_n289), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n496), .A2(new_n497), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(G900), .B2(G953), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n957), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n678), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(KEYINPUT62), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n968), .A2(new_n971), .A3(new_n678), .ZN(new_n972));
  NOR4_X1   g786(.A1(new_n747), .A2(new_n675), .A3(new_n834), .A4(new_n777), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n956), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n970), .A2(new_n783), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n964), .B1(new_n975), .B2(new_n219), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n967), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n219), .B1(G227), .B2(G900), .ZN(new_n980));
  INV_X1    g794(.A(new_n966), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n960), .B2(new_n219), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT126), .B1(new_n982), .B2(new_n976), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n979), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n980), .B1(new_n979), .B2(new_n983), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(G72));
  XNOR2_X1  g800(.A(new_n324), .B(KEYINPUT127), .ZN(new_n987));
  INV_X1    g801(.A(new_n944), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n960), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  AOI211_X1 g805(.A(new_n282), .B(new_n987), .C1(new_n989), .C2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n987), .A2(new_n282), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n975), .A2(new_n944), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(new_n994), .B2(new_n991), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n844), .A2(new_n855), .ZN(new_n996));
  INV_X1    g810(.A(new_n326), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n991), .B1(new_n997), .B2(new_n665), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n898), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n992), .A2(new_n995), .A3(new_n999), .ZN(G57));
endmodule


