//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944;
  XOR2_X1   g000(.A(G134gat), .B(G162gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT93), .ZN(new_n203));
  AND2_X1   g002(.A1(G232gat), .A2(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(KEYINPUT41), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n203), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G190gat), .B(G218gat), .Z(new_n207));
  NAND2_X1  g006(.A1(G43gat), .A2(G50gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G43gat), .A2(G50gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT15), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT85), .B(G43gat), .ZN(new_n212));
  INV_X1    g011(.A(G50gat), .ZN(new_n213));
  AOI211_X1 g012(.A(KEYINPUT15), .B(new_n209), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n215), .A2(KEYINPUT14), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(KEYINPUT14), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT84), .B(G36gat), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n216), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n211), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n220), .A2(new_n211), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226));
  INV_X1    g025(.A(G85gat), .ZN(new_n227));
  INV_X1    g026(.A(G92gat), .ZN(new_n228));
  AOI22_X1  g027(.A1(KEYINPUT8), .A2(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(new_n227), .B2(new_n228), .ZN(new_n231));
  NAND4_X1  g030(.A1(KEYINPUT94), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(G99gat), .B(G106gat), .Z(new_n234));
  OR2_X1    g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n237), .B(KEYINPUT95), .Z(new_n238));
  NAND2_X1  g037(.A1(new_n225), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n223), .ZN(new_n240));
  INV_X1    g039(.A(new_n237), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n240), .A2(new_n241), .B1(KEYINPUT41), .B2(new_n204), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n207), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n206), .B1(new_n243), .B2(KEYINPUT96), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT97), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n239), .A2(new_n207), .A3(new_n242), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(new_n243), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT97), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n248), .B(new_n206), .C1(new_n243), .C2(KEYINPUT96), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n245), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n247), .B1(new_n245), .B2(new_n249), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(G57gat), .B(G64gat), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT9), .ZN(new_n254));
  OR2_X1    g053(.A1(G71gat), .A2(G78gat), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n255), .A2(KEYINPUT90), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(KEYINPUT90), .ZN(new_n257));
  NAND2_X1  g056(.A1(G71gat), .A2(G78gat), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n254), .A2(new_n256), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n253), .A2(KEYINPUT91), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT9), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G57gat), .B(G64gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT91), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT21), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G231gat), .A2(G233gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(G127gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(G15gat), .B(G22gat), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n273), .A2(G1gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT16), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n275), .B2(G1gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(KEYINPUT86), .A2(G8gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(KEYINPUT86), .A2(G8gat), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT86), .ZN(new_n281));
  INV_X1    g080(.A(G8gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n268), .B2(new_n267), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n272), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT92), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(G155gat), .ZN(new_n289));
  XOR2_X1   g088(.A(G183gat), .B(G211gat), .Z(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n286), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n252), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT99), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT98), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n236), .B(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n235), .A2(new_n259), .A3(new_n266), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n235), .A2(new_n259), .A3(new_n266), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n236), .A2(new_n296), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT98), .B1(new_n233), .B2(new_n234), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n303), .A3(KEYINPUT99), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n299), .A2(new_n304), .B1(new_n267), .B2(new_n237), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G230gat), .A2(G233gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(G120gat), .B(G148gat), .Z(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT100), .ZN(new_n311));
  XNOR2_X1  g110(.A(G176gat), .B(G204gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n311), .B(new_n312), .Z(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT10), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n237), .A2(new_n267), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(new_n305), .B2(new_n316), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(new_n308), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n307), .B(KEYINPUT101), .Z(new_n321));
  OAI21_X1  g120(.A(new_n309), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n320), .B1(new_n322), .B2(new_n313), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n294), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325));
  XNOR2_X1  g124(.A(G155gat), .B(G162gat), .ZN(new_n326));
  INV_X1    g125(.A(G141gat), .ZN(new_n327));
  INV_X1    g126(.A(G148gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G162gat), .ZN(new_n332));
  INV_X1    g131(.A(G155gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT73), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G155gat), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n332), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT2), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n326), .B(new_n331), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n329), .A2(new_n338), .A3(new_n330), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n332), .A2(G155gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n333), .A2(G162gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n325), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G113gat), .B(G120gat), .ZN(new_n346));
  INV_X1    g145(.A(G127gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(G134gat), .ZN(new_n348));
  INV_X1    g147(.A(G134gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(G127gat), .ZN(new_n350));
  OAI22_X1  g149(.A1(new_n346), .A2(KEYINPUT1), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G120gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G113gat), .ZN(new_n353));
  INV_X1    g152(.A(G113gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G120gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G127gat), .B(G134gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n351), .A2(new_n359), .A3(KEYINPUT74), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT74), .B1(new_n351), .B2(new_n359), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n345), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n334), .A2(new_n336), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n338), .B1(new_n363), .B2(G162gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n326), .A2(new_n329), .A3(new_n330), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n325), .B(new_n344), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n339), .A2(KEYINPUT75), .A3(new_n325), .A4(new_n344), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n344), .B1(new_n364), .B2(new_n365), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n351), .A2(new_n359), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n351), .A2(new_n359), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT73), .B(G155gat), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT2), .B1(new_n378), .B2(new_n332), .ZN(new_n379));
  AND4_X1   g178(.A1(new_n341), .A2(new_n329), .A3(new_n342), .A4(new_n330), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n379), .A2(new_n380), .B1(new_n343), .B2(new_n340), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n377), .A2(new_n381), .A3(KEYINPUT4), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n371), .A2(new_n372), .A3(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n385));
  INV_X1    g184(.A(new_n361), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n351), .A2(new_n359), .A3(KEYINPUT74), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n374), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n377), .A2(new_n381), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n372), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n385), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT0), .ZN(new_n395));
  XNOR2_X1  g194(.A(G57gat), .B(G85gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  NAND4_X1  g196(.A1(new_n371), .A2(new_n372), .A3(new_n383), .A4(new_n385), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n393), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n397), .B1(new_n393), .B2(new_n398), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT77), .B1(new_n402), .B2(KEYINPUT6), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(KEYINPUT77), .A3(KEYINPUT6), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT27), .B(G183gat), .ZN(new_n409));
  INV_X1    g208(.A(G190gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n411));
  AND2_X1   g210(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n409), .B(new_n410), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G183gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT27), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G183gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n417), .A3(new_n410), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n412), .A2(new_n411), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(G169gat), .B2(G176gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(G169gat), .A2(G176gat), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n423), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n413), .A2(new_n420), .A3(new_n422), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G169gat), .A2(G176gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(G183gat), .A2(G190gat), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(KEYINPUT24), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT23), .ZN(new_n430));
  INV_X1    g229(.A(G169gat), .ZN(new_n431));
  INV_X1    g230(.A(G176gat), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n428), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n414), .A2(new_n410), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(KEYINPUT24), .A3(new_n427), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT25), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n428), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n433), .A2(new_n429), .ZN(new_n439));
  AND4_X1   g238(.A1(KEYINPUT25), .A2(new_n438), .A3(new_n439), .A4(new_n436), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n425), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n442), .B(KEYINPUT72), .Z(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n438), .A2(new_n439), .A3(new_n436), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT25), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n438), .A2(new_n439), .A3(new_n436), .A4(KEYINPUT25), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT29), .B1(new_n449), .B2(new_n425), .ZN(new_n450));
  INV_X1    g249(.A(new_n442), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n444), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G197gat), .B(G204gat), .ZN(new_n453));
  INV_X1    g252(.A(G211gat), .ZN(new_n454));
  INV_X1    g253(.A(G218gat), .ZN(new_n455));
  OAI22_X1  g254(.A1(new_n454), .A2(new_n455), .B1(KEYINPUT71), .B2(KEYINPUT22), .ZN(new_n456));
  AND2_X1   g255(.A1(KEYINPUT71), .A2(KEYINPUT22), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G211gat), .B(G218gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n452), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n460), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n441), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n443), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n441), .A2(new_n451), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G8gat), .B(G36gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(G64gat), .B(G92gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n472), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n461), .B2(new_n468), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n475), .A3(KEYINPUT30), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT30), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n469), .A2(new_n477), .A3(new_n472), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n408), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT3), .B1(new_n462), .B2(new_n463), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT29), .B1(new_n368), .B2(new_n369), .ZN(new_n482));
  OAI22_X1  g281(.A1(new_n481), .A2(new_n381), .B1(new_n462), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G228gat), .A2(G233gat), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n484), .B(G22gat), .Z(new_n485));
  OR2_X1    g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  XOR2_X1   g285(.A(G78gat), .B(G106gat), .Z(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT31), .B(G50gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT78), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n483), .A2(new_n485), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n486), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n489), .B(KEYINPUT78), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n486), .B2(new_n492), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT69), .ZN(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT66), .B(G71gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(G99gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G43gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G227gat), .A2(G233gat), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n503), .B(KEYINPUT64), .Z(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n441), .A2(new_n375), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n377), .B(new_n425), .C1(new_n437), .C2(new_n440), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n502), .B1(new_n508), .B2(KEYINPUT33), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT32), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n507), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n377), .B1(new_n449), .B2(new_n425), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n504), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT33), .ZN(new_n516));
  INV_X1    g315(.A(new_n502), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n515), .B(KEYINPUT32), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n498), .B1(new_n512), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT67), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n505), .A3(new_n507), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(KEYINPUT34), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n521), .A3(KEYINPUT34), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT34), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n506), .A2(new_n526), .A3(new_n505), .A4(new_n507), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n527), .A2(KEYINPUT68), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(KEYINPUT68), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n524), .A2(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n520), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n525), .ZN(new_n532));
  INV_X1    g331(.A(new_n529), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n527), .A2(KEYINPUT68), .ZN(new_n534));
  OAI22_X1  g333(.A1(new_n523), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n515), .A2(KEYINPUT32), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n515), .A2(new_n516), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(new_n502), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n518), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n535), .A2(new_n539), .A3(new_n498), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n497), .A2(new_n531), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT35), .B1(new_n480), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n479), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n543), .A2(KEYINPUT35), .ZN(new_n544));
  INV_X1    g343(.A(new_n497), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n535), .A2(new_n539), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n524), .A2(new_n525), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n528), .A2(new_n529), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n547), .A2(new_n548), .A3(new_n538), .A4(new_n518), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n393), .A2(new_n398), .ZN(new_n552));
  INV_X1    g351(.A(new_n397), .ZN(new_n553));
  AND4_X1   g352(.A1(KEYINPUT77), .A2(new_n552), .A3(KEYINPUT6), .A4(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(new_n405), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT80), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n393), .A2(KEYINPUT80), .A3(new_n398), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n553), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n401), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n551), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n542), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n371), .A2(new_n383), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n391), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n388), .A2(new_n372), .A3(new_n389), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(KEYINPUT39), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT39), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n568), .A3(new_n391), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n397), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT40), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n570), .A2(KEYINPUT79), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT79), .B1(new_n570), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n567), .A2(KEYINPUT40), .A3(new_n397), .A4(new_n569), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n559), .A2(new_n476), .A3(new_n478), .A4(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n497), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n474), .A2(KEYINPUT37), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n475), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT37), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(new_n469), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT38), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT38), .B1(new_n475), .B2(new_n578), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n466), .A2(new_n462), .A3(new_n467), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT81), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n452), .A2(new_n460), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT81), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n466), .A2(new_n588), .A3(new_n462), .A4(new_n467), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT37), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n584), .A2(new_n591), .B1(new_n472), .B2(new_n469), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n555), .A2(new_n560), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n583), .B1(new_n593), .B2(KEYINPUT82), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT82), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n555), .A2(new_n560), .A3(new_n592), .A4(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n577), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n480), .A2(new_n545), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n535), .A2(new_n539), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n547), .A2(new_n548), .B1(new_n538), .B2(new_n518), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT70), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n531), .A2(KEYINPUT36), .A3(new_n540), .ZN(new_n605));
  OAI211_X1 g404(.A(KEYINPUT70), .B(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n563), .B1(new_n597), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n284), .A2(new_n223), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n284), .A2(KEYINPUT87), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT87), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n280), .A2(new_n612), .A3(new_n283), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n610), .B1(new_n614), .B2(new_n225), .ZN(new_n615));
  NAND2_X1  g414(.A1(G229gat), .A2(G233gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(KEYINPUT18), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT88), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n284), .B(new_n223), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n616), .B(KEYINPUT13), .Z(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G113gat), .B(G141gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G197gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT11), .B(G169gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n617), .A2(new_n621), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT18), .B1(new_n615), .B2(new_n616), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n622), .B(new_n629), .C1(new_n631), .C2(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n609), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT89), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n609), .A2(KEYINPUT89), .A3(new_n636), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n324), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n408), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(G1gat), .Z(G1324gat));
  XOR2_X1   g443(.A(KEYINPUT16), .B(G8gat), .Z(new_n645));
  NAND3_X1  g444(.A1(new_n641), .A2(new_n543), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(KEYINPUT102), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n648), .A2(KEYINPUT102), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n282), .B1(new_n641), .B2(new_n543), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n646), .B1(new_n651), .B2(new_n647), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n650), .B2(new_n652), .ZN(G1325gat));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n606), .A2(new_n605), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT70), .B1(new_n550), .B2(new_n599), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n604), .A2(KEYINPUT103), .A3(new_n605), .A4(new_n606), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(G15gat), .B1(new_n642), .B2(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n550), .A2(G15gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n642), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT104), .ZN(G1326gat));
  NAND2_X1  g463(.A1(new_n641), .A2(new_n545), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT105), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT43), .B(G22gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  NOR2_X1   g467(.A1(new_n252), .A2(new_n292), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n323), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT106), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n639), .B2(new_n640), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n408), .A2(G29gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(KEYINPUT107), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(KEYINPUT107), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(KEYINPUT45), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n678));
  INV_X1    g477(.A(new_n252), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n609), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n678), .B1(new_n680), .B2(KEYINPUT44), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  AOI211_X1 g481(.A(KEYINPUT108), .B(new_n682), .C1(new_n609), .C2(new_n679), .ZN(new_n683));
  INV_X1    g482(.A(new_n563), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n657), .A2(new_n598), .A3(new_n658), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT109), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n593), .A2(KEYINPUT82), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n596), .A3(new_n582), .ZN(new_n688));
  INV_X1    g487(.A(new_n577), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n685), .A2(new_n686), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n657), .A2(new_n598), .A3(new_n658), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT109), .B1(new_n692), .B2(new_n597), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n684), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n682), .ZN(new_n695));
  OAI22_X1  g494(.A1(new_n681), .A2(new_n683), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n636), .ZN(new_n697));
  INV_X1    g496(.A(new_n323), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n697), .A2(new_n292), .A3(new_n698), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n408), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n677), .B1(new_n702), .B2(new_n219), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT45), .B1(new_n675), .B2(new_n676), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n703), .A2(new_n704), .ZN(G1328gat));
  NAND3_X1  g504(.A1(new_n672), .A2(new_n543), .A3(new_n218), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT46), .Z(new_n707));
  AND2_X1   g506(.A1(new_n700), .A2(new_n543), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n218), .B2(new_n708), .ZN(G1329gat));
  INV_X1    g508(.A(new_n212), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n700), .A2(new_n710), .A3(new_n659), .ZN(new_n711));
  INV_X1    g510(.A(new_n550), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n710), .B1(new_n672), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(KEYINPUT47), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n714), .A2(KEYINPUT47), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT111), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n716), .B(new_n718), .ZN(G1330gat));
  AOI21_X1  g518(.A(new_n213), .B1(new_n700), .B2(new_n545), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n497), .A2(G50gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT112), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n672), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g524(.A1(new_n636), .A2(new_n323), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n694), .A2(new_n293), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n408), .B(KEYINPUT113), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n543), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT49), .B(G64gat), .Z(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(G1333gat));
  INV_X1    g534(.A(G71gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n728), .A2(new_n736), .A3(new_n712), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n728), .A2(new_n659), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(new_n736), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g539(.A1(new_n728), .A2(new_n545), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n292), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n696), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n701), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n227), .B1(new_n745), .B2(KEYINPUT114), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(KEYINPUT114), .B2(new_n745), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n691), .A2(new_n693), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n563), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n669), .A2(new_n697), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT51), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n694), .A2(new_n753), .A3(new_n750), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n698), .A2(new_n701), .A3(new_n227), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT115), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n747), .B1(new_n755), .B2(new_n757), .ZN(G1336gat));
  AOI21_X1  g557(.A(new_n228), .B1(new_n744), .B2(new_n543), .ZN(new_n759));
  NOR4_X1   g558(.A1(new_n755), .A2(G92gat), .A3(new_n479), .A4(new_n323), .ZN(new_n760));
  OR3_X1    g559(.A1(new_n759), .A2(new_n760), .A3(KEYINPUT52), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT52), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1337gat));
  NAND3_X1  g562(.A1(new_n749), .A2(KEYINPUT51), .A3(new_n751), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n753), .B1(new_n694), .B2(new_n750), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(G99gat), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n766), .A2(new_n767), .A3(new_n712), .A4(new_n698), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n744), .A2(new_n659), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(new_n767), .ZN(G1338gat));
  NAND3_X1  g569(.A1(new_n696), .A2(new_n545), .A3(new_n743), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G106gat), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n497), .A2(G106gat), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n698), .B(new_n774), .C1(new_n752), .C2(new_n754), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(KEYINPUT116), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n766), .A2(new_n778), .A3(new_n698), .A4(new_n774), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n772), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT53), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n781), .B1(new_n780), .B2(KEYINPUT53), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n776), .B1(new_n782), .B2(new_n783), .ZN(G1339gat));
  INV_X1    g583(.A(new_n292), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n237), .A2(new_n267), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n297), .A2(new_n295), .A3(new_n298), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT99), .B1(new_n300), .B2(new_n303), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n316), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n317), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n321), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n314), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(new_n321), .A3(new_n790), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n794), .B(KEYINPUT54), .C1(new_n318), .C2(new_n308), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n320), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n793), .A2(new_n795), .A3(KEYINPUT55), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT118), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n320), .B1(new_n796), .B2(new_n797), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n804), .A3(new_n800), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n636), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n626), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n615), .A2(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n633), .A2(new_n628), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n698), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n679), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  AND4_X1   g610(.A1(new_n679), .A2(new_n802), .A3(new_n809), .A4(new_n805), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n785), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n294), .A2(new_n697), .A3(new_n323), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n815), .A2(new_n729), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n541), .A2(new_n543), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n636), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n815), .A2(new_n551), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n408), .A2(new_n543), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n822), .A2(new_n354), .A3(new_n697), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n819), .A2(new_n823), .ZN(G1340gat));
  AOI21_X1  g623(.A(G120gat), .B1(new_n818), .B2(new_n698), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n822), .A2(new_n352), .A3(new_n323), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n818), .B2(new_n292), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n820), .A2(G127gat), .A3(new_n292), .A4(new_n821), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(KEYINPUT119), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(KEYINPUT119), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(G1342gat));
  NAND3_X1  g631(.A1(new_n818), .A2(new_n349), .A3(new_n679), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n822), .B2(new_n252), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(G1343gat));
  NAND2_X1  g636(.A1(new_n660), .A2(new_n821), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n815), .A2(new_n545), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(KEYINPUT57), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n801), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n803), .A2(KEYINPUT120), .A3(new_n800), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n636), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n845), .A2(new_n846), .A3(new_n810), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n845), .B2(new_n810), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n252), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n812), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n292), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n814), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n545), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n841), .B1(KEYINPUT57), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n327), .B1(new_n854), .B2(new_n636), .ZN(new_n855));
  AND4_X1   g654(.A1(new_n545), .A2(new_n816), .A3(new_n479), .A4(new_n660), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n856), .A2(new_n327), .A3(new_n636), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT58), .B1(new_n855), .B2(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1344gat));
  NAND3_X1  g661(.A1(new_n856), .A2(new_n328), .A3(new_n698), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n865), .B1(new_n815), .B2(new_n545), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n845), .A2(new_n810), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT121), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n845), .A2(new_n846), .A3(new_n810), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n679), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871));
  OR3_X1    g670(.A1(new_n252), .A2(new_n871), .A3(new_n801), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n252), .B2(new_n801), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n809), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n785), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n814), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n497), .A2(KEYINPUT57), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n866), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n323), .B1(new_n838), .B2(KEYINPUT122), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n879), .B(new_n880), .C1(KEYINPUT122), .C2(new_n838), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n864), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  AOI211_X1 g681(.A(KEYINPUT59), .B(new_n328), .C1(new_n854), .C2(new_n698), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n863), .B1(new_n882), .B2(new_n883), .ZN(G1345gat));
  NAND3_X1  g683(.A1(new_n856), .A2(new_n378), .A3(new_n292), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n854), .A2(new_n292), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n887), .B2(new_n378), .ZN(G1346gat));
  AOI21_X1  g687(.A(G162gat), .B1(new_n856), .B2(new_n679), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n252), .A2(new_n332), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n854), .B2(new_n890), .ZN(G1347gat));
  OR2_X1    g690(.A1(new_n729), .A2(new_n479), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT124), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n820), .A2(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(new_n431), .A3(new_n697), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n701), .B1(new_n813), .B2(new_n814), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n541), .A2(new_n479), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(G169gat), .B1(new_n899), .B2(new_n636), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n896), .A2(new_n900), .ZN(G1348gat));
  OAI21_X1  g700(.A(G176gat), .B1(new_n895), .B2(new_n323), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n899), .A2(new_n432), .A3(new_n698), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1349gat));
  OAI21_X1  g703(.A(G183gat), .B1(new_n895), .B2(new_n785), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n899), .A2(new_n409), .A3(new_n292), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g707(.A1(new_n899), .A2(new_n410), .A3(new_n679), .ZN(new_n909));
  OAI21_X1  g708(.A(G190gat), .B1(new_n895), .B2(new_n252), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(KEYINPUT61), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(KEYINPUT61), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(G1351gat));
  AND4_X1   g712(.A1(new_n545), .A2(new_n897), .A3(new_n543), .A4(new_n660), .ZN(new_n914));
  AOI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n636), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n893), .A2(new_n659), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n879), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n636), .A2(G197gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(G1352gat));
  INV_X1    g718(.A(G204gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n914), .A2(new_n920), .A3(new_n698), .ZN(new_n921));
  AND2_X1   g720(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n922));
  NOR2_X1   g721(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n917), .A2(new_n698), .ZN(new_n925));
  OAI221_X1 g724(.A(new_n924), .B1(new_n922), .B2(new_n921), .C1(new_n925), .C2(new_n920), .ZN(G1353gat));
  NAND3_X1  g725(.A1(new_n914), .A2(new_n454), .A3(new_n292), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n292), .B1(new_n849), .B2(new_n874), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n878), .B1(new_n928), .B2(new_n852), .ZN(new_n929));
  INV_X1    g728(.A(new_n866), .ZN(new_n930));
  AND4_X1   g729(.A1(new_n292), .A2(new_n929), .A3(new_n930), .A4(new_n916), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n454), .B1(new_n931), .B2(KEYINPUT126), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n929), .A2(new_n930), .A3(new_n292), .A4(new_n916), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT63), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n879), .A2(KEYINPUT126), .A3(new_n292), .A4(new_n916), .ZN(new_n937));
  AND4_X1   g736(.A1(KEYINPUT63), .A2(new_n937), .A3(new_n935), .A4(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n927), .B1(new_n936), .B2(new_n938), .ZN(G1354gat));
  NOR2_X1   g738(.A1(new_n917), .A2(KEYINPUT127), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n879), .A2(KEYINPUT127), .A3(new_n916), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n679), .ZN(new_n942));
  OAI21_X1  g741(.A(G218gat), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n914), .A2(new_n455), .A3(new_n679), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1355gat));
endmodule


