//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n576, new_n577, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n636, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT65), .Z(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n454), .A2(new_n460), .B1(KEYINPUT66), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n462), .B1(KEYINPUT66), .B2(new_n461), .ZN(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT67), .Z(G319));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n465), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT68), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n468), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT69), .B1(new_n470), .B2(G2104), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(new_n472), .A3(KEYINPUT3), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n480), .A2(new_n482), .B1(new_n470), .B2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G137), .ZN(new_n484));
  NAND2_X1  g059(.A1(G101), .A2(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n479), .A2(new_n486), .ZN(G160));
  NAND2_X1  g062(.A1(new_n483), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n483), .A2(new_n467), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  NOR2_X1   g068(.A1(G100), .A2(G2105), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT70), .Z(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n490), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  NOR2_X1   g073(.A1(new_n472), .A2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G102), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n480), .A2(new_n482), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(G126), .A3(new_n471), .ZN(new_n503));
  NAND2_X1  g078(.A1(G114), .A2(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n505), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(new_n467), .A3(G138), .ZN(new_n508));
  NOR3_X1   g083(.A1(new_n474), .A2(KEYINPUT71), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n507), .A2(new_n467), .A3(G138), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n510), .B1(new_n465), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n502), .A2(G138), .A3(new_n467), .A4(new_n471), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n506), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G164));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT72), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n525), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n533));
  NAND2_X1  g108(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n533), .A2(G543), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n530), .A2(new_n531), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n532), .A2(new_n521), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G88), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n524), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(new_n541), .A3(G62), .ZN(new_n542));
  NAND2_X1  g117(.A1(G75), .A2(G543), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n544));
  INV_X1    g119(.A(G62), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT75), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n539), .B1(new_n547), .B2(G651), .ZN(G166));
  NAND3_X1  g123(.A1(new_n540), .A2(G63), .A3(G651), .ZN(new_n549));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT7), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n550), .A2(KEYINPUT7), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n523), .A2(G51), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G89), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n549), .B(new_n553), .C1(new_n554), .C2(new_n537), .ZN(G286));
  INV_X1    g130(.A(G286), .ZN(G168));
  INV_X1    g131(.A(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n540), .A2(G64), .ZN(new_n558));
  NAND2_X1  g133(.A1(G77), .A2(G543), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n523), .A2(G52), .ZN(new_n561));
  INV_X1    g136(.A(G90), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n537), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(G171));
  NAND2_X1  g139(.A1(new_n540), .A2(G56), .ZN(new_n565));
  NAND2_X1  g140(.A1(G68), .A2(G543), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n557), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n523), .A2(G43), .ZN(new_n568));
  INV_X1    g143(.A(G81), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n537), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G860), .ZN(G153));
  NAND3_X1  g147(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G36), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n574), .A2(new_n577), .ZN(G188));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n544), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n537), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n581), .A2(G651), .B1(new_n582), .B2(G91), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n523), .A2(G53), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT9), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(G299));
  OR2_X1    g161(.A1(new_n560), .A2(new_n563), .ZN(G301));
  INV_X1    g162(.A(G166), .ZN(G303));
  NAND2_X1  g163(.A1(new_n523), .A2(G49), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n582), .A2(G87), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n540), .B2(G74), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G288));
  NAND3_X1  g169(.A1(new_n521), .A2(G48), .A3(G543), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT78), .Z(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n544), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n596), .B1(new_n599), .B2(G651), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n540), .A2(KEYINPUT77), .A3(G86), .A4(new_n521), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n602));
  INV_X1    g177(.A(G86), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n537), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n600), .A2(new_n605), .ZN(G305));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n532), .A2(G60), .A3(new_n535), .A4(new_n536), .ZN(new_n609));
  NAND2_X1  g184(.A1(G72), .A2(G543), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n608), .B1(new_n611), .B2(G651), .ZN(new_n612));
  AOI211_X1 g187(.A(KEYINPUT79), .B(new_n557), .C1(new_n609), .C2(new_n610), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n582), .A2(G85), .B1(G47), .B2(new_n523), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n607), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n611), .A2(G651), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT79), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n611), .A2(new_n608), .A3(G651), .ZN(new_n619));
  AND4_X1   g194(.A1(new_n607), .A2(new_n618), .A3(new_n615), .A4(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(G290));
  NAND2_X1  g197(.A1(G79), .A2(G543), .ZN(new_n623));
  INV_X1    g198(.A(G66), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n544), .B2(new_n624), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n625), .A2(G651), .B1(G54), .B2(new_n523), .ZN(new_n626));
  INV_X1    g201(.A(G92), .ZN(new_n627));
  OAI21_X1  g202(.A(KEYINPUT10), .B1(new_n537), .B2(new_n627), .ZN(new_n628));
  OR3_X1    g203(.A1(new_n537), .A2(KEYINPUT10), .A3(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G868), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(G171), .ZN(G284));
  OAI21_X1  g208(.A(new_n632), .B1(new_n631), .B2(G171), .ZN(G321));
  NAND2_X1  g209(.A1(G286), .A2(G868), .ZN(new_n635));
  INV_X1    g210(.A(G299), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G868), .ZN(G297));
  OAI21_X1  g212(.A(new_n635), .B1(new_n636), .B2(G868), .ZN(G280));
  AND3_X1   g213(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n639));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(G860), .ZN(G148));
  OR2_X1    g216(.A1(new_n567), .A2(new_n570), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(new_n631), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n640), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n643), .B1(new_n645), .B2(new_n631), .ZN(G323));
  XNOR2_X1  g221(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g222(.A1(new_n489), .A2(G123), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n492), .A2(G135), .ZN(new_n649));
  NOR2_X1   g224(.A1(G99), .A2(G2105), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(new_n467), .B2(G111), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT81), .ZN(new_n653));
  INV_X1    g228(.A(G2096), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n465), .A2(new_n499), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT12), .Z(new_n657));
  XOR2_X1   g232(.A(KEYINPUT13), .B(G2100), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n659), .ZN(G156));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2435), .ZN(new_n662));
  XOR2_X1   g237(.A(G2427), .B(G2438), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT14), .ZN(new_n665));
  XOR2_X1   g240(.A(G2451), .B(G2454), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1341), .B(G1348), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2443), .B(G2446), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n670), .B(new_n671), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G14), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G401));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2072), .B(G2078), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT18), .Z(new_n679));
  XOR2_X1   g254(.A(new_n676), .B(KEYINPUT82), .Z(new_n680));
  OAI21_X1  g255(.A(KEYINPUT17), .B1(new_n680), .B2(new_n675), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(new_n677), .Z(new_n682));
  AND2_X1   g257(.A1(new_n680), .A2(new_n675), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n679), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(new_n654), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G2100), .ZN(G227));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n689), .A2(new_n690), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n696), .A2(new_n688), .A3(new_n691), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n694), .B(new_n697), .C1(new_n688), .C2(new_n696), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT85), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT84), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n702), .B(new_n705), .ZN(G229));
  NAND2_X1  g281(.A1(new_n492), .A2(G141), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n489), .A2(G129), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n499), .A2(G105), .ZN(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT26), .Z(new_n711));
  NAND4_X1  g286(.A1(new_n707), .A2(new_n708), .A3(new_n709), .A4(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G32), .B(new_n712), .S(G29), .Z(new_n713));
  XOR2_X1   g288(.A(KEYINPUT27), .B(G1996), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT92), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n717), .A2(KEYINPUT23), .A3(G20), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT23), .ZN(new_n719));
  INV_X1    g294(.A(G20), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G16), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n718), .B(new_n721), .C1(new_n636), .C2(new_n717), .ZN(new_n722));
  INV_X1    g297(.A(G1956), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G35), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G162), .B2(new_n725), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT95), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT29), .ZN(new_n729));
  INV_X1    g304(.A(G2090), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n724), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT96), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n639), .A2(G16), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G4), .B2(G16), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT89), .B(G1348), .Z(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT31), .B(G11), .Z(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(G160), .A2(G29), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT24), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(G34), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(G34), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n743), .A2(new_n744), .A3(new_n725), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n741), .A2(G2084), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n717), .A2(G5), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G171), .B2(new_n717), .ZN(new_n748));
  INV_X1    g323(.A(G1961), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n653), .A2(new_n725), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n735), .B2(new_n737), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n740), .A2(new_n746), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(G2084), .B1(new_n741), .B2(new_n745), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT94), .Z(new_n755));
  OR2_X1    g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n717), .A2(G19), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n571), .B2(new_n717), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT90), .ZN(new_n759));
  INV_X1    g334(.A(G1341), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n729), .B2(new_n730), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n492), .A2(G139), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(new_n467), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n499), .A2(G103), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n763), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  MUX2_X1   g344(.A(G33), .B(new_n769), .S(G29), .Z(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G2072), .Z(new_n771));
  NAND2_X1  g346(.A1(G164), .A2(G29), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G27), .B2(G29), .ZN(new_n773));
  INV_X1    g348(.A(G2078), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT28), .ZN(new_n776));
  INV_X1    g351(.A(G26), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G29), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(G29), .ZN(new_n779));
  OR2_X1    g354(.A1(G104), .A2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n780), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n781));
  INV_X1    g356(.A(G128), .ZN(new_n782));
  INV_X1    g357(.A(G140), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n781), .B1(new_n488), .B2(new_n782), .C1(new_n783), .C2(new_n491), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n779), .B1(new_n784), .B2(G29), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n778), .B1(new_n785), .B2(new_n776), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(G2067), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(G2067), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(G28), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(G28), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n790), .A2(new_n791), .A3(new_n725), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n775), .A2(new_n787), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n759), .B2(new_n760), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n762), .A2(new_n771), .A3(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n733), .A2(new_n756), .A3(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT36), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT88), .ZN(new_n798));
  NAND2_X1  g373(.A1(G166), .A2(G16), .ZN(new_n799));
  NOR2_X1   g374(.A1(G16), .A2(G22), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT87), .B(G1971), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n803), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n799), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n717), .B1(new_n600), .B2(new_n605), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n717), .A2(G6), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT32), .B(G1981), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OR3_X1    g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n808), .B2(new_n809), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n807), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n717), .A2(G23), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G288), .B2(G16), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  AOI211_X1 g395(.A(KEYINPUT33), .B(new_n816), .C1(G288), .C2(G16), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(G1976), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G1976), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n819), .B2(new_n821), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n798), .B1(new_n815), .B2(new_n826), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n804), .A2(new_n806), .B1(new_n812), .B2(new_n813), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n828), .A2(KEYINPUT88), .A3(new_n823), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT34), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT34), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n827), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n717), .A2(G24), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n621), .B2(new_n717), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n836), .A2(G1986), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(G1986), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n489), .A2(G119), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n492), .A2(G131), .ZN(new_n840));
  OR2_X1    g415(.A1(G95), .A2(G2105), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n841), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  MUX2_X1   g418(.A(G25), .B(new_n843), .S(G29), .Z(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT35), .B(G1991), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT86), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n844), .B(new_n846), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n837), .A2(new_n838), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n797), .B1(new_n834), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n827), .A2(new_n829), .A3(new_n832), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n832), .B1(new_n827), .B2(new_n829), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n797), .B(new_n848), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n716), .B(new_n796), .C1(new_n849), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n773), .A2(new_n774), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(G168), .A2(G16), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(G16), .B2(G21), .ZN(new_n858));
  XNOR2_X1  g433(.A(KEYINPUT93), .B(G1966), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n854), .A2(new_n856), .A3(new_n861), .ZN(G311));
  INV_X1    g437(.A(new_n733), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n756), .A2(new_n795), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n834), .A2(new_n848), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT36), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n865), .B1(new_n867), .B2(new_n852), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n868), .A2(new_n855), .A3(new_n860), .A4(new_n716), .ZN(G150));
  NAND2_X1  g444(.A1(new_n540), .A2(G67), .ZN(new_n870));
  NAND2_X1  g445(.A1(G80), .A2(G543), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n557), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n523), .A2(G55), .ZN(new_n873));
  INV_X1    g448(.A(G93), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(new_n537), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(G860), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT37), .Z(new_n877));
  NAND2_X1  g452(.A1(new_n639), .A2(G559), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT39), .ZN(new_n879));
  XNOR2_X1  g454(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n872), .A2(new_n875), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n571), .B1(new_n872), .B2(new_n875), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n881), .B(new_n885), .Z(new_n886));
  OAI21_X1  g461(.A(new_n877), .B1(new_n886), .B2(G860), .ZN(G145));
  XNOR2_X1  g462(.A(new_n517), .B(new_n784), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n712), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(new_n769), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n769), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G142), .ZN(new_n893));
  NOR2_X1   g468(.A1(G106), .A2(G2105), .ZN(new_n894));
  OAI21_X1  g469(.A(G2104), .B1(new_n467), .B2(G118), .ZN(new_n895));
  OAI22_X1  g470(.A1(new_n491), .A2(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(G130), .B2(new_n489), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(new_n657), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n843), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n892), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT99), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n890), .A2(new_n899), .A3(new_n891), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n901), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n497), .B(KEYINPUT98), .Z(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(new_n653), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(G160), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n903), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G37), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n902), .A3(new_n900), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g489(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n915));
  OR2_X1    g490(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n916));
  OAI21_X1  g491(.A(G166), .B1(new_n616), .B2(new_n620), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n618), .A2(new_n615), .A3(new_n619), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT80), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n614), .A2(new_n607), .A3(new_n615), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(G303), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(G305), .B(G288), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n917), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n922), .B1(new_n917), .B2(new_n921), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n915), .B(new_n916), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n917), .A2(new_n921), .ZN(new_n926));
  INV_X1    g501(.A(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n917), .A2(new_n921), .A3(new_n922), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n928), .A2(KEYINPUT100), .A3(KEYINPUT42), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n639), .A2(new_n636), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n630), .A2(G299), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT41), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n644), .A2(new_n883), .A3(new_n884), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n644), .B1(new_n884), .B2(new_n883), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n885), .A2(new_n645), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n934), .B1(new_n941), .B2(new_n936), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n931), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n942), .B1(new_n935), .B2(new_n939), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT101), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n948), .A2(new_n925), .A3(new_n949), .A4(new_n930), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT101), .B1(new_n931), .B2(new_n944), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n931), .A2(new_n944), .A3(KEYINPUT102), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n947), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G868), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n882), .A2(G868), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(G295));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n954), .B2(new_n956), .ZN(new_n959));
  AOI211_X1 g534(.A(KEYINPUT103), .B(new_n955), .C1(new_n953), .C2(G868), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(G331));
  NAND2_X1  g536(.A1(G301), .A2(G168), .ZN(new_n962));
  NAND2_X1  g537(.A1(G171), .A2(G286), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n885), .ZN(new_n965));
  INV_X1    g540(.A(new_n934), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n883), .A2(new_n962), .A3(new_n884), .A4(new_n963), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT41), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n934), .B(new_n969), .ZN(new_n970));
  AND4_X1   g545(.A1(new_n884), .A2(new_n962), .A3(new_n883), .A4(new_n963), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n884), .A2(new_n883), .B1(new_n962), .B2(new_n963), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n968), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n923), .A2(new_n924), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT104), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n965), .A2(new_n967), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n935), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n928), .A2(new_n929), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n968), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n974), .A2(new_n975), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n976), .A2(new_n911), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n973), .A2(new_n986), .A3(new_n966), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n987), .B(new_n975), .C1(new_n974), .C2(new_n986), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n988), .A2(new_n976), .A3(new_n911), .A4(new_n981), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(new_n984), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT44), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n983), .A2(new_n984), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n984), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n994), .B2(KEYINPUT44), .ZN(G397));
  OR2_X1    g570(.A1(G290), .A2(G1986), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n997));
  NAND2_X1  g572(.A1(G290), .A2(G1986), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT71), .B1(new_n474), .B2(new_n508), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n465), .A2(new_n511), .A3(new_n510), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(KEYINPUT4), .B2(new_n514), .ZN(new_n1004));
  INV_X1    g579(.A(new_n504), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n483), .B2(G126), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n500), .B1(new_n1006), .B2(new_n467), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1000), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n484), .A2(new_n485), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n467), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1012), .A2(G40), .A3(new_n468), .A4(new_n478), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(G290), .A2(KEYINPUT106), .A3(G1986), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n999), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n712), .B(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G2067), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n784), .B(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n843), .B(new_n845), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1014), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1016), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT107), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  OAI211_X1 g601(.A(KEYINPUT45), .B(new_n1000), .C1(new_n1004), .C2(new_n1007), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT116), .ZN(new_n1028));
  INV_X1    g603(.A(G40), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n479), .A2(new_n486), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n517), .A2(new_n1031), .A3(KEYINPUT45), .A4(new_n1000), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1028), .A2(new_n1010), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n859), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n506), .B2(new_n516), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1030), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI211_X1 g613(.A(KEYINPUT50), .B(G1384), .C1(new_n506), .C2(new_n516), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G2084), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1035), .A2(new_n1042), .A3(KEYINPUT121), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT121), .B1(new_n1035), .B2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT113), .B(G8), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G286), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1026), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1034), .A2(new_n1033), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1046), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1026), .B(new_n1047), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT123), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT45), .B1(new_n517), .B2(new_n1000), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(KEYINPUT116), .B2(new_n1027), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1032), .A2(new_n1030), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n859), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1038), .A2(new_n1039), .A3(G2084), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1046), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT123), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1058), .A2(new_n1059), .A3(new_n1026), .A4(new_n1047), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1052), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1035), .A2(new_n1042), .A3(KEYINPUT121), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1047), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1062), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI211_X1 g643(.A(KEYINPUT122), .B(new_n1047), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1048), .A2(new_n1061), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT110), .B(G2090), .Z(new_n1071));
  NAND2_X1  g646(.A1(new_n1040), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT111), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT111), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1040), .A2(new_n1074), .A3(new_n1071), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1027), .B(KEYINPUT109), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1053), .A2(KEYINPUT108), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1013), .B1(new_n1053), .B2(KEYINPUT108), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1073), .B(new_n1075), .C1(new_n1079), .C2(G1971), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(KEYINPUT55), .ZN(new_n1082));
  NAND3_X1  g657(.A1(G303), .A2(G8), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(KEYINPUT55), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1082), .ZN(new_n1085));
  INV_X1    g660(.A(G8), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1084), .B(new_n1085), .C1(G166), .C2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1080), .A2(new_n1089), .A3(G8), .ZN(new_n1090));
  INV_X1    g665(.A(G1981), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n600), .A2(new_n605), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n582), .A2(G86), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n600), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(KEYINPUT49), .B(new_n1092), .C1(new_n1094), .C2(new_n1091), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT49), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n600), .A2(new_n605), .A3(new_n1091), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1091), .B1(new_n600), .B2(new_n1093), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(new_n1050), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1095), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(G288), .A2(new_n824), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n591), .A2(new_n593), .A3(new_n592), .A4(G1976), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1104), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1046), .ZN(new_n1111));
  INV_X1    g686(.A(G288), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(G1976), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1113), .A2(KEYINPUT114), .A3(new_n1104), .A4(new_n1103), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1102), .A2(new_n1109), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1117));
  INV_X1    g692(.A(G1971), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1117), .A2(new_n1118), .B1(new_n1071), .B2(new_n1040), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1088), .B1(new_n1119), .B2(new_n1050), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1117), .B2(G2078), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1040), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n749), .ZN(new_n1124));
  OR2_X1    g699(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1125));
  NAND2_X1  g700(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(G40), .B1(new_n466), .B2(new_n467), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1053), .A2(new_n486), .A3(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1076), .A2(KEYINPUT53), .A3(new_n1129), .A4(new_n774), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1122), .A2(new_n1124), .A3(new_n1127), .A4(new_n1130), .ZN(new_n1131));
  AND4_X1   g706(.A1(new_n1090), .A2(new_n1116), .A3(new_n1120), .A4(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n774), .A2(KEYINPUT53), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1122), .B(new_n1124), .C1(new_n1033), .C2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1070), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1123), .A2(new_n723), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT56), .B(G2072), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1139), .B1(new_n1117), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n1143));
  XNOR2_X1  g718(.A(G299), .B(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1144), .A2(KEYINPUT119), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(KEYINPUT119), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1142), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1040), .A2(G1348), .B1(G2067), .B2(new_n1110), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n630), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1079), .A2(new_n1140), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1151), .A2(KEYINPUT118), .A3(new_n1139), .A4(new_n1144), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1144), .B(new_n1139), .C1(new_n1117), .C2(new_n1141), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT120), .B(G1341), .Z(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT58), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1117), .A2(G1996), .B1(new_n1100), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n571), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT59), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1147), .A2(KEYINPUT61), .A3(new_n1153), .ZN(new_n1163));
  OR3_X1    g738(.A1(new_n1148), .A2(KEYINPUT60), .A3(new_n630), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1149), .A2(new_n630), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1148), .A2(new_n639), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT60), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1144), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1142), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT61), .B1(new_n1156), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1157), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1070), .A2(KEYINPUT125), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1138), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1175));
  AND4_X1   g750(.A1(new_n1090), .A2(new_n1116), .A3(new_n1120), .A4(new_n1134), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1067), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(KEYINPUT122), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1066), .A2(new_n1062), .A3(new_n1067), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1180), .B(new_n1181), .C1(new_n1048), .C2(new_n1061), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1175), .A2(new_n1176), .A3(G171), .A4(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1058), .A2(G286), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1090), .A2(new_n1116), .A3(new_n1120), .A4(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(KEYINPUT117), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT117), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1185), .A2(new_n1189), .A3(new_n1186), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1115), .B(KEYINPUT115), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1080), .A2(G8), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1186), .B1(new_n1192), .B2(new_n1088), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1191), .A2(new_n1090), .A3(new_n1184), .A4(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1188), .A2(new_n1190), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1102), .A2(new_n824), .A3(new_n1112), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1111), .B1(new_n1196), .B2(new_n1092), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1090), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1197), .B1(new_n1191), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1183), .A2(new_n1195), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1025), .B1(new_n1174), .B2(new_n1200), .ZN(new_n1201));
  OR2_X1    g776(.A1(new_n843), .A2(new_n845), .ZN(new_n1202));
  OAI22_X1  g777(.A1(new_n1021), .A2(new_n1202), .B1(G2067), .B2(new_n784), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1203), .A2(new_n1014), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1020), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1014), .B1(new_n1205), .B2(new_n712), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1206), .B(KEYINPUT126), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1208), .B(KEYINPUT46), .Z(new_n1209));
  NOR2_X1   g784(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  XOR2_X1   g785(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1211));
  XNOR2_X1  g786(.A(new_n1210), .B(new_n1211), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n996), .A2(new_n1013), .A3(new_n1010), .ZN(new_n1213));
  XOR2_X1   g788(.A(new_n1213), .B(KEYINPUT48), .Z(new_n1214));
  AOI211_X1 g789(.A(new_n1204), .B(new_n1212), .C1(new_n1214), .C2(new_n1023), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1201), .A2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g791(.A1(new_n992), .A2(new_n463), .A3(new_n673), .A4(new_n993), .ZN(new_n1218));
  INV_X1    g792(.A(G227), .ZN(new_n1219));
  INV_X1    g793(.A(G229), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n913), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  NOR2_X1   g795(.A1(new_n1218), .A2(new_n1221), .ZN(G308));
  OR2_X1    g796(.A1(new_n1218), .A2(new_n1221), .ZN(G225));
endmodule


