//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n211));
  NAND4_X1  g0011(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n207), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n207), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n202), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n214), .B(new_n217), .C1(new_n220), .C2(new_n223), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G226), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XOR2_X1   g0034(.A(G50), .B(G58), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G351));
  NAND3_X1  g0040(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(new_n218), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n203), .A2(G20), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT8), .B(G58), .Z(new_n245));
  NAND2_X1  g0045(.A1(new_n219), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n245), .A2(new_n247), .B1(G150), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n243), .B1(new_n244), .B2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(new_n242), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(G20), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G50), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G50), .B2(new_n252), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G222), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G77), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G223), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n261), .B1(new_n262), .B2(new_n259), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  INV_X1    g0068(.A(new_n218), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n266), .A2(new_n274), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n275), .B1(G226), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n267), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT67), .B(G179), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G169), .ZN(new_n282));
  AOI211_X1 g0082(.A(new_n258), .B(new_n281), .C1(new_n282), .C2(new_n278), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n258), .A2(KEYINPUT9), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n267), .A2(G190), .A3(new_n277), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n278), .A2(G200), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n258), .A2(KEYINPUT9), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n284), .A2(new_n285), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  XOR2_X1   g0088(.A(KEYINPUT70), .B(KEYINPUT10), .Z(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT71), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(KEYINPUT10), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT72), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n283), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G68), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n248), .A2(G50), .B1(G20), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(new_n262), .B2(new_n246), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n242), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT11), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n253), .A2(new_n295), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT12), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n297), .A2(KEYINPUT11), .A3(new_n242), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n254), .A2(G68), .A3(new_n255), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n300), .A2(new_n302), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT3), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT3), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G33), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n307), .A2(new_n309), .A3(G232), .A4(G1698), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n307), .A2(new_n309), .A3(G226), .A4(new_n260), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G97), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n266), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n276), .A2(G238), .B1(new_n271), .B2(new_n274), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT13), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n316), .B1(new_n314), .B2(new_n315), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n305), .B1(new_n319), .B2(G190), .ZN(new_n320));
  INV_X1    g0120(.A(new_n318), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT73), .B1(new_n323), .B2(G200), .ZN(new_n324));
  OAI211_X1 g0124(.A(KEYINPUT73), .B(G200), .C1(new_n317), .C2(new_n318), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n320), .B(KEYINPUT74), .C1(new_n324), .C2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT73), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n319), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n325), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT74), .B1(new_n332), .B2(new_n320), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n319), .A2(G179), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n282), .B1(new_n321), .B2(new_n322), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XOR2_X1   g0138(.A(KEYINPUT75), .B(KEYINPUT14), .Z(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT76), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n336), .A2(KEYINPUT76), .A3(new_n339), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n338), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n305), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n334), .A2(new_n346), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n245), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n348));
  XNOR2_X1  g0148(.A(KEYINPUT15), .B(G87), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n246), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n242), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n254), .A2(G77), .A3(new_n255), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n351), .B(new_n352), .C1(G77), .C2(new_n252), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n259), .A2(G232), .A3(new_n260), .ZN(new_n354));
  INV_X1    g0154(.A(G107), .ZN(new_n355));
  INV_X1    g0155(.A(G238), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n354), .B1(new_n355), .B2(new_n259), .C1(new_n263), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n266), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n275), .B1(G244), .B2(new_n276), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT68), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT68), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n358), .A2(new_n362), .A3(new_n359), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n353), .B1(new_n364), .B2(G200), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n363), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G190), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n361), .A2(new_n282), .A3(new_n363), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n369), .A2(new_n353), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n279), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT69), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n373), .A2(KEYINPUT69), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n294), .A2(new_n347), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n307), .A2(new_n309), .A3(G226), .A4(G1698), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n307), .A2(new_n309), .A3(G223), .A4(new_n260), .ZN(new_n378));
  INV_X1    g0178(.A(G87), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n377), .B(new_n378), .C1(new_n306), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n266), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n276), .A2(G232), .B1(new_n271), .B2(new_n274), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT79), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT79), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n385), .A3(new_n382), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n282), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n381), .A2(new_n279), .A3(new_n382), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT18), .ZN(new_n392));
  INV_X1    g0192(.A(new_n254), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n245), .A2(new_n255), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n393), .A2(new_n394), .B1(new_n245), .B2(new_n252), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT16), .ZN(new_n397));
  AND2_X1   g0197(.A1(G58), .A2(G68), .ZN(new_n398));
  OAI21_X1  g0198(.A(G20), .B1(new_n398), .B2(new_n202), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT78), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n248), .A2(G159), .ZN(new_n402));
  OAI211_X1 g0202(.A(KEYINPUT78), .B(G20), .C1(new_n398), .C2(new_n202), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT77), .B(new_n405), .C1(new_n259), .C2(G20), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n406), .A2(G68), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n259), .B2(G20), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n307), .A2(new_n309), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT77), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI211_X1 g0212(.A(new_n397), .B(new_n404), .C1(new_n407), .C2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n295), .B1(new_n408), .B2(new_n410), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n397), .B1(new_n414), .B2(new_n404), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n242), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n396), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n391), .A2(new_n392), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n417), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT18), .B1(new_n390), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n383), .A2(G190), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n387), .B2(new_n330), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n417), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT17), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n404), .B1(new_n407), .B2(new_n412), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT16), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(new_n242), .A3(new_n415), .ZN(new_n427));
  AOI21_X1  g0227(.A(G200), .B1(new_n384), .B2(new_n386), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n427), .B(new_n396), .C1(new_n428), .C2(new_n421), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n418), .A2(new_n420), .A3(new_n424), .A4(new_n431), .ZN(new_n432));
  XOR2_X1   g0232(.A(new_n432), .B(KEYINPUT80), .Z(new_n433));
  NOR2_X1   g0233(.A1(new_n376), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT83), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n307), .A2(new_n309), .A3(G244), .A4(new_n260), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT4), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n260), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G283), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n307), .A2(new_n309), .A3(G250), .A4(G1698), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT82), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT82), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n259), .A2(new_n445), .A3(G250), .A4(G1698), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n436), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n251), .A2(G45), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n271), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n273), .A2(G1), .ZN(new_n455));
  INV_X1    g0255(.A(new_n452), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n450), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n436), .ZN(new_n458));
  INV_X1    g0258(.A(G257), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n454), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n435), .B1(new_n448), .B2(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n444), .A2(new_n446), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n266), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n460), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(KEYINPUT83), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n282), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n355), .B1(new_n408), .B2(new_n410), .ZN(new_n469));
  INV_X1    g0269(.A(G97), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(new_n355), .A3(KEYINPUT6), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT6), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G97), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n355), .A2(KEYINPUT81), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT81), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G107), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n471), .A2(new_n473), .A3(new_n475), .A4(new_n477), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n219), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n262), .A2(G20), .A3(G33), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n469), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  OR2_X1    g0283(.A1(new_n483), .A2(new_n243), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n252), .A2(G97), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n251), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n252), .A2(new_n486), .A3(new_n218), .A4(new_n241), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n485), .B1(new_n488), .B2(G97), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n448), .A2(new_n460), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n484), .A2(new_n489), .B1(new_n490), .B2(new_n279), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n468), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n461), .A2(G190), .A3(new_n466), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n489), .B1(new_n483), .B2(new_n243), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n330), .B1(new_n464), .B2(new_n465), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT84), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n493), .B2(new_n496), .ZN(new_n499));
  OAI211_X1 g0299(.A(KEYINPUT85), .B(new_n492), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n492), .B1(new_n498), .B2(new_n499), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT85), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT19), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n219), .B1(new_n312), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n379), .A2(new_n470), .A3(new_n355), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n505), .A2(KEYINPUT88), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT88), .B1(new_n505), .B2(new_n506), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n504), .B1(new_n246), .B2(new_n470), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT89), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n259), .A2(new_n219), .A3(G68), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT89), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(new_n504), .C1(new_n246), .C2(new_n470), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n242), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n349), .A2(new_n253), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n436), .A2(G274), .A3(new_n455), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n436), .A2(G250), .A3(new_n449), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT86), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT86), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n307), .A2(new_n309), .A3(G238), .A4(new_n260), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n307), .A2(new_n309), .A3(G244), .A4(G1698), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G116), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n266), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n524), .A2(G190), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n488), .A2(G87), .ZN(new_n531));
  INV_X1    g0331(.A(new_n523), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n529), .B1(new_n532), .B2(new_n521), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G200), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n518), .A2(new_n530), .A3(new_n531), .A4(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT87), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n533), .B2(new_n280), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n524), .A2(KEYINPUT87), .A3(new_n279), .A4(new_n529), .ZN(new_n538));
  INV_X1    g0338(.A(new_n349), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n488), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n516), .A2(new_n517), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n533), .A2(new_n282), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n537), .A2(new_n538), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n535), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n441), .B(new_n219), .C1(G33), .C2(new_n470), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT20), .ZN(new_n546));
  INV_X1    g0346(.A(G116), .ZN(new_n547));
  AOI22_X1  g0347(.A1(KEYINPUT90), .A2(new_n546), .B1(new_n547), .B2(G20), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n545), .A2(new_n548), .A3(new_n242), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n546), .A2(KEYINPUT90), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n252), .A2(new_n547), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n488), .B2(new_n547), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n549), .A2(new_n550), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n307), .A2(new_n309), .A3(G264), .A4(G1698), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n307), .A2(new_n309), .A3(G257), .A4(new_n260), .ZN(new_n558));
  INV_X1    g0358(.A(G303), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n557), .B(new_n558), .C1(new_n559), .C2(new_n259), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n266), .ZN(new_n561));
  XNOR2_X1  g0361(.A(KEYINPUT5), .B(G41), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n562), .A2(new_n455), .B1(new_n269), .B2(new_n270), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n563), .A2(G270), .B1(new_n271), .B2(new_n453), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n564), .A3(G190), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n561), .A2(new_n564), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n556), .B(new_n565), .C1(new_n566), .C2(new_n330), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n561), .A2(new_n564), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n555), .A2(new_n568), .A3(G169), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT21), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n566), .A2(G179), .A3(new_n555), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n555), .A2(new_n568), .A3(KEYINPUT21), .A4(G169), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n567), .A2(new_n571), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n544), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n457), .A2(G264), .A3(new_n436), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n454), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n307), .A2(new_n309), .A3(G257), .A4(G1698), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n307), .A2(new_n309), .A3(G250), .A4(new_n260), .ZN(new_n579));
  INV_X1    g0379(.A(G294), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n578), .B(new_n579), .C1(new_n306), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n266), .ZN(new_n582));
  INV_X1    g0382(.A(G190), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n577), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n454), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT91), .B1(new_n563), .B2(G264), .ZN(new_n586));
  AND4_X1   g0386(.A1(KEYINPUT91), .A2(new_n457), .A3(G264), .A4(new_n436), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n582), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT92), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n563), .A2(KEYINPUT91), .A3(G264), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT91), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n576), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT92), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n594), .A3(new_n582), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n585), .B1(new_n589), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n584), .B1(new_n596), .B2(G200), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n253), .A2(KEYINPUT25), .A3(new_n355), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT25), .B1(new_n253), .B2(new_n355), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n599), .A2(new_n600), .B1(new_n355), .B2(new_n487), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT24), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n259), .A2(new_n219), .A3(G87), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT22), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT23), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n219), .B2(G107), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n355), .A2(KEYINPUT23), .A3(G20), .ZN(new_n607));
  INV_X1    g0407(.A(new_n527), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n606), .A2(new_n607), .B1(new_n608), .B2(new_n219), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n602), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n604), .A2(new_n602), .A3(new_n609), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n601), .B1(new_n613), .B2(new_n242), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n597), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n593), .A2(new_n594), .A3(new_n582), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n594), .B1(new_n593), .B2(new_n582), .ZN(new_n617));
  OAI211_X1 g0417(.A(G179), .B(new_n454), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n577), .A2(new_n582), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G169), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n612), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n242), .B1(new_n622), .B2(new_n610), .ZN(new_n623));
  INV_X1    g0423(.A(new_n601), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n575), .A2(new_n615), .A3(new_n626), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n434), .A2(new_n500), .A3(new_n503), .A4(new_n627), .ZN(G372));
  INV_X1    g0428(.A(KEYINPUT93), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n541), .B(new_n542), .C1(new_n280), .C2(new_n533), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n468), .A2(new_n491), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n535), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n630), .B1(new_n633), .B2(KEYINPUT26), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  INV_X1    g0435(.A(new_n544), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n631), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n629), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n572), .A2(new_n573), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n626), .A2(new_n571), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n615), .A3(new_n632), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n501), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n637), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n632), .A2(new_n468), .A3(new_n491), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n635), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n645), .A2(new_n647), .A3(KEYINPUT93), .A4(new_n630), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n638), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n434), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT94), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n418), .A2(new_n420), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n372), .B1(new_n332), .B2(new_n320), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(new_n346), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n424), .A2(new_n431), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n291), .A2(new_n293), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n283), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n651), .A2(new_n658), .ZN(G369));
  NAND3_X1  g0459(.A1(new_n251), .A2(new_n219), .A3(G13), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(G213), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n615), .B(new_n626), .C1(new_n614), .C2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n621), .A2(new_n625), .A3(new_n665), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n639), .A2(new_n571), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n666), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT96), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n626), .A2(new_n665), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n555), .A2(new_n665), .ZN(new_n676));
  XOR2_X1   g0476(.A(new_n676), .B(KEYINPUT95), .Z(new_n677));
  NAND2_X1  g0477(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n574), .B2(new_n677), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n667), .B2(new_n668), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n675), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n215), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n506), .A2(G116), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n685), .A2(new_n251), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n223), .B2(new_n685), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT28), .Z(new_n690));
  NAND2_X1  g0490(.A1(new_n649), .A2(new_n666), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT29), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n642), .A2(KEYINPUT98), .A3(new_n643), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n631), .A2(new_n635), .A3(new_n636), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n630), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(KEYINPUT26), .B2(new_n633), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT98), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n641), .B2(new_n501), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n694), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(KEYINPUT29), .A3(new_n666), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n464), .A2(KEYINPUT83), .A3(new_n465), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT83), .B1(new_n464), .B2(new_n465), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n589), .A2(new_n595), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n561), .A2(new_n564), .A3(G179), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n533), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n705), .A2(KEYINPUT30), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n708), .B1(new_n616), .B2(new_n617), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n467), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n706), .A2(new_n454), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n533), .A2(new_n568), .A3(new_n279), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n490), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n709), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT31), .B1(new_n717), .B2(new_n665), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n706), .A2(new_n461), .A3(new_n466), .A4(new_n708), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n721), .A2(new_n710), .B1(new_n713), .B2(new_n715), .ZN(new_n722));
  AOI211_X1 g0522(.A(new_n720), .B(new_n666), .C1(new_n722), .C2(new_n709), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n719), .B1(new_n723), .B2(KEYINPUT97), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n503), .A2(new_n500), .A3(new_n627), .A4(new_n666), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n717), .A2(new_n665), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT97), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(new_n720), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n724), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n702), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n690), .B1(new_n731), .B2(G1), .ZN(G364));
  INV_X1    g0532(.A(G13), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n251), .B1(new_n734), .B2(G45), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n685), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n218), .B1(G20), .B2(new_n282), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT32), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n219), .A2(G179), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G190), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G159), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n279), .A2(new_n219), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n583), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G58), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n259), .B1(new_n741), .B2(new_n746), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n470), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n741), .B2(new_n746), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G87), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n742), .A2(new_n583), .A3(G200), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n757), .B(new_n760), .C1(new_n355), .C2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n747), .A2(G190), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n751), .B(new_n762), .C1(G50), .C2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n747), .A2(new_n583), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT101), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n747), .A2(new_n743), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n771), .A2(KEYINPUT100), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(KEYINPUT100), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n765), .B1(new_n295), .B2(new_n770), .C1(new_n262), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n776), .A2(new_n771), .B1(new_n749), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n744), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n259), .B1(new_n779), .B2(G329), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n580), .B2(new_n755), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n782), .A2(new_n761), .B1(new_n758), .B2(new_n559), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n778), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G326), .ZN(new_n785));
  XOR2_X1   g0585(.A(KEYINPUT33), .B(G317), .Z(new_n786));
  OAI221_X1 g0586(.A(new_n784), .B1(new_n785), .B2(new_n763), .C1(new_n770), .C2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n740), .B1(new_n775), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n739), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n684), .A2(new_n409), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n793), .A2(G355), .B1(new_n547), .B2(new_n684), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n236), .A2(G45), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT99), .Z(new_n796));
  NOR2_X1   g0596(.A1(new_n684), .A2(new_n259), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(G45), .B2(new_n222), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n794), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n738), .B(new_n788), .C1(new_n792), .C2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n791), .B(KEYINPUT102), .Z(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n679), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT103), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n679), .A2(G330), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n680), .A2(new_n738), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(G396));
  NAND3_X1  g0606(.A1(new_n370), .A2(new_n371), .A3(new_n666), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n353), .A2(new_n665), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n365), .B2(new_n367), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n370), .A2(new_n371), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n691), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n811), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n649), .A2(new_n666), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n737), .B1(new_n815), .B2(new_n730), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n730), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n739), .A2(new_n789), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n738), .B1(new_n262), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n409), .B1(new_n744), .B2(new_n776), .ZN(new_n820));
  INV_X1    g0620(.A(new_n761), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G87), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n355), .B2(new_n758), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n820), .B(new_n823), .C1(G97), .C2(new_n754), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n824), .B1(new_n580), .B2(new_n749), .C1(new_n559), .C2(new_n763), .ZN(new_n825));
  INV_X1    g0625(.A(new_n774), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(G116), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n770), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G283), .ZN(new_n829));
  INV_X1    g0629(.A(new_n749), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n764), .A2(G137), .B1(new_n830), .B2(G143), .ZN(new_n831));
  INV_X1    g0631(.A(G150), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n774), .B2(new_n745), .C1(new_n832), .C2(new_n770), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT34), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n259), .B1(new_n744), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(G50), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n837), .A2(new_n758), .B1(new_n761), .B2(new_n295), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n836), .B(new_n838), .C1(G58), .C2(new_n754), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n827), .A2(new_n829), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n819), .B1(new_n740), .B2(new_n840), .C1(new_n813), .C2(new_n790), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n817), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G384));
  NOR2_X1   g0643(.A1(new_n734), .A2(new_n251), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT113), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n242), .B1(new_n425), .B2(KEYINPUT16), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT106), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n413), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(KEYINPUT106), .B(new_n242), .C1(new_n425), .C2(KEYINPUT16), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n395), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(new_n663), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n432), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT107), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n429), .B1(new_n850), .B2(new_n663), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n850), .A2(new_n390), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n853), .B(KEYINPUT37), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n391), .A2(new_n417), .ZN(new_n857));
  XNOR2_X1  g0657(.A(KEYINPUT108), .B(KEYINPUT37), .ZN(new_n858));
  INV_X1    g0658(.A(new_n663), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n417), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n857), .A2(new_n429), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n412), .A2(G68), .A3(new_n406), .ZN(new_n863));
  INV_X1    g0663(.A(new_n404), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT16), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n847), .B1(new_n865), .B2(new_n243), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n426), .A3(new_n849), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n396), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n423), .B1(new_n868), .B2(new_n859), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n391), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n853), .B1(new_n871), .B2(KEYINPUT37), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n852), .B1(new_n862), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n854), .B2(new_n855), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT107), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n861), .A3(new_n856), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n874), .B1(new_n432), .B2(new_n851), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n873), .A2(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n723), .A2(new_n718), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n725), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT112), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n344), .B1(new_n328), .B2(new_n333), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n305), .A2(new_n665), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n885), .B1(new_n332), .B2(new_n320), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n344), .B2(new_n345), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n811), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n881), .A2(new_n882), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n882), .B1(new_n881), .B2(new_n889), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n879), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n845), .B1(new_n892), .B2(KEYINPUT40), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n878), .B1(new_n862), .B2(new_n872), .ZN(new_n894));
  INV_X1    g0694(.A(new_n852), .ZN(new_n895));
  AND4_X1   g0695(.A1(new_n857), .A2(new_n429), .A3(new_n858), .A4(new_n860), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n869), .B2(new_n870), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n898), .B2(new_n853), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n895), .B1(new_n899), .B2(new_n876), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n894), .B1(new_n900), .B2(KEYINPUT38), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n881), .A2(new_n889), .A3(new_n882), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n881), .A2(new_n889), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT112), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(KEYINPUT113), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n893), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n894), .A2(KEYINPUT110), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT110), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n877), .A2(new_n910), .A3(new_n878), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT109), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n655), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n424), .A2(KEYINPUT109), .A3(new_n431), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n913), .A2(new_n652), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n857), .A2(new_n429), .A3(new_n860), .ZN(new_n916));
  INV_X1    g0716(.A(new_n858), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n915), .A2(new_n860), .B1(new_n896), .B2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n909), .A2(new_n911), .B1(new_n919), .B2(new_n874), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n881), .A2(new_n889), .A3(KEYINPUT40), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n908), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n434), .A2(new_n881), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  INV_X1    g0725(.A(G330), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n652), .A2(new_n859), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n807), .B(KEYINPUT104), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT105), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n814), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n886), .A2(new_n888), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n920), .B2(KEYINPUT39), .ZN(new_n936));
  INV_X1    g0736(.A(new_n346), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(new_n665), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n929), .B1(new_n934), .B2(new_n879), .C1(new_n936), .C2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n693), .A2(new_n434), .A3(new_n701), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n658), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT111), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n941), .B(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n844), .B1(new_n928), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n928), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n479), .A2(new_n480), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(KEYINPUT35), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(KEYINPUT35), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n949), .A2(G116), .A3(new_n220), .A4(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n222), .A2(new_n262), .A3(new_n398), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(G68), .B2(new_n201), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n733), .A2(G1), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n947), .B(new_n952), .C1(new_n954), .C2(new_n955), .ZN(G367));
  NAND2_X1  g0756(.A1(new_n797), .A2(new_n232), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n791), .B(new_n739), .C1(new_n684), .C2(new_n539), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n738), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n518), .A2(new_n531), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n665), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n632), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n630), .B2(new_n961), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n755), .A2(new_n295), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G58), .B2(new_n759), .ZN(new_n965));
  INV_X1    g0765(.A(G137), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n259), .B1(new_n744), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G77), .B2(new_n821), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n965), .B(new_n968), .C1(new_n832), .C2(new_n749), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G143), .B2(new_n764), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n745), .B2(new_n770), .C1(new_n201), .C2(new_n774), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n259), .B1(new_n779), .B2(G317), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n470), .B2(new_n761), .C1(new_n355), .C2(new_n755), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G311), .B2(new_n764), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n758), .A2(new_n547), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n749), .A2(new_n559), .B1(KEYINPUT46), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(KEYINPUT46), .B2(new_n975), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n782), .B2(new_n774), .C1(new_n580), .C2(new_n770), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n971), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT47), .Z(new_n981));
  OAI221_X1 g0781(.A(new_n959), .B1(new_n963), .B2(new_n801), .C1(new_n981), .C2(new_n740), .ZN(new_n982));
  INV_X1    g0782(.A(new_n731), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n494), .A2(new_n665), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n501), .A2(new_n984), .B1(new_n492), .B2(new_n666), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n675), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT45), .Z(new_n987));
  NOR2_X1   g0787(.A1(new_n675), .A2(new_n985), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(new_n682), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n669), .B(new_n680), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(new_n672), .Z(new_n993));
  AOI21_X1  g0793(.A(new_n983), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n685), .B(KEYINPUT41), .Z(new_n995));
  OAI21_X1  g0795(.A(new_n735), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT116), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n673), .A2(new_n985), .ZN(new_n1000));
  OR3_X1    g0800(.A1(new_n1000), .A2(KEYINPUT114), .A3(KEYINPUT42), .ZN(new_n1001));
  OAI21_X1  g0801(.A(KEYINPUT114), .B1(new_n1000), .B2(KEYINPUT42), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n621), .B(new_n625), .C1(new_n498), .C2(new_n499), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n665), .B1(new_n1004), .B2(new_n492), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n1000), .B2(KEYINPUT42), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n998), .B(new_n999), .C1(new_n1003), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT115), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1003), .A2(new_n1006), .A3(new_n998), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n997), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1012), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1014), .A2(KEYINPUT116), .A3(new_n1010), .A4(new_n1009), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n681), .A2(new_n985), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n996), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1017), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n982), .B1(new_n1019), .B2(new_n1020), .ZN(G387));
  NAND2_X1  g0821(.A1(new_n993), .A2(new_n736), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n409), .B1(new_n744), .B2(new_n785), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n764), .A2(G322), .B1(new_n830), .B2(G317), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n774), .B2(new_n559), .C1(new_n776), .C2(new_n770), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G294), .A2(new_n759), .B1(new_n754), .B2(G283), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT49), .Z(new_n1031));
  AOI211_X1 g0831(.A(new_n1023), .B(new_n1031), .C1(G116), .C2(new_n821), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n259), .B1(new_n744), .B2(new_n832), .C1(new_n470), .C2(new_n761), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n755), .A2(new_n349), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(G77), .C2(new_n759), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n771), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G50), .A2(new_n830), .B1(new_n1036), .B2(G68), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1035), .B(new_n1037), .C1(new_n745), .C2(new_n763), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n245), .B2(new_n828), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n739), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n797), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n245), .A2(new_n837), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT50), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  AOI211_X1 g0844(.A(G45), .B(new_n687), .C1(G68), .C2(G77), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1041), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1046), .A2(KEYINPUT117), .B1(G45), .B2(new_n229), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(KEYINPUT117), .B2(new_n1046), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n793), .A2(new_n687), .B1(new_n355), .B2(new_n684), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT118), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n1052), .A2(new_n791), .A3(new_n739), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n738), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1040), .B(new_n1055), .C1(new_n669), .C2(new_n801), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n731), .A2(new_n993), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n685), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n731), .A2(new_n993), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1022), .B(new_n1056), .C1(new_n1059), .C2(new_n1060), .ZN(G393));
  OR2_X1    g0861(.A1(new_n991), .A2(KEYINPUT119), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n991), .A2(KEYINPUT119), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n736), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1058), .B1(new_n991), .B2(new_n1057), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1057), .B2(new_n991), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n985), .A2(G20), .A3(new_n790), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT120), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1041), .A2(new_n239), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n792), .B1(new_n215), .B2(new_n470), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n737), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n755), .A2(new_n547), .B1(new_n758), .B2(new_n782), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n409), .B1(new_n744), .B2(new_n777), .C1(new_n355), .C2(new_n761), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n580), .B2(new_n771), .ZN(new_n1075));
  INV_X1    g0875(.A(G317), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n763), .A2(new_n1076), .B1(new_n749), .B2(new_n776), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT121), .B(KEYINPUT52), .Z(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n559), .B2(new_n770), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n763), .A2(new_n832), .B1(new_n749), .B2(new_n745), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT51), .Z(new_n1082));
  AOI21_X1  g0882(.A(new_n409), .B1(new_n779), .B2(G143), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n759), .A2(G68), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n754), .A2(G77), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1083), .A2(new_n822), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n826), .B2(new_n245), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n201), .B2(new_n770), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1080), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1071), .B1(new_n1089), .B2(new_n739), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1068), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1064), .A2(new_n1066), .A3(new_n1091), .ZN(G390));
  NAND2_X1  g0892(.A1(new_n934), .A2(new_n939), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n936), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n730), .A2(new_n811), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n926), .B1(new_n725), .B2(new_n880), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n889), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1095), .B(new_n933), .C1(KEYINPUT122), .C2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n920), .A2(new_n938), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n700), .A2(new_n666), .A3(new_n813), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n930), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n933), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1094), .A2(new_n1098), .A3(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1093), .A2(new_n936), .B1(new_n1102), .B2(new_n1099), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1096), .A2(KEYINPUT122), .A3(new_n889), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(new_n735), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n936), .A2(new_n789), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n818), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n737), .B1(new_n245), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n828), .A2(G107), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n826), .A2(G97), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n761), .A2(new_n295), .B1(new_n744), .B2(new_n580), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT124), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G283), .B2(new_n764), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n760), .A2(new_n1085), .A3(new_n409), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G116), .B2(new_n830), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1112), .A2(new_n1113), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT54), .B(G143), .Z(new_n1120));
  AOI22_X1  g0920(.A1(new_n826), .A2(new_n1120), .B1(G159), .B2(new_n754), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n966), .B2(new_n770), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT123), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n409), .B1(new_n779), .B2(G125), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n201), .B2(new_n761), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G132), .B2(new_n830), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n759), .A2(G150), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT53), .Z(new_n1128));
  INV_X1    g0928(.A(G128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1126), .B(new_n1128), .C1(new_n1129), .C2(new_n763), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1119), .B1(new_n1123), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1111), .B1(new_n1131), .B2(new_n739), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1109), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1108), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1097), .B1(new_n1095), .B2(new_n933), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n932), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1095), .A2(new_n933), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1096), .A2(new_n813), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n933), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1137), .A2(new_n930), .A3(new_n1100), .A4(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1136), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n434), .A2(new_n1096), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n942), .A2(new_n658), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1107), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1144), .B1(new_n1136), .B2(new_n1141), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1104), .B(new_n1148), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1147), .A2(new_n685), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1134), .A2(new_n1150), .ZN(G378));
  NOR2_X1   g0951(.A1(new_n258), .A2(new_n663), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT126), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n294), .B(new_n1154), .ZN(new_n1155));
  XOR2_X1   g0955(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1155), .B(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n789), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n355), .A2(new_n749), .B1(new_n771), .B2(new_n349), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n272), .B(new_n409), .C1(new_n744), .C2(new_n782), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n750), .A2(new_n761), .B1(new_n758), .B2(new_n262), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1160), .A2(new_n964), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n470), .B2(new_n770), .C1(new_n547), .C2(new_n763), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT58), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G50), .B1(new_n306), .B2(new_n272), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n259), .B2(G41), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n759), .A2(new_n1120), .B1(new_n754), .B2(G150), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n749), .B2(new_n1129), .C1(new_n966), .C2(new_n771), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n770), .A2(new_n835), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(G125), .C2(new_n764), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n821), .A2(G159), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G33), .B(G41), .C1(new_n779), .C2(G124), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1165), .B(new_n1167), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n740), .B1(new_n1178), .B2(KEYINPUT125), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(KEYINPUT125), .B2(new_n1178), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n818), .A2(new_n201), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1159), .A2(new_n737), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1158), .ZN(new_n1184));
  OAI21_X1  g0984(.A(G330), .B1(new_n920), .B2(new_n921), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1184), .B1(new_n908), .B2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1158), .C1(new_n893), .C2(new_n907), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n940), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n905), .A2(KEYINPUT113), .A3(new_n906), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT113), .B1(new_n905), .B2(new_n906), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1186), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n1158), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n908), .A2(new_n1186), .A3(new_n1184), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n1194), .A3(new_n941), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1189), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1183), .B1(new_n1196), .B2(new_n736), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1189), .A2(new_n1195), .B1(new_n1149), .B2(new_n1145), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n685), .B1(new_n1198), .B2(KEYINPUT57), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT127), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1189), .A2(new_n1200), .A3(new_n1195), .ZN(new_n1201));
  OAI211_X1 g1001(.A(KEYINPUT127), .B(new_n940), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT57), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1149), .B2(new_n1145), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1197), .B1(new_n1199), .B2(new_n1205), .ZN(G375));
  INV_X1    g1006(.A(new_n995), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1136), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1146), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n409), .B1(new_n744), .B2(new_n559), .C1(new_n262), .C2(new_n761), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1210), .B(new_n1034), .C1(G97), .C2(new_n759), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n782), .B2(new_n749), .C1(new_n580), .C2(new_n763), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G107), .B2(new_n826), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n828), .A2(G116), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n828), .A2(new_n1120), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n966), .A2(new_n749), .B1(new_n771), .B2(new_n832), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n763), .A2(new_n835), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n755), .A2(new_n837), .B1(new_n758), .B2(new_n745), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n259), .B1(new_n744), .B2(new_n1129), .C1(new_n750), .C2(new_n761), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1213), .A2(new_n1214), .B1(new_n1215), .B2(new_n1220), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n737), .B1(G68), .B2(new_n1110), .C1(new_n1221), .C2(new_n740), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1139), .B2(new_n789), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n1142), .B2(new_n736), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1209), .A2(new_n1224), .ZN(G381));
  NOR4_X1   g1025(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n1224), .A3(new_n1209), .ZN(new_n1227));
  OR4_X1    g1027(.A1(G387), .A2(new_n1227), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1028(.A(G378), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n664), .A2(G213), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G407), .B(G213), .C1(G375), .C2(new_n1232), .ZN(G409));
  OAI211_X1 g1033(.A(G378), .B(new_n1197), .C1(new_n1199), .C2(new_n1205), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1149), .A2(new_n1145), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1196), .A2(new_n1207), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1182), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1201), .A2(new_n736), .A3(new_n1202), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1229), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1234), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1230), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1208), .B1(new_n1148), .B2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1136), .A2(new_n1141), .A3(KEYINPUT60), .A4(new_n1144), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n685), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1224), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n842), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(G384), .A3(new_n1224), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1231), .A2(G2897), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1249), .A2(G2897), .A3(new_n1231), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT61), .B1(new_n1241), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1241), .B2(new_n1249), .ZN(new_n1258));
  INV_X1    g1058(.A(G390), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G387), .A2(new_n1259), .ZN(new_n1260));
  XOR2_X1   g1060(.A(G393), .B(G396), .Z(new_n1261));
  INV_X1    g1061(.A(new_n1020), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(new_n996), .A3(new_n1018), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n982), .A3(G390), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1260), .A2(new_n1261), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1261), .B1(new_n1260), .B2(new_n1264), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1231), .B1(new_n1234), .B2(new_n1239), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1268), .A2(KEYINPUT63), .A3(new_n1250), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1256), .A2(new_n1258), .A3(new_n1267), .A4(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT62), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1268), .A2(new_n1271), .A3(new_n1250), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1268), .B2(new_n1254), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1271), .B1(new_n1268), .B2(new_n1250), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1270), .B1(new_n1276), .B2(new_n1267), .ZN(G405));
  AND2_X1   g1077(.A1(G375), .A2(new_n1229), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1234), .ZN(new_n1279));
  OR3_X1    g1079(.A1(new_n1278), .A2(new_n1279), .A3(new_n1250), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1250), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1267), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1280), .A2(new_n1267), .A3(new_n1281), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(G402));
endmodule


