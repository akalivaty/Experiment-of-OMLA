//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT67), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G567), .B1(G2106), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NOR3_X1   g045(.A1(new_n470), .A2(new_n462), .A3(G2105), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT69), .B1(new_n467), .B2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G101), .ZN(new_n474));
  OAI22_X1  g049(.A1(new_n468), .A2(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n476), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n467), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n475), .A2(new_n478), .ZN(G160));
  INV_X1    g054(.A(new_n468), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n466), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT70), .B(G114), .ZN(new_n490));
  OAI211_X1 g065(.A(G2104), .B(new_n489), .C1(new_n490), .C2(new_n467), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n466), .A2(G126), .A3(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n467), .A2(G138), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n496));
  AOI21_X1  g071(.A(KEYINPUT3), .B1(new_n464), .B2(G2104), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n463), .B2(new_n465), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT71), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n500), .A2(KEYINPUT4), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n476), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n493), .B1(new_n503), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n507), .A2(KEYINPUT6), .A3(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT6), .B1(new_n507), .B2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(G50), .A2(new_n512), .B1(new_n515), .B2(G88), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n516), .A2(KEYINPUT73), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(G166));
  NAND2_X1  g099(.A1(new_n515), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n512), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n528), .A2(new_n529), .B1(new_n513), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n525), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(G651), .A2(new_n538), .B1(new_n515), .B2(G90), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n512), .A2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n518), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n512), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n515), .A2(G81), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n512), .A2(new_n554), .A3(G53), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n514), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(G651), .A2(new_n559), .B1(new_n515), .B2(G91), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G168), .ZN(G286));
  INV_X1    g137(.A(G166), .ZN(G303));
  NAND2_X1  g138(.A1(new_n515), .A2(G87), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n512), .A2(G49), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  AOI22_X1  g142(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n518), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT76), .ZN(new_n570));
  AOI22_X1  g145(.A1(G48), .A2(new_n512), .B1(new_n515), .B2(G86), .ZN(new_n571));
  OR3_X1    g146(.A1(new_n568), .A2(KEYINPUT76), .A3(new_n518), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n518), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(KEYINPUT77), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(KEYINPUT77), .ZN(new_n578));
  AOI22_X1  g153(.A1(G47), .A2(new_n512), .B1(new_n515), .B2(G85), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n515), .A2(G92), .ZN(new_n582));
  XOR2_X1   g157(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT79), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n582), .A2(new_n584), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n514), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(G651), .A2(new_n589), .B1(new_n512), .B2(G54), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n581), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n581), .B1(new_n592), .B2(G868), .ZN(G321));
  NOR2_X1   g169(.A1(G299), .A2(G868), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(G868), .B2(G168), .ZN(G280));
  XOR2_X1   g171(.A(G280), .B(KEYINPUT80), .Z(G297));
  INV_X1    g172(.A(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n592), .B1(new_n598), .B2(G860), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT81), .ZN(G148));
  OAI21_X1  g175(.A(KEYINPUT82), .B1(new_n548), .B2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n592), .A2(new_n598), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  MUX2_X1   g178(.A(KEYINPUT82), .B(new_n601), .S(new_n603), .Z(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g180(.A(new_n473), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n476), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  INV_X1    g184(.A(G2100), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n614));
  INV_X1    g189(.A(G111), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n613), .A2(new_n614), .B1(new_n615), .B2(G2105), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n614), .B2(new_n613), .ZN(new_n617));
  INV_X1    g192(.A(G135), .ZN(new_n618));
  INV_X1    g193(.A(G123), .ZN(new_n619));
  OAI221_X1 g194(.A(new_n617), .B1(new_n468), .B2(new_n618), .C1(new_n619), .C2(new_n482), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND3_X1  g196(.A1(new_n611), .A2(new_n612), .A3(new_n621), .ZN(G156));
  INV_X1    g197(.A(KEYINPUT14), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n626), .B2(new_n625), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2451), .B(G2454), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  XOR2_X1   g205(.A(G1341), .B(G1348), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n628), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2443), .B(G2446), .Z(new_n634));
  OAI21_X1  g209(.A(G14), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n633), .ZN(G401));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2072), .B(G2078), .Z(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT18), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(KEYINPUT17), .ZN(new_n643));
  INV_X1    g218(.A(new_n637), .ZN(new_n644));
  INV_X1    g219(.A(new_n638), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n640), .A3(new_n645), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(new_n639), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n642), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT84), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(G227));
  XNOR2_X1  g227(.A(G1991), .B(G1996), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT88), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  AND2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n660), .A2(new_n661), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  MUX2_X1   g242(.A(new_n667), .B(new_n666), .S(new_n659), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT85), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1981), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G1986), .ZN(new_n672));
  INV_X1    g247(.A(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(G1986), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  AND3_X1   g253(.A1(new_n672), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n678), .B1(new_n672), .B2(new_n676), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n657), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n674), .A2(new_n675), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n671), .A2(G1986), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n677), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n672), .A2(new_n676), .A3(new_n678), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(new_n656), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(new_n686), .ZN(G229));
  NAND2_X1  g262(.A1(new_n573), .A2(G16), .ZN(new_n688));
  OR2_X1    g263(.A1(G6), .A2(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(KEYINPUT32), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT32), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n688), .A2(new_n692), .A3(new_n689), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1981), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n696));
  NAND2_X1  g271(.A1(G303), .A2(G16), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G22), .ZN(new_n700));
  AND3_X1   g275(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n698), .B1(new_n697), .B2(new_n700), .ZN(new_n702));
  MUX2_X1   g277(.A(G23), .B(G288), .S(G16), .Z(new_n703));
  XOR2_X1   g278(.A(KEYINPUT33), .B(G1976), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NOR3_X1   g280(.A1(new_n701), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n695), .A2(new_n696), .A3(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(G16), .A2(G24), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G290), .B2(new_n699), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(new_n675), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G25), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n467), .A2(G107), .ZN(new_n713));
  OAI21_X1  g288(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n483), .A2(G119), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n480), .A2(G131), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n712), .B1(new_n719), .B2(new_n711), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT35), .B(G1991), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n709), .A2(new_n675), .ZN(new_n723));
  AND4_X1   g298(.A1(new_n707), .A2(new_n710), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n695), .A2(new_n706), .ZN(new_n725));
  AOI21_X1  g300(.A(KEYINPUT89), .B1(new_n725), .B2(KEYINPUT34), .ZN(new_n726));
  AND3_X1   g301(.A1(new_n725), .A2(KEYINPUT89), .A3(KEYINPUT34), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(KEYINPUT90), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n724), .B(new_n730), .C1(new_n726), .C2(new_n727), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n729), .A2(KEYINPUT36), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G171), .A2(new_n699), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G5), .B2(new_n699), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G19), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n548), .B2(G16), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n734), .A2(new_n735), .B1(G1341), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n711), .A2(G27), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G164), .B2(new_n711), .ZN(new_n740));
  OAI221_X1 g315(.A(new_n738), .B1(G1341), .B2(new_n737), .C1(G2078), .C2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT24), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(G34), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(G34), .ZN(new_n745));
  AOI21_X1  g320(.A(G29), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G160), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(G29), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n711), .A2(G33), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT25), .Z(new_n752));
  INV_X1    g327(.A(G139), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n752), .B1(new_n753), .B2(new_n468), .C1(new_n467), .C2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n750), .B1(new_n755), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2072), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n749), .A2(G2084), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT92), .B(G2067), .Z(new_n759));
  AND3_X1   g334(.A1(new_n711), .A2(KEYINPUT28), .A3(G26), .ZN(new_n760));
  AOI21_X1  g335(.A(KEYINPUT28), .B1(new_n711), .B2(G26), .ZN(new_n761));
  NOR2_X1   g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT91), .Z(new_n763));
  OAI211_X1 g338(.A(new_n763), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n480), .A2(G140), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n483), .A2(G128), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n760), .B(new_n761), .C1(new_n767), .C2(G29), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI221_X1 g344(.A(new_n758), .B1(new_n759), .B2(new_n769), .C1(new_n734), .C2(new_n735), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT30), .B(G28), .ZN(new_n771));
  OR2_X1    g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  NAND2_X1  g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n771), .A2(new_n711), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n620), .B2(new_n711), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n769), .B2(new_n759), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n776), .B1(new_n757), .B2(new_n756), .C1(G2084), .C2(new_n749), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n741), .A2(new_n770), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n699), .A2(G20), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT23), .Z(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G299), .B2(G16), .ZN(new_n781));
  INV_X1    g356(.A(G1956), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n711), .A2(G35), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G162), .B2(new_n711), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT29), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(G2090), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(G2090), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n740), .A2(G2078), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n783), .A2(new_n787), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G16), .A2(G21), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G168), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1966), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n711), .A2(G32), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n480), .A2(G141), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n483), .A2(G129), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n606), .A2(G105), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT26), .Z(new_n800));
  NAND4_X1  g375(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n795), .B1(new_n802), .B2(new_n711), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT27), .B(G1996), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n592), .A2(G16), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G4), .B2(G16), .ZN(new_n807));
  INV_X1    g382(.A(G1348), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n808), .B2(new_n807), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n778), .A2(new_n790), .A3(new_n794), .A4(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT93), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n732), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(KEYINPUT36), .B1(new_n729), .B2(new_n731), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(G311));
  INV_X1    g390(.A(new_n814), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n816), .A2(new_n812), .A3(new_n732), .ZN(G150));
  XNOR2_X1  g392(.A(KEYINPUT97), .B(G860), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n592), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT95), .B(G93), .Z(new_n822));
  AOI22_X1  g397(.A1(G55), .A2(new_n512), .B1(new_n515), .B2(new_n822), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  OR3_X1    g399(.A1(new_n824), .A2(KEYINPUT94), .A3(new_n518), .ZN(new_n825));
  OAI21_X1  g400(.A(KEYINPUT94), .B1(new_n824), .B2(new_n518), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(KEYINPUT96), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(KEYINPUT96), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n828), .A2(new_n547), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n548), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n821), .B(new_n832), .Z(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n819), .B1(new_n834), .B2(KEYINPUT39), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(KEYINPUT39), .B2(new_n834), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n828), .A2(new_n829), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n819), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(G145));
  XNOR2_X1  g415(.A(G164), .B(new_n767), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n802), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(new_n755), .Z(new_n843));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n480), .A2(G142), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n483), .A2(G130), .ZN(new_n846));
  OR2_X1    g421(.A1(G106), .A2(G2105), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n847), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n719), .A2(KEYINPUT99), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n718), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n608), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n853), .A2(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n849), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n856), .A2(new_n849), .A3(new_n857), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n843), .B1(new_n844), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n858), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n842), .B(new_n755), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT101), .ZN(new_n866));
  XNOR2_X1  g441(.A(G160), .B(KEYINPUT98), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G162), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n867), .A2(G162), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n620), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  INV_X1    g447(.A(new_n620), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n873), .A3(new_n868), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT102), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n862), .A2(new_n866), .A3(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT100), .B(G37), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n843), .A2(new_n861), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n864), .A2(new_n865), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT103), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n877), .A4(new_n878), .ZN(new_n886));
  XNOR2_X1  g461(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n887), .B1(new_n883), .B2(new_n886), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(G395));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n891));
  NAND2_X1  g466(.A1(G299), .A2(new_n592), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n591), .A2(new_n556), .A3(new_n560), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT41), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n894), .A2(KEYINPUT106), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(KEYINPUT106), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n892), .A2(KEYINPUT105), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(KEYINPUT105), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n893), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n895), .B(new_n896), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n832), .B(new_n602), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n899), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n907));
  XOR2_X1   g482(.A(G290), .B(G288), .Z(new_n908));
  NAND2_X1  g483(.A1(G303), .A2(G305), .ZN(new_n909));
  NAND2_X1  g484(.A1(G166), .A2(new_n573), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n909), .A2(new_n910), .ZN(new_n914));
  INV_X1    g489(.A(new_n908), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT107), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(KEYINPUT109), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n903), .A2(new_n905), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n907), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(G868), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n922), .B1(new_n907), .B2(new_n924), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n891), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n927), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n929), .A2(KEYINPUT110), .A3(G868), .A4(new_n925), .ZN(new_n930));
  INV_X1    g505(.A(new_n837), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n928), .B(new_n930), .C1(G868), .C2(new_n931), .ZN(G295));
  OAI211_X1 g507(.A(new_n928), .B(new_n930), .C1(G868), .C2(new_n931), .ZN(G331));
  NAND2_X1  g508(.A1(new_n921), .A2(KEYINPUT111), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n830), .A2(new_n831), .A3(G168), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(G168), .B1(new_n830), .B2(new_n831), .ZN(new_n937));
  OAI21_X1  g512(.A(G301), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n937), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(G171), .A3(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n904), .B1(new_n941), .B2(new_n900), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n913), .A2(new_n920), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n892), .A2(new_n893), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n938), .A2(new_n940), .A3(KEYINPUT41), .A4(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n934), .A2(new_n942), .A3(new_n944), .A4(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n901), .A2(new_n940), .A3(new_n938), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n941), .A2(new_n899), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n921), .ZN(new_n950));
  AND4_X1   g525(.A1(KEYINPUT43), .A2(new_n947), .A3(new_n878), .A4(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G37), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n948), .A2(new_n949), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n954), .A2(new_n934), .A3(new_n944), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT43), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n947), .A2(new_n958), .A3(new_n878), .A4(new_n950), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n958), .B1(new_n953), .B2(new_n955), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n957), .B1(new_n962), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT4), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(new_n498), .B2(new_n499), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n966), .A2(new_n502), .B1(new_n476), .B2(new_n504), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n964), .B1(new_n967), .B2(new_n493), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(G160), .A2(G40), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n767), .B(G2067), .Z(new_n974));
  INV_X1    g549(.A(G1996), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n801), .B(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n721), .A3(new_n719), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n767), .A2(G2067), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n973), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OR3_X1    g555(.A1(new_n973), .A2(G1986), .A3(G290), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n718), .B(new_n721), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n977), .A2(new_n984), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n981), .A2(new_n982), .B1(new_n972), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n980), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT46), .B1(new_n972), .B2(new_n975), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n988), .B(KEYINPUT127), .Z(new_n989));
  AOI21_X1  g564(.A(new_n801), .B1(KEYINPUT46), .B2(new_n975), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n974), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n973), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n993), .B2(new_n992), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(G164), .B2(G1384), .ZN(new_n997));
  AND2_X1   g572(.A1(G160), .A2(G40), .ZN(new_n998));
  OAI211_X1 g573(.A(KEYINPUT112), .B(new_n964), .C1(new_n967), .C2(new_n493), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n1000), .A2(G8), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT115), .B(G1981), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n573), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n512), .A2(G48), .ZN(new_n1004));
  INV_X1    g579(.A(new_n515), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT116), .B(G86), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n569), .B(new_n1004), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G1981), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1003), .A2(KEYINPUT49), .A3(new_n1008), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1001), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1976), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G288), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT114), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1001), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(G288), .B2(new_n1014), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1013), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(KEYINPUT52), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n997), .A2(new_n1024), .A3(new_n999), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n971), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G2090), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(KEYINPUT45), .B(new_n964), .C1(new_n967), .C2(new_n493), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1030), .A2(new_n998), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n970), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n698), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1023), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(G166), .B2(new_n1023), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n522), .A2(KEYINPUT55), .A3(G8), .A4(new_n523), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1035), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1035), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1034), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OR2_X1    g620(.A1(G288), .A2(G1976), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1003), .B1(new_n1013), .B2(new_n1046), .ZN(new_n1047));
  XOR2_X1   g622(.A(new_n1001), .B(KEYINPUT117), .Z(new_n1048));
  AOI22_X1  g623(.A1(new_n1022), .A2(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT120), .B(KEYINPUT63), .Z(new_n1050));
  NAND3_X1  g625(.A1(new_n1044), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n997), .A2(new_n999), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT50), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n998), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n1028), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1033), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1041), .B1(new_n1057), .B2(G8), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1051), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1030), .A2(new_n998), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n1052), .B2(new_n969), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT118), .B1(new_n1061), .B2(G1966), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT45), .B1(new_n997), .B2(new_n999), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1063), .B(new_n793), .C1(new_n1064), .C2(new_n1060), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT119), .B(G2084), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1027), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1023), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G168), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1050), .B1(new_n1059), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1042), .B1(new_n1034), .B2(KEYINPUT121), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(KEYINPUT121), .B2(new_n1034), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1044), .A2(new_n1020), .A3(KEYINPUT63), .A4(new_n1021), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1070), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1049), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1059), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n534), .A2(G8), .A3(new_n535), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1079), .A2(KEYINPUT123), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(KEYINPUT123), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1069), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1080), .A2(KEYINPUT124), .A3(new_n1081), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT51), .B1(new_n1069), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1086), .B1(new_n1091), .B2(KEYINPUT125), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT125), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1093), .B(KEYINPUT51), .C1(new_n1069), .C2(new_n1090), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1084), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G2078), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1061), .A2(KEYINPUT53), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1032), .B2(G2078), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n735), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1078), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1091), .A2(KEYINPUT125), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1086), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1094), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1084), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1102), .A2(G171), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(KEYINPUT62), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n1112));
  XNOR2_X1  g687(.A(G299), .B(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1024), .B1(new_n997), .B2(new_n999), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n782), .B1(new_n1114), .B2(new_n1054), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1031), .A2(new_n970), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(G1348), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1000), .A2(G2067), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(new_n591), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1113), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1118), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1118), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(new_n1123), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n970), .A2(new_n975), .A3(new_n998), .A4(new_n1030), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT58), .B(G1341), .Z(new_n1131));
  NAND2_X1  g706(.A1(new_n1000), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n548), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1121), .A2(KEYINPUT60), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n592), .A3(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(G299), .B(KEYINPUT57), .ZN(new_n1142));
  AOI21_X1  g717(.A(G1956), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1031), .A2(new_n970), .A3(new_n1116), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(KEYINPUT61), .A3(new_n1118), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1127), .A2(new_n1137), .A3(new_n1141), .A4(new_n1146), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1135), .A2(new_n1136), .B1(new_n1138), .B2(new_n592), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1124), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1096), .A2(KEYINPUT53), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1099), .B(new_n1101), .C1(new_n1150), .C2(new_n1032), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1110), .B1(G171), .B2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT126), .B(KEYINPUT54), .Z(new_n1153));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1151), .B2(G171), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1102), .A2(G171), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1152), .A2(new_n1153), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1111), .B1(new_n1149), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1109), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1077), .B1(new_n1104), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n985), .ZN(new_n1161));
  XNOR2_X1  g736(.A(G290), .B(new_n675), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n973), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n995), .B1(new_n1160), .B2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g739(.A(G319), .ZN(new_n1166));
  NOR3_X1   g740(.A1(G227), .A2(new_n1166), .A3(G401), .ZN(new_n1167));
  NAND3_X1  g741(.A1(new_n681), .A2(new_n686), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g742(.A1(new_n953), .A2(new_n955), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n1169), .A2(KEYINPUT43), .ZN(new_n1170));
  AOI221_X4 g744(.A(new_n1168), .B1(new_n883), .B2(new_n886), .C1(new_n1170), .C2(new_n959), .ZN(G308));
  AOI21_X1  g745(.A(new_n1168), .B1(new_n883), .B2(new_n886), .ZN(new_n1172));
  OAI21_X1  g746(.A(new_n1172), .B1(new_n961), .B2(new_n960), .ZN(G225));
endmodule


