

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721;

  XNOR2_X1 U371 ( .A(n349), .B(n348), .ZN(G63) );
  INV_X1 U372 ( .A(KEYINPUT120), .ZN(n348) );
  NOR2_X1 U373 ( .A1(n706), .A2(n611), .ZN(n610) );
  XNOR2_X1 U374 ( .A(n351), .B(n350), .ZN(n717) );
  INV_X1 U375 ( .A(n499), .ZN(n350) );
  XNOR2_X1 U376 ( .A(n352), .B(KEYINPUT103), .ZN(n462) );
  OR2_X1 U377 ( .A1(n484), .A2(n513), .ZN(n352) );
  NOR2_X1 U378 ( .A1(G902), .A2(n685), .ZN(n436) );
  XNOR2_X1 U379 ( .A(n362), .B(G119), .ZN(n364) );
  XNOR2_X1 U380 ( .A(G116), .B(G113), .ZN(n363) );
  NAND2_X1 U381 ( .A1(n680), .A2(n681), .ZN(n349) );
  XNOR2_X2 U382 ( .A(n377), .B(n376), .ZN(n514) );
  NAND2_X1 U383 ( .A1(n498), .A2(n516), .ZN(n351) );
  INV_X1 U384 ( .A(G953), .ZN(n707) );
  XOR2_X2 U385 ( .A(n473), .B(KEYINPUT1), .Z(n563) );
  INV_X2 U386 ( .A(KEYINPUT3), .ZN(n362) );
  NOR2_X2 U387 ( .A1(n574), .A2(n560), .ZN(n561) );
  XNOR2_X2 U388 ( .A(n557), .B(n556), .ZN(n574) );
  XNOR2_X2 U389 ( .A(n494), .B(KEYINPUT6), .ZN(n573) );
  XNOR2_X2 U390 ( .A(n463), .B(KEYINPUT41), .ZN(n498) );
  XNOR2_X1 U391 ( .A(n551), .B(n355), .ZN(n568) );
  XOR2_X2 U392 ( .A(G137), .B(G140), .Z(n428) );
  XNOR2_X1 U393 ( .A(n677), .B(KEYINPUT119), .ZN(n678) );
  XNOR2_X1 U394 ( .A(KEYINPUT16), .B(G122), .ZN(n365) );
  XNOR2_X1 U395 ( .A(G143), .B(G128), .ZN(n382) );
  XNOR2_X1 U396 ( .A(n694), .B(n367), .ZN(n371) );
  XNOR2_X1 U397 ( .A(n451), .B(n450), .ZN(n547) );
  XNOR2_X1 U398 ( .A(KEYINPUT85), .B(KEYINPUT33), .ZN(n450) );
  XNOR2_X1 U399 ( .A(n401), .B(n400), .ZN(n618) );
  XNOR2_X1 U400 ( .A(n693), .B(n361), .ZN(n414) );
  XNOR2_X1 U401 ( .A(n441), .B(KEYINPUT70), .ZN(n361) );
  XOR2_X1 U402 ( .A(KEYINPUT89), .B(n428), .Z(n702) );
  XNOR2_X1 U403 ( .A(n434), .B(KEYINPUT25), .ZN(n435) );
  NOR2_X1 U404 ( .A1(n582), .A2(n473), .ZN(n474) );
  XNOR2_X1 U405 ( .A(n356), .B(n372), .ZN(n625) );
  XNOR2_X1 U406 ( .A(n371), .B(n370), .ZN(n356) );
  XNOR2_X1 U407 ( .A(KEYINPUT65), .B(KEYINPUT0), .ZN(n545) );
  XNOR2_X1 U408 ( .A(n432), .B(n431), .ZN(n685) );
  XNOR2_X1 U409 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U410 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U411 ( .A(n702), .B(n357), .ZN(n413) );
  INV_X1 U412 ( .A(KEYINPUT35), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n568), .B(G122), .ZN(G24) );
  NAND2_X1 U414 ( .A1(n555), .A2(n354), .ZN(n556) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n586) );
  INV_X1 U416 ( .A(KEYINPUT88), .ZN(n353) );
  NAND2_X1 U417 ( .A1(n579), .A2(n354), .ZN(n580) );
  XNOR2_X2 U418 ( .A(n546), .B(n545), .ZN(n354) );
  NAND2_X1 U419 ( .A1(n625), .A2(n611), .ZN(n377) );
  XNOR2_X1 U420 ( .A(n620), .B(n619), .ZN(n622) );
  XNOR2_X1 U421 ( .A(n426), .B(n425), .ZN(n432) );
  XNOR2_X1 U422 ( .A(n390), .B(n366), .ZN(n367) );
  XNOR2_X2 U423 ( .A(n364), .B(n363), .ZN(n440) );
  AND2_X1 U424 ( .A1(G227), .A2(n707), .ZN(n357) );
  XOR2_X1 U425 ( .A(G104), .B(G107), .Z(n358) );
  INV_X1 U426 ( .A(n651), .ZN(n566) );
  NOR2_X1 U427 ( .A1(n571), .A2(n582), .ZN(n458) );
  XNOR2_X1 U428 ( .A(n399), .B(n398), .ZN(n400) );
  NOR2_X1 U429 ( .A1(n406), .A2(n520), .ZN(n552) );
  NOR2_X1 U430 ( .A1(n536), .A2(n534), .ZN(n509) );
  XNOR2_X1 U431 ( .A(n424), .B(KEYINPUT24), .ZN(n425) );
  AND2_X2 U432 ( .A1(n616), .A2(n615), .ZN(n676) );
  BUF_X1 U433 ( .A(n676), .Z(n683) );
  BUF_X1 U434 ( .A(n514), .Z(n536) );
  NOR2_X2 U435 ( .A1(n622), .A2(n687), .ZN(n624) );
  XNOR2_X1 U436 ( .A(n608), .B(n607), .ZN(G75) );
  XNOR2_X1 U437 ( .A(KEYINPUT74), .B(G110), .ZN(n359) );
  XNOR2_X1 U438 ( .A(n358), .B(n359), .ZN(n693) );
  INV_X1 U439 ( .A(KEYINPUT4), .ZN(n360) );
  XNOR2_X1 U440 ( .A(n360), .B(G101), .ZN(n441) );
  XNOR2_X1 U441 ( .A(n414), .B(KEYINPUT75), .ZN(n372) );
  XNOR2_X2 U442 ( .A(n440), .B(n365), .ZN(n694) );
  XOR2_X2 U443 ( .A(G146), .B(G125), .Z(n390) );
  XOR2_X1 U444 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n366) );
  NAND2_X1 U445 ( .A1(G224), .A2(n707), .ZN(n368) );
  XNOR2_X1 U446 ( .A(n368), .B(KEYINPUT86), .ZN(n369) );
  XOR2_X1 U447 ( .A(n369), .B(n382), .Z(n370) );
  XNOR2_X1 U448 ( .A(G902), .B(KEYINPUT15), .ZN(n611) );
  XOR2_X1 U449 ( .A(KEYINPUT87), .B(KEYINPUT77), .Z(n375) );
  INV_X1 U450 ( .A(G902), .ZN(n416) );
  INV_X1 U451 ( .A(G237), .ZN(n373) );
  NAND2_X1 U452 ( .A1(n416), .A2(n373), .ZN(n379) );
  NAND2_X1 U453 ( .A1(G210), .A2(n379), .ZN(n374) );
  XOR2_X1 U454 ( .A(n375), .B(n374), .Z(n376) );
  INV_X1 U455 ( .A(KEYINPUT38), .ZN(n378) );
  XNOR2_X1 U456 ( .A(n514), .B(n378), .ZN(n484) );
  NAND2_X1 U457 ( .A1(n379), .A2(G214), .ZN(n507) );
  INV_X1 U458 ( .A(n507), .ZN(n513) );
  NAND2_X1 U459 ( .A1(n484), .A2(n513), .ZN(n407) );
  XNOR2_X1 U460 ( .A(G116), .B(G107), .ZN(n380) );
  XNOR2_X1 U461 ( .A(n380), .B(KEYINPUT9), .ZN(n381) );
  XOR2_X1 U462 ( .A(n381), .B(KEYINPUT7), .Z(n384) );
  XNOR2_X1 U463 ( .A(n382), .B(G134), .ZN(n412) );
  XNOR2_X1 U464 ( .A(n412), .B(G122), .ZN(n383) );
  XNOR2_X1 U465 ( .A(n384), .B(n383), .ZN(n388) );
  NAND2_X1 U466 ( .A1(G234), .A2(n707), .ZN(n386) );
  XOR2_X1 U467 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n385) );
  XNOR2_X1 U468 ( .A(n386), .B(n385), .ZN(n427) );
  NAND2_X1 U469 ( .A1(G217), .A2(n427), .ZN(n387) );
  XOR2_X1 U470 ( .A(n388), .B(n387), .Z(n677) );
  NOR2_X1 U471 ( .A1(G902), .A2(n677), .ZN(n389) );
  XNOR2_X1 U472 ( .A(n389), .B(G478), .ZN(n522) );
  INV_X1 U473 ( .A(n522), .ZN(n406) );
  XNOR2_X1 U474 ( .A(KEYINPUT13), .B(KEYINPUT95), .ZN(n403) );
  XOR2_X2 U475 ( .A(KEYINPUT10), .B(n390), .Z(n701) );
  XOR2_X1 U476 ( .A(n701), .B(G104), .Z(n401) );
  XOR2_X1 U477 ( .A(KEYINPUT12), .B(G122), .Z(n392) );
  XNOR2_X1 U478 ( .A(G113), .B(G140), .ZN(n391) );
  XNOR2_X1 U479 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U480 ( .A(KEYINPUT94), .B(KEYINPUT11), .Z(n394) );
  NOR2_X1 U481 ( .A1(G953), .A2(G237), .ZN(n437) );
  NAND2_X1 U482 ( .A1(G214), .A2(n437), .ZN(n393) );
  XNOR2_X1 U483 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U484 ( .A(n396), .B(n395), .ZN(n399) );
  INV_X1 U485 ( .A(KEYINPUT67), .ZN(n397) );
  XNOR2_X1 U486 ( .A(n397), .B(G131), .ZN(n411) );
  XNOR2_X1 U487 ( .A(n411), .B(G143), .ZN(n398) );
  NOR2_X1 U488 ( .A1(G902), .A2(n618), .ZN(n402) );
  XNOR2_X1 U489 ( .A(n403), .B(n402), .ZN(n405) );
  INV_X1 U490 ( .A(G475), .ZN(n404) );
  XNOR2_X1 U491 ( .A(n405), .B(n404), .ZN(n520) );
  NAND2_X1 U492 ( .A1(n407), .A2(n552), .ZN(n410) );
  NAND2_X1 U493 ( .A1(n520), .A2(n522), .ZN(n657) );
  OR2_X1 U494 ( .A1(n520), .A2(n522), .ZN(n653) );
  XNOR2_X1 U495 ( .A(n653), .B(KEYINPUT96), .ZN(n531) );
  NAND2_X1 U496 ( .A1(n657), .A2(n531), .ZN(n517) );
  NAND2_X1 U497 ( .A1(n462), .A2(n517), .ZN(n409) );
  NAND2_X1 U498 ( .A1(n410), .A2(n409), .ZN(n452) );
  XNOR2_X1 U499 ( .A(n412), .B(n411), .ZN(n705) );
  XNOR2_X1 U500 ( .A(n705), .B(G146), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U502 ( .A(n446), .B(n415), .ZN(n672) );
  NAND2_X1 U503 ( .A1(n672), .A2(n416), .ZN(n418) );
  XOR2_X1 U504 ( .A(KEYINPUT68), .B(G469), .Z(n417) );
  XNOR2_X2 U505 ( .A(n418), .B(n417), .ZN(n473) );
  INV_X1 U506 ( .A(n563), .ZN(n571) );
  XOR2_X1 U507 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n420) );
  NAND2_X1 U508 ( .A1(G234), .A2(n611), .ZN(n419) );
  XNOR2_X1 U509 ( .A(n420), .B(n419), .ZN(n433) );
  NAND2_X1 U510 ( .A1(n433), .A2(G221), .ZN(n421) );
  XOR2_X1 U511 ( .A(KEYINPUT21), .B(n421), .Z(n489) );
  XNOR2_X1 U512 ( .A(KEYINPUT92), .B(n489), .ZN(n553) );
  XNOR2_X1 U513 ( .A(n701), .B(KEYINPUT90), .ZN(n426) );
  XOR2_X1 U514 ( .A(KEYINPUT23), .B(G110), .Z(n423) );
  XNOR2_X1 U515 ( .A(G119), .B(G128), .ZN(n422) );
  XOR2_X1 U516 ( .A(n423), .B(n422), .Z(n424) );
  NAND2_X1 U517 ( .A1(n427), .A2(G221), .ZN(n430) );
  XNOR2_X1 U518 ( .A(n428), .B(KEYINPUT69), .ZN(n429) );
  NAND2_X1 U519 ( .A1(G217), .A2(n433), .ZN(n434) );
  XNOR2_X2 U520 ( .A(n436), .B(n435), .ZN(n562) );
  NAND2_X1 U521 ( .A1(n553), .A2(n562), .ZN(n582) );
  NAND2_X1 U522 ( .A1(n437), .A2(G210), .ZN(n438) );
  XNOR2_X1 U523 ( .A(n438), .B(KEYINPUT93), .ZN(n439) );
  XNOR2_X1 U524 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U525 ( .A(G137), .B(KEYINPUT5), .Z(n442) );
  XNOR2_X1 U526 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U527 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U528 ( .A(n446), .B(n445), .ZN(n637) );
  OR2_X1 U529 ( .A1(n637), .A2(G902), .ZN(n449) );
  INV_X1 U530 ( .A(KEYINPUT72), .ZN(n447) );
  XNOR2_X1 U531 ( .A(n447), .B(G472), .ZN(n448) );
  XNOR2_X2 U532 ( .A(n449), .B(n448), .ZN(n494) );
  NAND2_X1 U533 ( .A1(n458), .A2(n573), .ZN(n451) );
  INV_X1 U534 ( .A(n547), .ZN(n602) );
  NAND2_X1 U535 ( .A1(n452), .A2(n602), .ZN(n466) );
  AND2_X1 U536 ( .A1(n571), .A2(n582), .ZN(n453) );
  XNOR2_X1 U537 ( .A(n453), .B(KEYINPUT50), .ZN(n454) );
  INV_X1 U538 ( .A(n494), .ZN(n581) );
  NOR2_X1 U539 ( .A1(n454), .A2(n581), .ZN(n457) );
  XNOR2_X1 U540 ( .A(KEYINPUT98), .B(n562), .ZN(n572) );
  NOR2_X1 U541 ( .A1(n572), .A2(n489), .ZN(n455) );
  XNOR2_X1 U542 ( .A(n455), .B(KEYINPUT49), .ZN(n456) );
  NAND2_X1 U543 ( .A1(n457), .A2(n456), .ZN(n460) );
  INV_X1 U544 ( .A(n458), .ZN(n459) );
  OR2_X1 U545 ( .A1(n494), .A2(n459), .ZN(n578) );
  AND2_X1 U546 ( .A1(n460), .A2(n578), .ZN(n461) );
  XNOR2_X1 U547 ( .A(KEYINPUT51), .B(n461), .ZN(n464) );
  NAND2_X1 U548 ( .A1(n462), .A2(n552), .ZN(n463) );
  NAND2_X1 U549 ( .A1(n464), .A2(n498), .ZN(n465) );
  NAND2_X1 U550 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U551 ( .A(n467), .B(KEYINPUT115), .ZN(n468) );
  XNOR2_X1 U552 ( .A(KEYINPUT52), .B(n468), .ZN(n471) );
  NAND2_X1 U553 ( .A1(G234), .A2(G237), .ZN(n469) );
  XNOR2_X1 U554 ( .A(n469), .B(KEYINPUT14), .ZN(n477) );
  NAND2_X1 U555 ( .A1(G952), .A2(n477), .ZN(n470) );
  NOR2_X1 U556 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U557 ( .A1(G953), .A2(n472), .ZN(n606) );
  XNOR2_X1 U558 ( .A(n474), .B(KEYINPUT100), .ZN(n483) );
  OR2_X1 U559 ( .A1(n494), .A2(n513), .ZN(n475) );
  XNOR2_X1 U560 ( .A(n475), .B(KEYINPUT30), .ZN(n481) );
  OR2_X1 U561 ( .A1(n707), .A2(G902), .ZN(n476) );
  NAND2_X1 U562 ( .A1(n477), .A2(n476), .ZN(n479) );
  NOR2_X1 U563 ( .A1(G953), .A2(G952), .ZN(n478) );
  NOR2_X1 U564 ( .A1(n479), .A2(n478), .ZN(n542) );
  NAND2_X1 U565 ( .A1(G953), .A2(G900), .ZN(n480) );
  NAND2_X1 U566 ( .A1(n542), .A2(n480), .ZN(n490) );
  NOR2_X1 U567 ( .A1(n481), .A2(n490), .ZN(n482) );
  NAND2_X1 U568 ( .A1(n483), .A2(n482), .ZN(n519) );
  OR2_X1 U569 ( .A1(n519), .A2(n484), .ZN(n485) );
  XNOR2_X2 U570 ( .A(n485), .B(KEYINPUT39), .ZN(n533) );
  INV_X1 U571 ( .A(n657), .ZN(n660) );
  NAND2_X1 U572 ( .A1(n533), .A2(n660), .ZN(n488) );
  INV_X1 U573 ( .A(KEYINPUT102), .ZN(n486) );
  XNOR2_X1 U574 ( .A(n486), .B(KEYINPUT40), .ZN(n487) );
  XNOR2_X1 U575 ( .A(n488), .B(n487), .ZN(n635) );
  INV_X1 U576 ( .A(n562), .ZN(n493) );
  INV_X1 U577 ( .A(n489), .ZN(n491) );
  NOR2_X1 U578 ( .A1(n491), .A2(n490), .ZN(n492) );
  NAND2_X1 U579 ( .A1(n493), .A2(n492), .ZN(n504) );
  NOR2_X1 U580 ( .A1(n504), .A2(n494), .ZN(n495) );
  XNOR2_X1 U581 ( .A(n495), .B(KEYINPUT28), .ZN(n497) );
  XNOR2_X1 U582 ( .A(n473), .B(KEYINPUT101), .ZN(n496) );
  AND2_X1 U583 ( .A1(n497), .A2(n496), .ZN(n516) );
  XNOR2_X1 U584 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n499) );
  NOR2_X2 U585 ( .A1(n635), .A2(n717), .ZN(n502) );
  XNOR2_X1 U586 ( .A(KEYINPUT82), .B(KEYINPUT46), .ZN(n501) );
  XNOR2_X1 U587 ( .A(n502), .B(n501), .ZN(n529) );
  INV_X1 U588 ( .A(n573), .ZN(n503) );
  NOR2_X1 U589 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U590 ( .A(n505), .B(KEYINPUT99), .ZN(n506) );
  NOR2_X1 U591 ( .A1(n657), .A2(n506), .ZN(n508) );
  NAND2_X1 U592 ( .A1(n508), .A2(n507), .ZN(n534) );
  XNOR2_X1 U593 ( .A(KEYINPUT36), .B(n509), .ZN(n510) );
  AND2_X1 U594 ( .A1(n510), .A2(n563), .ZN(n512) );
  INV_X1 U595 ( .A(KEYINPUT105), .ZN(n511) );
  XNOR2_X1 U596 ( .A(n512), .B(n511), .ZN(n718) );
  OR2_X2 U597 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X2 U598 ( .A(n515), .B(KEYINPUT19), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n544), .A2(n516), .ZN(n656) );
  INV_X1 U600 ( .A(n517), .ZN(n588) );
  NOR2_X1 U601 ( .A1(n656), .A2(n588), .ZN(n518) );
  XNOR2_X1 U602 ( .A(n518), .B(KEYINPUT47), .ZN(n526) );
  INV_X1 U603 ( .A(n519), .ZN(n525) );
  INV_X1 U604 ( .A(n520), .ZN(n521) );
  NOR2_X1 U605 ( .A1(n522), .A2(n521), .ZN(n549) );
  INV_X1 U606 ( .A(n549), .ZN(n523) );
  NOR2_X1 U607 ( .A1(n536), .A2(n523), .ZN(n524) );
  NAND2_X1 U608 ( .A1(n525), .A2(n524), .ZN(n633) );
  NAND2_X1 U609 ( .A1(n526), .A2(n633), .ZN(n527) );
  NOR2_X1 U610 ( .A1(n718), .A2(n527), .ZN(n528) );
  NAND2_X1 U611 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U612 ( .A(n530), .B(KEYINPUT48), .ZN(n539) );
  INV_X1 U613 ( .A(n531), .ZN(n532) );
  NAND2_X1 U614 ( .A1(n533), .A2(n532), .ZN(n667) );
  OR2_X1 U615 ( .A1(n534), .A2(n563), .ZN(n535) );
  XNOR2_X1 U616 ( .A(n535), .B(KEYINPUT43), .ZN(n537) );
  NAND2_X1 U617 ( .A1(n537), .A2(n536), .ZN(n669) );
  NAND2_X1 U618 ( .A1(n667), .A2(n669), .ZN(n538) );
  NOR2_X2 U619 ( .A1(n539), .A2(n538), .ZN(n609) );
  NOR2_X1 U620 ( .A1(n609), .A2(KEYINPUT2), .ZN(n540) );
  XNOR2_X1 U621 ( .A(n540), .B(KEYINPUT78), .ZN(n596) );
  NAND2_X1 U622 ( .A1(G898), .A2(G953), .ZN(n541) );
  AND2_X1 U623 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U624 ( .A1(n544), .A2(n543), .ZN(n546) );
  NOR2_X1 U625 ( .A1(n547), .A2(n586), .ZN(n548) );
  XNOR2_X1 U626 ( .A(n548), .B(KEYINPUT34), .ZN(n550) );
  NAND2_X1 U627 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U628 ( .A(KEYINPUT22), .B(KEYINPUT73), .Z(n557) );
  NAND2_X1 U629 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U630 ( .A(KEYINPUT97), .B(n554), .ZN(n555) );
  OR2_X1 U631 ( .A1(n572), .A2(n573), .ZN(n558) );
  NOR2_X1 U632 ( .A1(n571), .A2(n558), .ZN(n559) );
  XOR2_X1 U633 ( .A(KEYINPUT76), .B(n559), .Z(n560) );
  XOR2_X1 U634 ( .A(KEYINPUT32), .B(n561), .Z(n720) );
  NOR2_X1 U635 ( .A1(n574), .A2(n562), .ZN(n565) );
  NOR2_X1 U636 ( .A1(n563), .A2(n581), .ZN(n564) );
  AND2_X1 U637 ( .A1(n565), .A2(n564), .ZN(n651) );
  AND2_X1 U638 ( .A1(n720), .A2(n566), .ZN(n567) );
  NAND2_X1 U639 ( .A1(n568), .A2(n567), .ZN(n570) );
  NOR2_X1 U640 ( .A1(KEYINPUT71), .A2(KEYINPUT44), .ZN(n569) );
  XNOR2_X1 U641 ( .A(n570), .B(n569), .ZN(n593) );
  NAND2_X1 U642 ( .A1(KEYINPUT71), .A2(KEYINPUT44), .ZN(n591) );
  NAND2_X1 U643 ( .A1(n572), .A2(n571), .ZN(n577) );
  NOR2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U645 ( .A(n575), .B(KEYINPUT83), .ZN(n576) );
  NOR2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n643) );
  INV_X1 U647 ( .A(n578), .ZN(n579) );
  XNOR2_X1 U648 ( .A(n580), .B(KEYINPUT31), .ZN(n664) );
  NOR2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n584) );
  INV_X1 U650 ( .A(n473), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n645) );
  NOR2_X1 U653 ( .A1(n664), .A2(n645), .ZN(n587) );
  NOR2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U655 ( .A1(n643), .A2(n589), .ZN(n590) );
  AND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X2 U658 ( .A(n594), .B(KEYINPUT45), .ZN(n688) );
  NOR2_X1 U659 ( .A1(n688), .A2(KEYINPUT2), .ZN(n595) );
  NOR2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U661 ( .A1(n609), .A2(KEYINPUT2), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n597), .B(KEYINPUT81), .ZN(n598) );
  NAND2_X1 U663 ( .A1(n688), .A2(n598), .ZN(n615) );
  AND2_X1 U664 ( .A1(n599), .A2(n615), .ZN(n601) );
  INV_X1 U665 ( .A(KEYINPUT79), .ZN(n600) );
  XNOR2_X1 U666 ( .A(n601), .B(n600), .ZN(n604) );
  AND2_X1 U667 ( .A1(n498), .A2(n602), .ZN(n603) );
  NOR2_X1 U668 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U669 ( .A1(n606), .A2(n605), .ZN(n608) );
  INV_X1 U670 ( .A(KEYINPUT53), .ZN(n607) );
  INV_X1 U671 ( .A(n609), .ZN(n706) );
  NAND2_X1 U672 ( .A1(n688), .A2(n610), .ZN(n614) );
  XOR2_X1 U673 ( .A(n611), .B(KEYINPUT80), .Z(n612) );
  NAND2_X1 U674 ( .A1(n612), .A2(KEYINPUT2), .ZN(n613) );
  NAND2_X1 U675 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U676 ( .A1(n676), .A2(G475), .ZN(n620) );
  XOR2_X1 U677 ( .A(KEYINPUT59), .B(KEYINPUT64), .Z(n617) );
  INV_X1 U678 ( .A(G952), .ZN(n621) );
  AND2_X1 U679 ( .A1(n621), .A2(G953), .ZN(n687) );
  XNOR2_X1 U680 ( .A(KEYINPUT60), .B(KEYINPUT118), .ZN(n623) );
  XNOR2_X1 U681 ( .A(n624), .B(n623), .ZN(G60) );
  INV_X1 U682 ( .A(n687), .ZN(n681) );
  NAND2_X1 U683 ( .A1(n676), .A2(G210), .ZN(n629) );
  XOR2_X1 U684 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n627) );
  XNOR2_X1 U685 ( .A(n625), .B(KEYINPUT84), .ZN(n626) );
  XNOR2_X1 U686 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U687 ( .A(n629), .B(n628), .ZN(n630) );
  AND2_X1 U688 ( .A1(n681), .A2(n630), .ZN(n632) );
  XNOR2_X1 U689 ( .A(KEYINPUT56), .B(KEYINPUT116), .ZN(n631) );
  XNOR2_X1 U690 ( .A(n632), .B(n631), .ZN(G51) );
  XNOR2_X1 U691 ( .A(n633), .B(G143), .ZN(G45) );
  XOR2_X1 U692 ( .A(G131), .B(KEYINPUT126), .Z(n634) );
  XNOR2_X1 U693 ( .A(n635), .B(n634), .ZN(G33) );
  NAND2_X1 U694 ( .A1(n676), .A2(G472), .ZN(n639) );
  XNOR2_X1 U695 ( .A(KEYINPUT106), .B(KEYINPUT62), .ZN(n636) );
  XNOR2_X1 U696 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U697 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X2 U698 ( .A1(n640), .A2(n687), .ZN(n642) );
  XNOR2_X1 U699 ( .A(KEYINPUT107), .B(KEYINPUT63), .ZN(n641) );
  XNOR2_X1 U700 ( .A(n642), .B(n641), .ZN(G57) );
  XOR2_X1 U701 ( .A(G101), .B(n643), .Z(G3) );
  NAND2_X1 U702 ( .A1(n645), .A2(n660), .ZN(n644) );
  XNOR2_X1 U703 ( .A(n644), .B(G104), .ZN(G6) );
  XOR2_X1 U704 ( .A(KEYINPUT109), .B(KEYINPUT27), .Z(n647) );
  INV_X1 U705 ( .A(n653), .ZN(n663) );
  NAND2_X1 U706 ( .A1(n645), .A2(n663), .ZN(n646) );
  XNOR2_X1 U707 ( .A(n647), .B(n646), .ZN(n648) );
  XOR2_X1 U708 ( .A(n648), .B(KEYINPUT26), .Z(n650) );
  XNOR2_X1 U709 ( .A(G107), .B(KEYINPUT108), .ZN(n649) );
  XNOR2_X1 U710 ( .A(n650), .B(n649), .ZN(G9) );
  XOR2_X1 U711 ( .A(G110), .B(n651), .Z(n652) );
  XNOR2_X1 U712 ( .A(KEYINPUT110), .B(n652), .ZN(G12) );
  NOR2_X1 U713 ( .A1(n653), .A2(n656), .ZN(n655) );
  XNOR2_X1 U714 ( .A(G128), .B(KEYINPUT29), .ZN(n654) );
  XNOR2_X1 U715 ( .A(n655), .B(n654), .ZN(G30) );
  NOR2_X1 U716 ( .A1(n657), .A2(n656), .ZN(n659) );
  XNOR2_X1 U717 ( .A(G146), .B(KEYINPUT111), .ZN(n658) );
  XNOR2_X1 U718 ( .A(n659), .B(n658), .ZN(G48) );
  NAND2_X1 U719 ( .A1(n664), .A2(n660), .ZN(n661) );
  XNOR2_X1 U720 ( .A(n661), .B(KEYINPUT112), .ZN(n662) );
  XNOR2_X1 U721 ( .A(G113), .B(n662), .ZN(G15) );
  XOR2_X1 U722 ( .A(G116), .B(KEYINPUT113), .Z(n666) );
  NAND2_X1 U723 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U724 ( .A(n666), .B(n665), .ZN(G18) );
  XNOR2_X1 U725 ( .A(n667), .B(G134), .ZN(n668) );
  XNOR2_X1 U726 ( .A(KEYINPUT114), .B(n668), .ZN(G36) );
  XNOR2_X1 U727 ( .A(G140), .B(n669), .ZN(G42) );
  NAND2_X1 U728 ( .A1(n683), .A2(G469), .ZN(n674) );
  XOR2_X1 U729 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n670) );
  XNOR2_X1 U730 ( .A(n670), .B(KEYINPUT117), .ZN(n671) );
  XNOR2_X1 U731 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U732 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U733 ( .A1(n687), .A2(n675), .ZN(G54) );
  NAND2_X1 U734 ( .A1(n676), .A2(G478), .ZN(n679) );
  XNOR2_X1 U735 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U736 ( .A1(n683), .A2(G217), .ZN(n684) );
  XNOR2_X1 U737 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U738 ( .A1(n687), .A2(n686), .ZN(G66) );
  NAND2_X1 U739 ( .A1(n707), .A2(n688), .ZN(n692) );
  NAND2_X1 U740 ( .A1(G953), .A2(G224), .ZN(n689) );
  XNOR2_X1 U741 ( .A(KEYINPUT61), .B(n689), .ZN(n690) );
  NAND2_X1 U742 ( .A1(n690), .A2(G898), .ZN(n691) );
  NAND2_X1 U743 ( .A1(n692), .A2(n691), .ZN(n699) );
  XNOR2_X1 U744 ( .A(G101), .B(n693), .ZN(n695) );
  XNOR2_X1 U745 ( .A(n694), .B(n695), .ZN(n697) );
  NOR2_X1 U746 ( .A1(G898), .A2(n707), .ZN(n696) );
  NOR2_X1 U747 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U748 ( .A(n699), .B(n698), .ZN(n700) );
  XOR2_X1 U749 ( .A(KEYINPUT121), .B(n700), .Z(G69) );
  XNOR2_X1 U750 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U751 ( .A(n703), .B(KEYINPUT4), .ZN(n704) );
  XNOR2_X1 U752 ( .A(n705), .B(n704), .ZN(n710) );
  XNOR2_X1 U753 ( .A(n706), .B(n710), .ZN(n708) );
  NAND2_X1 U754 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U755 ( .A(KEYINPUT122), .B(n709), .ZN(n716) );
  XNOR2_X1 U756 ( .A(G227), .B(n710), .ZN(n711) );
  NAND2_X1 U757 ( .A1(n711), .A2(G900), .ZN(n712) );
  XOR2_X1 U758 ( .A(KEYINPUT123), .B(n712), .Z(n713) );
  NAND2_X1 U759 ( .A1(G953), .A2(n713), .ZN(n714) );
  XNOR2_X1 U760 ( .A(KEYINPUT124), .B(n714), .ZN(n715) );
  NAND2_X1 U761 ( .A1(n716), .A2(n715), .ZN(G72) );
  XOR2_X1 U762 ( .A(n717), .B(G137), .Z(G39) );
  XNOR2_X1 U763 ( .A(G125), .B(n718), .ZN(n719) );
  XNOR2_X1 U764 ( .A(n719), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U765 ( .A(n720), .B(G119), .Z(n721) );
  XNOR2_X1 U766 ( .A(KEYINPUT125), .B(n721), .ZN(G21) );
endmodule

