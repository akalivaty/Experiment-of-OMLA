//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT69), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n192), .A2(KEYINPUT16), .A3(G140), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n193), .B1(new_n187), .B2(KEYINPUT16), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  OR2_X1    g012(.A1(new_n198), .A2(KEYINPUT23), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(KEYINPUT23), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n199), .A2(new_n200), .B1(new_n201), .B2(G128), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT68), .B(G110), .Z(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(new_n198), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT24), .B(G110), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n202), .A2(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OR2_X1    g021(.A1(new_n196), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n194), .B(new_n188), .ZN(new_n209));
  INV_X1    g023(.A(G110), .ZN(new_n210));
  OAI22_X1  g024(.A1(new_n202), .A2(new_n210), .B1(new_n205), .B2(new_n206), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G953), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(G221), .A3(G234), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(KEYINPUT22), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n216), .B(G137), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n208), .A2(new_n217), .A3(new_n212), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G217), .ZN(new_n222));
  INV_X1    g036(.A(G902), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(G234), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G902), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n226), .A2(KEYINPUT70), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n219), .A2(new_n223), .A3(new_n220), .ZN(new_n228));
  OR2_X1    g042(.A1(new_n228), .A2(KEYINPUT25), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(KEYINPUT25), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(new_n224), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(KEYINPUT70), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(G472), .A2(G902), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G143), .B(G146), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(G128), .ZN(new_n238));
  OR2_X1    g052(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n239));
  INV_X1    g053(.A(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n239), .A2(new_n240), .A3(G146), .A4(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n188), .A2(G143), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n197), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n238), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT11), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G137), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT11), .A3(G134), .ZN(new_n252));
  INV_X1    g066(.A(G131), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(G137), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n250), .A2(new_n252), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n251), .A2(G134), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n249), .A2(G137), .ZN(new_n257));
  OAI21_X1  g071(.A(G131), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n255), .A2(new_n258), .A3(KEYINPUT64), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT64), .B1(new_n255), .B2(new_n258), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n247), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n250), .A2(new_n254), .A3(new_n252), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G131), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT0), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(new_n197), .ZN(new_n266));
  NOR2_X1   g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n245), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n236), .B1(new_n265), .B2(new_n197), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n264), .A2(new_n255), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT66), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n272), .B(new_n247), .C1(new_n259), .C2(new_n260), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n262), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(G116), .B(G119), .Z(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT2), .B(G113), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n255), .A2(new_n258), .ZN(new_n280));
  AOI21_X1  g094(.A(G128), .B1(new_n243), .B2(new_n244), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n197), .B1(new_n239), .B2(new_n241), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n236), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n280), .B1(new_n283), .B2(new_n242), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n284), .A2(new_n270), .A3(new_n275), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n276), .A2(new_n279), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n284), .A2(new_n270), .ZN(new_n288));
  INV_X1    g102(.A(new_n279), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(G101), .ZN(new_n292));
  NOR2_X1   g106(.A1(G237), .A2(G953), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G210), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n292), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n287), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(KEYINPUT31), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT67), .ZN(new_n300));
  AOI211_X1 g114(.A(new_n289), .B(new_n285), .C1(new_n274), .C2(new_n275), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(new_n296), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n287), .A2(KEYINPUT67), .A3(new_n297), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n299), .B1(new_n304), .B2(KEYINPUT31), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n290), .B(KEYINPUT28), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n274), .A2(new_n279), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n295), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n235), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT32), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n285), .B1(new_n274), .B2(new_n275), .ZN(new_n314));
  AOI211_X1 g128(.A(new_n300), .B(new_n296), .C1(new_n314), .C2(new_n279), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT67), .B1(new_n287), .B2(new_n297), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT31), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n299), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n310), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n234), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT32), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n287), .A2(new_n290), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n309), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n306), .A2(new_n307), .A3(new_n295), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n279), .B1(new_n284), .B2(new_n270), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n306), .A2(new_n329), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n330), .A2(new_n326), .A3(new_n309), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G902), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G472), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n233), .B1(new_n322), .B2(new_n334), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT9), .B(G234), .Z(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n337), .A2(new_n222), .A3(G953), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT86), .ZN(new_n340));
  INV_X1    g154(.A(G116), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(G122), .ZN(new_n342));
  INV_X1    g156(.A(G122), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT86), .A3(G116), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G107), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n341), .A2(G122), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G128), .B(G143), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(G134), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(KEYINPUT14), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n343), .A2(KEYINPUT86), .A3(G116), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT86), .B1(new_n343), .B2(G116), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT87), .ZN(new_n356));
  OR2_X1    g170(.A1(new_n347), .A2(KEYINPUT14), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT87), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n345), .A2(new_n358), .A3(new_n352), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AOI211_X1 g174(.A(new_n349), .B(new_n351), .C1(new_n360), .C2(G107), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n345), .A2(new_n347), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G107), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n363), .A2(new_n348), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n350), .A2(new_n249), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n350), .A2(KEYINPUT13), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n240), .A2(G128), .ZN(new_n367));
  OAI21_X1  g181(.A(G134), .B1(new_n367), .B2(KEYINPUT13), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n365), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n339), .B1(new_n361), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n360), .A2(G107), .ZN(new_n372));
  INV_X1    g186(.A(new_n351), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n348), .A3(new_n373), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n364), .A2(new_n369), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(new_n338), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT88), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(KEYINPUT88), .B(new_n339), .C1(new_n361), .C2(new_n370), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n223), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G478), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n381), .A2(KEYINPUT90), .A3(KEYINPUT15), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(KEYINPUT15), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT90), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n380), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT91), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR4_X1   g202(.A1(new_n380), .A2(KEYINPUT91), .A3(new_n382), .A4(new_n385), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT89), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n380), .A2(new_n390), .A3(new_n383), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n390), .B1(new_n380), .B2(new_n383), .ZN(new_n392));
  OAI22_X1  g206(.A1(new_n388), .A2(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G237), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n214), .A3(G214), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n240), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n293), .A2(G143), .A3(G214), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT17), .A3(G131), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(new_n253), .A3(new_n397), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT83), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(G131), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n396), .A2(new_n403), .A3(new_n253), .A4(new_n397), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n209), .B(new_n399), .C1(new_n405), .C2(KEYINPUT17), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n187), .A2(new_n188), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n191), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT18), .A2(G131), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n398), .B(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G113), .B(G122), .ZN(new_n413));
  INV_X1    g227(.A(G104), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT84), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT84), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n406), .A2(new_n411), .A3(new_n418), .A4(new_n415), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n187), .B(KEYINPUT19), .Z(new_n421));
  OAI211_X1 g235(.A(new_n405), .B(new_n195), .C1(G146), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n411), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n416), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n426));
  NOR2_X1   g240(.A1(G475), .A2(G902), .ZN(new_n427));
  XOR2_X1   g241(.A(new_n427), .B(KEYINPUT85), .Z(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n425), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n431));
  AOI22_X1  g245(.A1(new_n417), .A2(new_n419), .B1(new_n416), .B2(new_n423), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n431), .B1(new_n432), .B2(new_n428), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  OR2_X1    g248(.A1(KEYINPUT92), .A2(G952), .ZN(new_n435));
  NAND2_X1  g249(.A1(KEYINPUT92), .A2(G952), .ZN(new_n436));
  AOI21_X1  g250(.A(G953), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(G234), .A2(G237), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(KEYINPUT21), .B(G898), .Z(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(G902), .A3(G953), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G475), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n412), .A2(new_n416), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n420), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n449), .B2(new_n223), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n434), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n393), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G469), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n264), .A2(new_n255), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT3), .B1(new_n414), .B2(G107), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT3), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n346), .A3(G104), .ZN(new_n458));
  INV_X1    g272(.A(G101), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n414), .A2(G107), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n456), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n346), .A2(G104), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n414), .A2(G107), .ZN(new_n463));
  OAI21_X1  g277(.A(G101), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n247), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n464), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n240), .A2(KEYINPUT1), .A3(G146), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(new_n283), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n455), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT12), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n268), .A2(new_n269), .ZN(new_n472));
  NAND2_X1  g286(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G101), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n473), .B1(new_n475), .B2(new_n461), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n474), .A2(G101), .B1(KEYINPUT71), .B2(KEYINPUT4), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n238), .A2(new_n246), .A3(new_n468), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n465), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT10), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n455), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n247), .A2(new_n465), .A3(KEYINPUT10), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n478), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G110), .B(G140), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n214), .A2(G227), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n486), .B(new_n487), .Z(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n471), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n478), .A2(new_n482), .A3(new_n484), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n455), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n488), .B1(new_n492), .B2(new_n485), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n454), .B(new_n223), .C1(new_n490), .C2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n488), .ZN(new_n495));
  INV_X1    g309(.A(new_n485), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n495), .B1(new_n471), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT72), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n489), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n485), .A2(KEYINPUT72), .A3(new_n488), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n492), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n501), .A3(G469), .ZN(new_n502));
  NAND2_X1  g316(.A1(G469), .A2(G902), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n494), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(G221), .B1(new_n337), .B2(G902), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G214), .B1(G237), .B2(G902), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n507), .B(KEYINPUT73), .Z(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  XOR2_X1   g323(.A(G110), .B(G122), .Z(new_n510));
  OAI21_X1  g324(.A(new_n279), .B1(new_n476), .B2(new_n477), .ZN(new_n511));
  OR2_X1    g325(.A1(new_n277), .A2(new_n278), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n201), .A3(G116), .ZN(new_n514));
  OAI211_X1 g328(.A(G113), .B(new_n514), .C1(new_n277), .C2(new_n513), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n465), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n511), .A2(KEYINPUT74), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT74), .B1(new_n511), .B2(new_n516), .ZN(new_n518));
  OAI211_X1 g332(.A(KEYINPUT75), .B(new_n510), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n510), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n511), .A2(new_n516), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT74), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n511), .A2(KEYINPUT74), .A3(new_n516), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n511), .A2(new_n520), .A3(new_n516), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n526), .A2(KEYINPUT75), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n519), .B(KEYINPUT6), .C1(new_n525), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n247), .A2(new_n192), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n472), .A2(G125), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT77), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT78), .B(G224), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G953), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n532), .B(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n510), .B1(new_n517), .B2(new_n518), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT76), .B1(new_n536), .B2(KEYINPUT6), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT76), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT6), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n525), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n528), .A2(new_n535), .A3(new_n537), .A4(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n529), .A2(new_n530), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n534), .A2(KEYINPUT80), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n534), .A2(KEYINPUT80), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT81), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT7), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n542), .B1(new_n548), .B2(new_n534), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n465), .A2(KEYINPUT79), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n515), .A2(new_n512), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n510), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n547), .A2(new_n526), .A3(new_n549), .A4(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n541), .A2(new_n223), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G210), .B1(G237), .B2(G902), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n541), .A2(new_n223), .A3(new_n555), .A4(new_n557), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n509), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n453), .A2(new_n506), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n335), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT93), .B(G101), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(G3));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n559), .A2(new_n560), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n566), .B1(new_n567), .B2(new_n507), .ZN(new_n568));
  INV_X1    g382(.A(new_n507), .ZN(new_n569));
  AOI211_X1 g383(.A(KEYINPUT94), .B(new_n569), .C1(new_n559), .C2(new_n560), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT33), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n378), .A2(new_n572), .A3(new_n379), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n371), .A2(new_n376), .A3(KEYINPUT33), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n223), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G478), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n380), .A2(G478), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n450), .B1(new_n433), .B2(new_n430), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(new_n445), .ZN(new_n585));
  INV_X1    g399(.A(G472), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n319), .B2(new_n223), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n587), .A2(new_n311), .A3(new_n233), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n571), .A2(new_n585), .A3(new_n506), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT34), .B(G104), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT96), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n589), .B(new_n591), .ZN(G6));
  INV_X1    g406(.A(new_n431), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n425), .B2(new_n429), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n432), .A2(new_n431), .A3(new_n428), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT97), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n425), .A2(new_n593), .A3(new_n429), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n433), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n450), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n393), .A3(new_n446), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n600), .A2(new_n393), .A3(KEYINPUT98), .A4(new_n446), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n605), .A2(new_n506), .A3(new_n588), .A4(new_n571), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n606), .B(KEYINPUT35), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G107), .ZN(G9));
  NAND3_X1  g422(.A1(new_n453), .A2(new_n506), .A3(new_n561), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n319), .A2(new_n223), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n218), .A2(KEYINPUT36), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n213), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n225), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n231), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n611), .A2(new_n320), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT99), .B(KEYINPUT37), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G110), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n617), .B(new_n619), .ZN(G12));
  AND3_X1   g434(.A1(new_n319), .A2(new_n312), .A3(new_n234), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n312), .B1(new_n319), .B2(new_n234), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n334), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n567), .A2(new_n507), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT94), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n567), .A2(new_n566), .A3(new_n507), .ZN(new_n626));
  AND4_X1   g440(.A1(new_n623), .A2(new_n625), .A3(new_n506), .A4(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(G900), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n440), .B1(new_n628), .B2(new_n444), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n600), .A2(new_n393), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n627), .A2(new_n615), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G128), .ZN(G30));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n567), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT38), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n569), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n290), .A2(new_n329), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n304), .B1(new_n295), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n586), .B1(new_n639), .B2(new_n223), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n313), .B2(new_n321), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n629), .B(KEYINPUT39), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n506), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(KEYINPUT40), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n641), .A2(new_n615), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n393), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n582), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n644), .A2(KEYINPUT40), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n637), .A2(new_n646), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G143), .ZN(G45));
  NOR4_X1   g465(.A1(new_n579), .A2(new_n580), .A3(new_n582), .A4(new_n629), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n627), .A2(new_n615), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT101), .B(G146), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G48));
  OR2_X1    g469(.A1(new_n490), .A2(new_n493), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n454), .B1(new_n656), .B2(new_n223), .ZN(new_n657));
  INV_X1    g471(.A(new_n494), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n505), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n568), .A2(new_n570), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n335), .A3(new_n585), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT41), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G113), .ZN(G15));
  NAND3_X1  g478(.A1(new_n661), .A2(new_n605), .A3(new_n335), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G116), .ZN(G18));
  NAND4_X1  g480(.A1(new_n661), .A2(new_n623), .A3(new_n453), .A4(new_n615), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G119), .ZN(G21));
  NOR2_X1   g482(.A1(new_n660), .A2(new_n445), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n625), .A2(new_n626), .A3(new_n648), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n233), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n330), .A2(new_n309), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n235), .B1(new_n305), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(KEYINPUT102), .B1(new_n610), .B2(G472), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n677), .B(new_n586), .C1(new_n319), .C2(new_n223), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n672), .B(new_n675), .C1(new_n676), .C2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(G902), .B1(new_n305), .B2(new_n310), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n677), .B1(new_n682), .B2(new_n586), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n610), .A2(KEYINPUT102), .A3(G472), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n674), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT103), .B1(new_n685), .B2(new_n672), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n669), .B(new_n671), .C1(new_n681), .C2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT104), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G122), .ZN(G24));
  INV_X1    g503(.A(new_n660), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n571), .A2(new_n652), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n683), .A2(new_n684), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n615), .A4(new_n675), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n693), .B1(new_n685), .B2(new_n615), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n691), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT106), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  XNOR2_X1  g513(.A(new_n503), .B(KEYINPUT107), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n502), .A2(KEYINPUT108), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n502), .A2(KEYINPUT108), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n494), .B(new_n700), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n505), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n559), .A2(new_n560), .A3(new_n507), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n623), .A2(new_n706), .A3(new_n652), .A4(new_n672), .ZN(new_n707));
  NAND2_X1  g521(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n707), .A2(new_n710), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n707), .A2(new_n710), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n710), .B1(new_n707), .B2(new_n708), .ZN(new_n717));
  OAI21_X1  g531(.A(KEYINPUT110), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT111), .B(G131), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G33));
  NAND4_X1  g535(.A1(new_n623), .A2(new_n706), .A3(new_n631), .A4(new_n672), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G134), .ZN(G36));
  OR2_X1    g537(.A1(new_n579), .A2(new_n580), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT113), .ZN(new_n725));
  OR3_X1    g539(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT113), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n582), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n582), .B(KEYINPUT114), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(KEYINPUT43), .A3(new_n581), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n587), .A2(new_n311), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n735), .A3(new_n615), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n705), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n497), .A2(new_n501), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT45), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(G469), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n742), .A2(KEYINPUT46), .A3(new_n700), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT46), .B1(new_n742), .B2(new_n700), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n658), .ZN(new_n745));
  INV_X1    g559(.A(new_n505), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n745), .A2(new_n746), .A3(new_n642), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n733), .A2(KEYINPUT44), .A3(new_n735), .A4(new_n615), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n738), .A2(new_n739), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n745), .B2(new_n746), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n744), .A2(new_n658), .ZN(new_n753));
  OAI211_X1 g567(.A(KEYINPUT47), .B(new_n505), .C1(new_n753), .C2(new_n743), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n623), .A2(new_n672), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n652), .A3(new_n739), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G140), .ZN(G42));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n724), .B1(new_n759), .B2(new_n659), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n641), .A2(new_n672), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n505), .B(new_n508), .C1(new_n659), .C2(new_n759), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n636), .A2(new_n731), .A3(new_n760), .A4(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n739), .A2(new_n690), .A3(new_n440), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n582), .A3(new_n724), .ZN(new_n767));
  INV_X1    g581(.A(new_n765), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n733), .B(new_n768), .C1(new_n695), .C2(new_n696), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n657), .A2(new_n505), .A3(new_n658), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n739), .B1(new_n755), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n439), .B1(new_n729), .B2(new_n732), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n679), .A2(new_n680), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n692), .A2(KEYINPUT103), .A3(new_n672), .A4(new_n675), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n767), .B(new_n769), .C1(new_n771), .C2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n772), .A2(new_n775), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n636), .A2(new_n569), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n690), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n778), .A2(KEYINPUT50), .A3(new_n690), .A4(new_n779), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n777), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n437), .B1(new_n784), .B2(KEYINPUT51), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n785), .B1(KEYINPUT51), .B2(new_n784), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n787));
  INV_X1    g601(.A(new_n719), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n627), .B(new_n615), .C1(new_n631), .C2(new_n652), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n641), .A2(new_n615), .A3(new_n629), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n671), .A2(new_n790), .A3(new_n505), .A4(new_n703), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n697), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT52), .ZN(new_n793));
  INV_X1    g607(.A(new_n615), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n393), .A2(new_n794), .A3(new_n629), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n623), .A2(new_n506), .A3(new_n795), .A4(new_n739), .ZN(new_n796));
  INV_X1    g610(.A(new_n600), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n722), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n706), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n615), .B(new_n675), .C1(new_n676), .C2(new_n678), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT105), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n799), .B1(new_n801), .B2(new_n694), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n798), .B1(new_n802), .B2(new_n652), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n697), .A2(new_n789), .A3(new_n791), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n788), .A2(new_n793), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n807));
  INV_X1    g621(.A(new_n669), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n808), .B(new_n670), .C1(new_n773), .C2(new_n774), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n661), .B(new_n335), .C1(new_n605), .C2(new_n585), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n667), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n807), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n687), .A2(KEYINPUT115), .A3(new_n667), .A4(new_n810), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n588), .A2(new_n506), .A3(new_n561), .A4(new_n446), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT116), .B1(new_n581), .B2(new_n583), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n579), .A2(new_n580), .A3(new_n582), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n623), .A2(new_n672), .ZN(new_n820));
  OAI22_X1  g634(.A1(new_n815), .A2(new_n819), .B1(new_n820), .B2(new_n609), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n611), .A2(new_n320), .A3(new_n672), .A4(new_n506), .ZN(new_n822));
  INV_X1    g636(.A(new_n561), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n393), .A2(new_n446), .A3(new_n582), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT117), .B1(new_n825), .B2(new_n617), .ZN(new_n826));
  INV_X1    g640(.A(new_n616), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n562), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n824), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n588), .A2(new_n829), .A3(new_n506), .A4(new_n561), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n821), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n814), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n787), .B1(new_n806), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n793), .A2(new_n805), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n652), .B(new_n706), .C1(new_n695), .C2(new_n696), .ZN(new_n837));
  INV_X1    g651(.A(new_n798), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n719), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n815), .ZN(new_n841));
  INV_X1    g655(.A(new_n819), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n841), .A2(new_n842), .B1(new_n335), .B2(new_n562), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n825), .A2(new_n617), .A3(KEYINPUT117), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n831), .B1(new_n828), .B2(new_n830), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n812), .B2(new_n813), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n836), .A2(KEYINPUT53), .A3(new_n840), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n835), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT54), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n766), .A2(new_n583), .A3(new_n581), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n787), .B1(new_n712), .B2(new_n714), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n793), .A2(new_n805), .A3(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n803), .A2(new_n833), .A3(KEYINPUT118), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT118), .B1(new_n803), .B2(new_n833), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n809), .A2(new_n811), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n853), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n835), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n786), .A2(new_n850), .A3(new_n851), .A4(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n778), .A2(new_n661), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n733), .A2(new_n335), .A3(new_n768), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(KEYINPUT48), .Z(new_n864));
  NOR3_X1   g678(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(G952), .A2(G953), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n764), .B1(new_n865), .B2(new_n866), .ZN(G75));
  NOR2_X1   g681(.A1(new_n214), .A2(G952), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n528), .A2(new_n537), .A3(new_n540), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(new_n535), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT55), .Z(new_n871));
  NAND2_X1  g685(.A1(new_n835), .A2(new_n858), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(G210), .A3(G902), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OR2_X1    g689(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n876));
  NAND2_X1  g690(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n873), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT120), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n873), .A2(new_n881), .A3(new_n876), .A4(new_n878), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n868), .B(new_n875), .C1(new_n880), .C2(new_n882), .ZN(G51));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT118), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n839), .B2(new_n846), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n803), .A2(new_n833), .A3(KEYINPUT118), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n793), .A2(new_n805), .A3(new_n852), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n847), .A2(new_n840), .A3(new_n805), .A4(new_n793), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n857), .A2(new_n890), .B1(new_n891), .B2(new_n787), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n892), .A2(new_n223), .A3(new_n742), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n700), .B(KEYINPUT57), .Z(new_n894));
  AND3_X1   g708(.A1(new_n835), .A2(new_n858), .A3(new_n859), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n859), .B1(new_n835), .B2(new_n858), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n893), .B1(new_n897), .B2(new_n656), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n884), .B1(new_n898), .B2(new_n868), .ZN(new_n899));
  INV_X1    g713(.A(new_n868), .ZN(new_n900));
  INV_X1    g714(.A(new_n656), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n872), .A2(KEYINPUT54), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n860), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n901), .B1(new_n903), .B2(new_n894), .ZN(new_n904));
  OAI211_X1 g718(.A(KEYINPUT121), .B(new_n900), .C1(new_n904), .C2(new_n893), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n899), .A2(new_n905), .ZN(G54));
  NAND4_X1  g720(.A1(new_n872), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n907), .A2(new_n432), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n432), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(new_n868), .ZN(G60));
  NAND2_X1  g724(.A1(new_n573), .A2(new_n574), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT122), .Z(new_n912));
  NAND2_X1  g726(.A1(G478), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT59), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n903), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n850), .A2(new_n860), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n916), .A2(new_n914), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n900), .B(new_n915), .C1(new_n917), .C2(new_n912), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(G63));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n920));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT60), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n920), .B1(new_n872), .B2(new_n923), .ZN(new_n924));
  AOI211_X1 g738(.A(KEYINPUT123), .B(new_n922), .C1(new_n835), .C2(new_n858), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n613), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT123), .B1(new_n892), .B2(new_n922), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n872), .A2(new_n920), .A3(new_n923), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n221), .B(KEYINPUT124), .Z(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n926), .A2(new_n930), .A3(new_n900), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n926), .A2(new_n930), .A3(KEYINPUT61), .A4(new_n900), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(G66));
  OAI21_X1  g749(.A(G953), .B1(new_n442), .B2(new_n533), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n847), .B2(G953), .ZN(new_n937));
  INV_X1    g751(.A(G898), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n869), .B1(new_n938), .B2(G953), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n937), .B(new_n939), .Z(G69));
  XNOR2_X1  g754(.A(new_n314), .B(new_n421), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n214), .A2(G900), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n738), .A2(new_n739), .A3(new_n748), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n820), .B2(new_n670), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n747), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n697), .A2(new_n789), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n947), .A2(new_n757), .A3(new_n722), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n788), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n943), .B1(new_n949), .B2(new_n214), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n719), .B1(new_n945), .B2(new_n747), .ZN(new_n953));
  AOI21_X1  g767(.A(G953), .B1(new_n953), .B2(new_n948), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n954), .A2(KEYINPUT125), .A3(new_n943), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n942), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n214), .B1(G227), .B2(G900), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n650), .A2(new_n947), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n842), .B1(new_n582), .B2(new_n393), .ZN(new_n962));
  OR4_X1    g776(.A1(new_n820), .A2(new_n962), .A3(new_n644), .A4(new_n705), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n749), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n961), .A2(new_n757), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n942), .B1(new_n965), .B2(new_n214), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n956), .A2(new_n958), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n950), .A2(new_n951), .ZN(new_n969));
  OAI21_X1  g783(.A(KEYINPUT125), .B1(new_n954), .B2(new_n943), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n941), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n957), .B1(new_n971), .B2(new_n966), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n968), .A2(new_n972), .ZN(G72));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT63), .Z(new_n975));
  XNOR2_X1  g789(.A(new_n325), .B(KEYINPUT127), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n304), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n849), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n961), .A2(new_n757), .A3(new_n847), .A4(new_n964), .ZN(new_n979));
  AOI211_X1 g793(.A(new_n309), .B(new_n323), .C1(new_n979), .C2(new_n975), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n946), .A2(new_n788), .A3(new_n847), .A4(new_n948), .ZN(new_n981));
  AOI211_X1 g795(.A(new_n295), .B(new_n324), .C1(new_n981), .C2(new_n975), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT126), .B1(new_n982), .B2(new_n868), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n975), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n984), .A2(new_n309), .A3(new_n323), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT126), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n985), .A2(new_n986), .A3(new_n900), .ZN(new_n987));
  AOI211_X1 g801(.A(new_n978), .B(new_n980), .C1(new_n983), .C2(new_n987), .ZN(G57));
endmodule


