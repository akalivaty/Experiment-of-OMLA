

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736;

  BUF_X1 U366 ( .A(G101), .Z(n345) );
  NOR2_X1 U367 ( .A1(n565), .A2(n564), .ZN(n402) );
  NAND2_X2 U368 ( .A1(n416), .A2(n415), .ZN(n414) );
  XNOR2_X2 U369 ( .A(n720), .B(n452), .ZN(n692) );
  XNOR2_X2 U370 ( .A(n358), .B(n552), .ZN(n565) );
  NOR2_X2 U371 ( .A1(n734), .A2(n352), .ZN(n578) );
  XNOR2_X2 U372 ( .A(n412), .B(n411), .ZN(n734) );
  INV_X1 U373 ( .A(G953), .ZN(n722) );
  XNOR2_X2 U374 ( .A(n444), .B(n349), .ZN(n551) );
  INV_X2 U375 ( .A(n437), .ZN(n439) );
  XNOR2_X2 U376 ( .A(G128), .B(KEYINPUT76), .ZN(n437) );
  OR2_X2 U377 ( .A1(n692), .A2(G902), .ZN(n376) );
  XNOR2_X2 U378 ( .A(n536), .B(KEYINPUT1), .ZN(n600) );
  NOR2_X1 U379 ( .A1(n598), .A2(n597), .ZN(n396) );
  AND2_X1 U380 ( .A1(n382), .A2(n379), .ZN(n378) );
  AND2_X1 U381 ( .A1(n581), .A2(n387), .ZN(n386) );
  AND2_X1 U382 ( .A1(n580), .A2(n353), .ZN(n387) );
  AND2_X1 U383 ( .A1(n583), .A2(n732), .ZN(n404) );
  AND2_X1 U384 ( .A1(n679), .A2(n560), .ZN(n546) );
  XNOR2_X1 U385 ( .A(n509), .B(n362), .ZN(n577) );
  XNOR2_X1 U386 ( .A(n504), .B(n405), .ZN(n712) );
  XNOR2_X1 U387 ( .A(n407), .B(n406), .ZN(n504) );
  XNOR2_X1 U388 ( .A(n461), .B(n446), .ZN(n418) );
  XNOR2_X1 U389 ( .A(n445), .B(G131), .ZN(n461) );
  INV_X1 U390 ( .A(KEYINPUT79), .ZN(n423) );
  XNOR2_X1 U391 ( .A(G119), .B(KEYINPUT3), .ZN(n406) );
  NAND2_X1 U392 ( .A1(n432), .A2(n431), .ZN(n407) );
  XNOR2_X1 U393 ( .A(G104), .B(G110), .ZN(n427) );
  NOR2_X1 U394 ( .A1(n721), .A2(n421), .ZN(n366) );
  XOR2_X1 U395 ( .A(G902), .B(KEYINPUT15), .Z(n641) );
  XNOR2_X1 U396 ( .A(n501), .B(n368), .ZN(n367) );
  INV_X1 U397 ( .A(KEYINPUT5), .ZN(n368) );
  XOR2_X1 U398 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n502) );
  AND2_X1 U399 ( .A1(n550), .A2(n351), .ZN(n359) );
  NOR2_X1 U400 ( .A1(n398), .A2(n397), .ZN(n381) );
  XNOR2_X1 U401 ( .A(n433), .B(n372), .ZN(n371) );
  XOR2_X1 U402 ( .A(G146), .B(G125), .Z(n433) );
  XNOR2_X1 U403 ( .A(KEYINPUT18), .B(KEYINPUT89), .ZN(n434) );
  XOR2_X1 U404 ( .A(KEYINPUT17), .B(KEYINPUT75), .Z(n435) );
  INV_X1 U405 ( .A(KEYINPUT4), .ZN(n440) );
  INV_X1 U406 ( .A(G472), .ZN(n362) );
  XNOR2_X1 U407 ( .A(KEYINPUT16), .B(G122), .ZN(n405) );
  XNOR2_X1 U408 ( .A(n364), .B(n463), .ZN(n662) );
  XNOR2_X1 U409 ( .A(n462), .B(n350), .ZN(n364) );
  XNOR2_X1 U410 ( .A(n428), .B(n711), .ZN(n451) );
  AND2_X1 U411 ( .A1(n513), .A2(n611), .ZN(n517) );
  BUF_X1 U412 ( .A(n551), .Z(n530) );
  XNOR2_X1 U413 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n574) );
  NOR2_X1 U414 ( .A1(G953), .A2(G237), .ZN(n500) );
  XNOR2_X1 U415 ( .A(G146), .B(KEYINPUT68), .ZN(n445) );
  NAND2_X1 U416 ( .A1(G234), .A2(G237), .ZN(n476) );
  INV_X1 U417 ( .A(KEYINPUT33), .ZN(n413) );
  OR2_X1 U418 ( .A1(G237), .A2(G902), .ZN(n512) );
  INV_X1 U419 ( .A(n688), .ZN(n380) );
  XNOR2_X1 U420 ( .A(n401), .B(KEYINPUT10), .ZN(n719) );
  XNOR2_X1 U421 ( .A(G140), .B(G125), .ZN(n401) );
  XOR2_X1 U422 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n456) );
  XNOR2_X1 U423 ( .A(KEYINPUT101), .B(KEYINPUT99), .ZN(n455) );
  XNOR2_X1 U424 ( .A(G143), .B(G113), .ZN(n457) );
  XOR2_X1 U425 ( .A(G122), .B(G104), .Z(n458) );
  NAND2_X1 U426 ( .A1(n424), .A2(n422), .ZN(n419) );
  NOR2_X1 U427 ( .A1(n640), .A2(n423), .ZN(n422) );
  XNOR2_X1 U428 ( .A(n367), .B(n502), .ZN(n506) );
  XOR2_X1 U429 ( .A(KEYINPUT95), .B(KEYINPUT24), .Z(n492) );
  XNOR2_X1 U430 ( .A(G137), .B(G110), .ZN(n491) );
  XNOR2_X1 U431 ( .A(n719), .B(n400), .ZN(n489) );
  INV_X1 U432 ( .A(KEYINPUT94), .ZN(n400) );
  XNOR2_X1 U433 ( .A(G128), .B(G146), .ZN(n486) );
  XOR2_X1 U434 ( .A(G122), .B(G107), .Z(n468) );
  XNOR2_X1 U435 ( .A(G134), .B(G116), .ZN(n467) );
  INV_X1 U436 ( .A(KEYINPUT92), .ZN(n417) );
  XOR2_X1 U437 ( .A(KEYINPUT93), .B(G140), .Z(n449) );
  XNOR2_X1 U438 ( .A(n447), .B(n370), .ZN(n441) );
  XNOR2_X1 U439 ( .A(n436), .B(n371), .ZN(n370) );
  NOR2_X1 U440 ( .A1(n542), .A2(n541), .ZN(n545) );
  XNOR2_X1 U441 ( .A(n663), .B(KEYINPUT59), .ZN(n664) );
  NOR2_X1 U442 ( .A1(n369), .A2(n514), .ZN(n515) );
  XNOR2_X1 U443 ( .A(n518), .B(n363), .ZN(n519) );
  XNOR2_X1 U444 ( .A(KEYINPUT84), .B(KEYINPUT36), .ZN(n363) );
  INV_X1 U445 ( .A(KEYINPUT32), .ZN(n411) );
  AND2_X1 U446 ( .A1(n598), .A2(n347), .ZN(n410) );
  NOR2_X1 U447 ( .A1(n554), .A2(n555), .ZN(n679) );
  XNOR2_X1 U448 ( .A(n374), .B(KEYINPUT81), .ZN(n373) );
  AND2_X1 U449 ( .A1(n388), .A2(n585), .ZN(n375) );
  OR2_X1 U450 ( .A1(n415), .A2(n409), .ZN(n346) );
  AND2_X1 U451 ( .A1(n388), .A2(n603), .ZN(n347) );
  AND2_X1 U452 ( .A1(n373), .A2(n409), .ZN(n348) );
  XOR2_X1 U453 ( .A(n443), .B(KEYINPUT77), .Z(n349) );
  XOR2_X1 U454 ( .A(n454), .B(n453), .Z(n350) );
  XOR2_X1 U455 ( .A(KEYINPUT47), .B(n558), .Z(n351) );
  AND2_X1 U456 ( .A1(n584), .A2(n410), .ZN(n352) );
  NOR2_X1 U457 ( .A1(n348), .A2(n593), .ZN(n353) );
  AND2_X1 U458 ( .A1(n420), .A2(n366), .ZN(n354) );
  XOR2_X1 U459 ( .A(G469), .B(KEYINPUT69), .Z(n355) );
  INV_X1 U460 ( .A(n598), .ZN(n409) );
  OR2_X1 U461 ( .A1(n567), .A2(KEYINPUT34), .ZN(n356) );
  BUF_X2 U462 ( .A(n600), .Z(n369) );
  XNOR2_X1 U463 ( .A(KEYINPUT66), .B(n642), .ZN(n357) );
  INV_X1 U464 ( .A(KEYINPUT80), .ZN(n397) );
  XOR2_X1 U465 ( .A(KEYINPUT88), .B(n652), .Z(n690) );
  NOR2_X1 U466 ( .A1(n730), .A2(n735), .ZN(n548) );
  AND2_X1 U467 ( .A1(n359), .A2(n549), .ZN(n399) );
  NAND2_X1 U468 ( .A1(n577), .A2(n611), .ZN(n521) );
  NOR2_X1 U469 ( .A1(n576), .A2(n346), .ZN(n408) );
  NAND2_X1 U470 ( .A1(n551), .A2(n611), .ZN(n358) );
  XOR2_X2 U471 ( .A(G101), .B(KEYINPUT67), .Z(n503) );
  AND2_X1 U472 ( .A1(n360), .A2(n690), .ZN(G63) );
  XNOR2_X1 U473 ( .A(n697), .B(n361), .ZN(n360) );
  INV_X1 U474 ( .A(n698), .ZN(n361) );
  XNOR2_X2 U475 ( .A(n496), .B(n365), .ZN(n598) );
  NOR2_X1 U476 ( .A1(n699), .A2(G902), .ZN(n365) );
  NAND2_X1 U477 ( .A1(n384), .A2(n383), .ZN(n382) );
  XNOR2_X1 U478 ( .A(n399), .B(KEYINPUT48), .ZN(n384) );
  NAND2_X1 U479 ( .A1(n354), .A2(n419), .ZN(n643) );
  INV_X1 U480 ( .A(n689), .ZN(n398) );
  NAND2_X1 U481 ( .A1(n722), .A2(G224), .ZN(n372) );
  XNOR2_X2 U482 ( .A(n466), .B(n440), .ZN(n447) );
  XNOR2_X2 U483 ( .A(n439), .B(n438), .ZN(n466) );
  NAND2_X1 U484 ( .A1(n584), .A2(n375), .ZN(n374) );
  XNOR2_X1 U485 ( .A(n369), .B(KEYINPUT87), .ZN(n576) );
  NOR2_X1 U486 ( .A1(n579), .A2(KEYINPUT44), .ZN(n583) );
  XNOR2_X1 U487 ( .A(n578), .B(KEYINPUT83), .ZN(n579) );
  NAND2_X1 U488 ( .A1(n396), .A2(n536), .ZN(n591) );
  XNOR2_X2 U489 ( .A(n376), .B(n355), .ZN(n536) );
  NAND2_X2 U490 ( .A1(n378), .A2(n377), .ZN(n721) );
  OR2_X1 U491 ( .A1(n384), .A2(n397), .ZN(n377) );
  NOR2_X1 U492 ( .A1(n381), .A2(n380), .ZN(n379) );
  NOR2_X1 U493 ( .A1(n689), .A2(KEYINPUT80), .ZN(n383) );
  XNOR2_X2 U494 ( .A(n385), .B(n594), .ZN(n708) );
  NAND2_X1 U495 ( .A1(n403), .A2(n386), .ZN(n385) );
  INV_X1 U496 ( .A(n369), .ZN(n388) );
  NAND2_X1 U497 ( .A1(n389), .A2(n394), .ZN(n570) );
  NAND2_X1 U498 ( .A1(n392), .A2(n390), .ZN(n389) );
  NAND2_X1 U499 ( .A1(n610), .A2(n391), .ZN(n390) );
  INV_X1 U500 ( .A(KEYINPUT34), .ZN(n391) );
  NAND2_X1 U501 ( .A1(n393), .A2(n356), .ZN(n392) );
  INV_X1 U502 ( .A(n610), .ZN(n393) );
  XNOR2_X2 U503 ( .A(n414), .B(n413), .ZN(n610) );
  AND2_X1 U504 ( .A1(n395), .A2(n569), .ZN(n394) );
  NAND2_X1 U505 ( .A1(n567), .A2(KEYINPUT34), .ZN(n395) );
  NAND2_X1 U506 ( .A1(n600), .A2(n396), .ZN(n587) );
  NOR2_X1 U507 ( .A1(n369), .A2(n396), .ZN(n601) );
  XNOR2_X2 U508 ( .A(G143), .B(KEYINPUT65), .ZN(n438) );
  OR2_X2 U509 ( .A1(n644), .A2(n645), .ZN(n425) );
  OR2_X2 U510 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U511 ( .A(n402), .B(n566), .ZN(n573) );
  XNOR2_X1 U512 ( .A(n404), .B(KEYINPUT71), .ZN(n403) );
  NAND2_X1 U513 ( .A1(n584), .A2(n408), .ZN(n412) );
  INV_X1 U514 ( .A(n585), .ZN(n415) );
  XNOR2_X1 U515 ( .A(n587), .B(KEYINPUT105), .ZN(n416) );
  XNOR2_X2 U516 ( .A(n508), .B(n417), .ZN(n720) );
  XNOR2_X2 U517 ( .A(n447), .B(n418), .ZN(n508) );
  NAND2_X1 U518 ( .A1(n708), .A2(n423), .ZN(n420) );
  AND2_X1 U519 ( .A1(n640), .A2(n423), .ZN(n421) );
  INV_X1 U520 ( .A(n708), .ZN(n424) );
  BUF_X1 U521 ( .A(n610), .Z(n630) );
  XOR2_X1 U522 ( .A(n492), .B(n491), .Z(n426) );
  XNOR2_X1 U523 ( .A(n503), .B(KEYINPUT70), .ZN(n428) );
  NAND2_X1 U524 ( .A1(n615), .A2(n520), .ZN(n572) );
  XNOR2_X1 U525 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U526 ( .A(n493), .B(n426), .ZN(n494) );
  INV_X1 U527 ( .A(KEYINPUT72), .ZN(n543) );
  XNOR2_X1 U528 ( .A(n495), .B(n494), .ZN(n699) );
  XNOR2_X1 U529 ( .A(n543), .B(KEYINPUT39), .ZN(n544) );
  XNOR2_X1 U530 ( .A(n692), .B(n693), .ZN(n694) );
  XNOR2_X1 U531 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U532 ( .A(n639), .B(n638), .ZN(G75) );
  INV_X1 U533 ( .A(KEYINPUT2), .ZN(n645) );
  XNOR2_X1 U534 ( .A(n427), .B(G107), .ZN(n711) );
  INV_X1 U535 ( .A(G116), .ZN(n429) );
  NAND2_X1 U536 ( .A1(G113), .A2(n429), .ZN(n432) );
  INV_X1 U537 ( .A(G113), .ZN(n430) );
  NAND2_X1 U538 ( .A1(n430), .A2(G116), .ZN(n431) );
  XNOR2_X1 U539 ( .A(n451), .B(n712), .ZN(n442) );
  XNOR2_X1 U540 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U541 ( .A(n442), .B(n441), .ZN(n647) );
  OR2_X2 U542 ( .A1(n647), .A2(n641), .ZN(n444) );
  AND2_X1 U543 ( .A1(G210), .A2(n512), .ZN(n443) );
  XOR2_X1 U544 ( .A(G134), .B(G137), .Z(n446) );
  NAND2_X1 U545 ( .A1(G227), .A2(n722), .ZN(n448) );
  XNOR2_X1 U546 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U547 ( .A(KEYINPUT13), .B(G475), .ZN(n465) );
  XOR2_X1 U548 ( .A(KEYINPUT102), .B(KEYINPUT12), .Z(n454) );
  NAND2_X1 U549 ( .A1(G214), .A2(n500), .ZN(n453) );
  XNOR2_X1 U550 ( .A(n456), .B(n455), .ZN(n460) );
  XNOR2_X1 U551 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U552 ( .A(n460), .B(n459), .Z(n463) );
  XNOR2_X1 U553 ( .A(n719), .B(n461), .ZN(n462) );
  NOR2_X1 U554 ( .A1(G902), .A2(n662), .ZN(n464) );
  XNOR2_X1 U555 ( .A(n465), .B(n464), .ZN(n531) );
  INV_X1 U556 ( .A(n531), .ZN(n554) );
  XNOR2_X1 U557 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U558 ( .A(n466), .B(n469), .ZN(n474) );
  XOR2_X1 U559 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n472) );
  NAND2_X1 U560 ( .A1(G234), .A2(n722), .ZN(n470) );
  XOR2_X1 U561 ( .A(KEYINPUT8), .B(n470), .Z(n490) );
  NAND2_X1 U562 ( .A1(G217), .A2(n490), .ZN(n471) );
  XNOR2_X1 U563 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U564 ( .A(n474), .B(n473), .ZN(n698) );
  NOR2_X1 U565 ( .A1(G902), .A2(n698), .ZN(n475) );
  XOR2_X1 U566 ( .A(G478), .B(n475), .Z(n555) );
  INV_X1 U567 ( .A(n679), .ZN(n556) );
  XNOR2_X1 U568 ( .A(KEYINPUT14), .B(n476), .ZN(n479) );
  NAND2_X1 U569 ( .A1(G902), .A2(n479), .ZN(n561) );
  OR2_X1 U570 ( .A1(n722), .A2(n561), .ZN(n477) );
  XOR2_X1 U571 ( .A(KEYINPUT107), .B(n477), .Z(n478) );
  NOR2_X1 U572 ( .A1(G900), .A2(n478), .ZN(n481) );
  NAND2_X1 U573 ( .A1(n479), .A2(G952), .ZN(n480) );
  XNOR2_X1 U574 ( .A(n480), .B(KEYINPUT90), .ZN(n628) );
  NOR2_X1 U575 ( .A1(G953), .A2(n628), .ZN(n563) );
  NOR2_X1 U576 ( .A1(n481), .A2(n563), .ZN(n523) );
  XOR2_X1 U577 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n484) );
  INV_X1 U578 ( .A(n641), .ZN(n640) );
  NAND2_X1 U579 ( .A1(n640), .A2(G234), .ZN(n482) );
  XNOR2_X1 U580 ( .A(n482), .B(KEYINPUT20), .ZN(n497) );
  NAND2_X1 U581 ( .A1(G217), .A2(n497), .ZN(n483) );
  XNOR2_X1 U582 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U583 ( .A(KEYINPUT74), .B(n485), .ZN(n496) );
  XNOR2_X1 U584 ( .A(n486), .B(KEYINPUT23), .ZN(n487) );
  XNOR2_X1 U585 ( .A(G119), .B(n487), .ZN(n488) );
  XNOR2_X1 U586 ( .A(n489), .B(n488), .ZN(n495) );
  NAND2_X1 U587 ( .A1(G221), .A2(n490), .ZN(n493) );
  NAND2_X1 U588 ( .A1(G221), .A2(n497), .ZN(n498) );
  XOR2_X1 U589 ( .A(KEYINPUT21), .B(n498), .Z(n520) );
  NAND2_X1 U590 ( .A1(n598), .A2(n520), .ZN(n499) );
  NOR2_X1 U591 ( .A1(n523), .A2(n499), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n500), .A2(G210), .ZN(n501) );
  XNOR2_X1 U593 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U594 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U595 ( .A(n508), .B(n507), .ZN(n656) );
  NOR2_X1 U596 ( .A1(G902), .A2(n656), .ZN(n509) );
  XOR2_X1 U597 ( .A(KEYINPUT6), .B(KEYINPUT104), .Z(n510) );
  XOR2_X1 U598 ( .A(n577), .B(n510), .Z(n585) );
  NAND2_X1 U599 ( .A1(n534), .A2(n415), .ZN(n511) );
  NOR2_X1 U600 ( .A1(n556), .A2(n511), .ZN(n513) );
  NAND2_X1 U601 ( .A1(G214), .A2(n512), .ZN(n611) );
  XOR2_X1 U602 ( .A(KEYINPUT108), .B(n517), .Z(n514) );
  XNOR2_X1 U603 ( .A(n515), .B(KEYINPUT43), .ZN(n516) );
  NOR2_X1 U604 ( .A1(n530), .A2(n516), .ZN(n689) );
  NAND2_X1 U605 ( .A1(n517), .A2(n530), .ZN(n518) );
  NOR2_X1 U606 ( .A1(n576), .A2(n519), .ZN(n685) );
  INV_X1 U607 ( .A(n520), .ZN(n597) );
  XNOR2_X1 U608 ( .A(n591), .B(KEYINPUT109), .ZN(n525) );
  XNOR2_X1 U609 ( .A(n521), .B(KEYINPUT30), .ZN(n522) );
  NOR2_X1 U610 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U611 ( .A1(n525), .A2(n524), .ZN(n542) );
  NAND2_X1 U612 ( .A1(n531), .A2(n555), .ZN(n526) );
  XNOR2_X1 U613 ( .A(KEYINPUT106), .B(n526), .ZN(n568) );
  NOR2_X1 U614 ( .A1(n542), .A2(n568), .ZN(n527) );
  NAND2_X1 U615 ( .A1(n530), .A2(n527), .ZN(n528) );
  XNOR2_X1 U616 ( .A(KEYINPUT110), .B(n528), .ZN(n736) );
  XOR2_X1 U617 ( .A(n736), .B(KEYINPUT78), .Z(n529) );
  NOR2_X1 U618 ( .A1(n685), .A2(n529), .ZN(n550) );
  XNOR2_X1 U619 ( .A(KEYINPUT38), .B(n530), .ZN(n541) );
  INV_X1 U620 ( .A(n541), .ZN(n612) );
  NAND2_X1 U621 ( .A1(n612), .A2(n611), .ZN(n618) );
  NOR2_X1 U622 ( .A1(n531), .A2(n555), .ZN(n615) );
  INV_X1 U623 ( .A(n615), .ZN(n532) );
  NOR2_X1 U624 ( .A1(n618), .A2(n532), .ZN(n533) );
  XNOR2_X1 U625 ( .A(n533), .B(KEYINPUT41), .ZN(n629) );
  AND2_X1 U626 ( .A1(n577), .A2(n534), .ZN(n535) );
  XNOR2_X1 U627 ( .A(n535), .B(KEYINPUT28), .ZN(n538) );
  XOR2_X1 U628 ( .A(n536), .B(KEYINPUT111), .Z(n537) );
  NAND2_X1 U629 ( .A1(n538), .A2(n537), .ZN(n553) );
  NOR2_X1 U630 ( .A1(n629), .A2(n553), .ZN(n540) );
  XNOR2_X1 U631 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n539) );
  XNOR2_X1 U632 ( .A(n540), .B(n539), .ZN(n730) );
  XNOR2_X1 U633 ( .A(n545), .B(n544), .ZN(n560) );
  XNOR2_X1 U634 ( .A(n546), .B(KEYINPUT40), .ZN(n735) );
  XNOR2_X1 U635 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n547) );
  XNOR2_X1 U636 ( .A(n548), .B(n547), .ZN(n549) );
  INV_X1 U637 ( .A(KEYINPUT19), .ZN(n552) );
  NOR2_X1 U638 ( .A1(n553), .A2(n565), .ZN(n677) );
  NAND2_X1 U639 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U640 ( .A1(n556), .A2(n559), .ZN(n557) );
  XOR2_X1 U641 ( .A(KEYINPUT103), .B(n557), .Z(n586) );
  NAND2_X1 U642 ( .A1(n677), .A2(n586), .ZN(n558) );
  INV_X1 U643 ( .A(n559), .ZN(n681) );
  NAND2_X1 U644 ( .A1(n681), .A2(n560), .ZN(n688) );
  INV_X1 U645 ( .A(n721), .ZN(n596) );
  XNOR2_X1 U646 ( .A(G898), .B(KEYINPUT91), .ZN(n707) );
  NAND2_X1 U647 ( .A1(G953), .A2(n707), .ZN(n714) );
  NOR2_X1 U648 ( .A1(n561), .A2(n714), .ZN(n562) );
  NOR2_X1 U649 ( .A1(n563), .A2(n562), .ZN(n564) );
  INV_X1 U650 ( .A(KEYINPUT0), .ZN(n566) );
  BUF_X1 U651 ( .A(n573), .Z(n567) );
  INV_X1 U652 ( .A(n568), .ZN(n569) );
  XNOR2_X1 U653 ( .A(n570), .B(KEYINPUT35), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n582), .A2(KEYINPUT44), .ZN(n571) );
  XNOR2_X1 U655 ( .A(n571), .B(KEYINPUT82), .ZN(n581) );
  XNOR2_X2 U656 ( .A(n575), .B(n574), .ZN(n584) );
  INV_X1 U657 ( .A(n577), .ZN(n603) );
  NAND2_X1 U658 ( .A1(n579), .A2(KEYINPUT44), .ZN(n580) );
  INV_X1 U659 ( .A(n582), .ZN(n732) );
  INV_X1 U660 ( .A(n586), .ZN(n617) );
  INV_X1 U661 ( .A(n567), .ZN(n589) );
  NOR2_X1 U662 ( .A1(n603), .A2(n587), .ZN(n607) );
  NAND2_X1 U663 ( .A1(n589), .A2(n607), .ZN(n588) );
  XNOR2_X1 U664 ( .A(n588), .B(KEYINPUT31), .ZN(n682) );
  NAND2_X1 U665 ( .A1(n603), .A2(n589), .ZN(n590) );
  NOR2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n670) );
  NOR2_X1 U667 ( .A1(n682), .A2(n670), .ZN(n592) );
  NOR2_X1 U668 ( .A1(n617), .A2(n592), .ZN(n593) );
  INV_X1 U669 ( .A(KEYINPUT45), .ZN(n594) );
  INV_X1 U670 ( .A(n708), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n644) );
  XNOR2_X1 U672 ( .A(n645), .B(n644), .ZN(n635) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n599), .B(KEYINPUT49), .ZN(n605) );
  XOR2_X1 U675 ( .A(KEYINPUT50), .B(n601), .Z(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U679 ( .A(KEYINPUT51), .B(n608), .Z(n609) );
  NOR2_X1 U680 ( .A1(n629), .A2(n609), .ZN(n625) );
  NOR2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U682 ( .A(KEYINPUT116), .B(n613), .Z(n614) );
  NAND2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U684 ( .A(n616), .B(KEYINPUT117), .ZN(n620) );
  NOR2_X1 U685 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U686 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U687 ( .A(n621), .B(KEYINPUT118), .ZN(n622) );
  NOR2_X1 U688 ( .A1(n630), .A2(n622), .ZN(n623) );
  XOR2_X1 U689 ( .A(KEYINPUT119), .B(n623), .Z(n624) );
  NOR2_X1 U690 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U691 ( .A(n626), .B(KEYINPUT52), .ZN(n627) );
  NOR2_X1 U692 ( .A1(n628), .A2(n627), .ZN(n633) );
  NOR2_X1 U693 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U694 ( .A(KEYINPUT120), .B(n631), .ZN(n632) );
  NOR2_X1 U695 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U696 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U697 ( .A1(G953), .A2(n636), .ZN(n639) );
  INV_X1 U698 ( .A(KEYINPUT53), .ZN(n637) );
  XNOR2_X1 U699 ( .A(n637), .B(KEYINPUT121), .ZN(n638) );
  NAND2_X1 U700 ( .A1(n641), .A2(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U701 ( .A1(n643), .A2(n357), .ZN(n646) );
  AND2_X2 U702 ( .A1(n646), .A2(n425), .ZN(n691) );
  NAND2_X1 U703 ( .A1(G210), .A2(n691), .ZN(n651) );
  XOR2_X1 U704 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n649) );
  XNOR2_X1 U705 ( .A(n647), .B(KEYINPUT85), .ZN(n648) );
  XNOR2_X1 U706 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U707 ( .A(n651), .B(n650), .ZN(n653) );
  NOR2_X1 U708 ( .A1(G952), .A2(n722), .ZN(n652) );
  NAND2_X1 U709 ( .A1(n653), .A2(n690), .ZN(n655) );
  INV_X1 U710 ( .A(KEYINPUT56), .ZN(n654) );
  XNOR2_X1 U711 ( .A(n655), .B(n654), .ZN(G51) );
  NAND2_X1 U712 ( .A1(G472), .A2(n691), .ZN(n659) );
  XOR2_X1 U713 ( .A(n656), .B(KEYINPUT62), .Z(n657) );
  XNOR2_X1 U714 ( .A(n657), .B(KEYINPUT86), .ZN(n658) );
  XNOR2_X1 U715 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U716 ( .A1(n660), .A2(n690), .ZN(n661) );
  XNOR2_X1 U717 ( .A(n661), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U718 ( .A1(n691), .A2(G475), .ZN(n665) );
  XNOR2_X1 U719 ( .A(n662), .B(KEYINPUT122), .ZN(n663) );
  XNOR2_X1 U720 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U721 ( .A1(n666), .A2(n690), .ZN(n668) );
  INV_X1 U722 ( .A(KEYINPUT60), .ZN(n667) );
  XNOR2_X1 U723 ( .A(n668), .B(n667), .ZN(G60) );
  XOR2_X1 U724 ( .A(n345), .B(n348), .Z(G3) );
  NAND2_X1 U725 ( .A1(n670), .A2(n679), .ZN(n669) );
  XNOR2_X1 U726 ( .A(n669), .B(G104), .ZN(G6) );
  XOR2_X1 U727 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n672) );
  NAND2_X1 U728 ( .A1(n670), .A2(n681), .ZN(n671) );
  XNOR2_X1 U729 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U730 ( .A(G107), .B(n673), .ZN(G9) );
  XOR2_X1 U731 ( .A(G110), .B(n352), .Z(G12) );
  XOR2_X1 U732 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n675) );
  NAND2_X1 U733 ( .A1(n677), .A2(n681), .ZN(n674) );
  XNOR2_X1 U734 ( .A(n675), .B(n674), .ZN(n676) );
  XOR2_X1 U735 ( .A(G128), .B(n676), .Z(G30) );
  NAND2_X1 U736 ( .A1(n677), .A2(n679), .ZN(n678) );
  XNOR2_X1 U737 ( .A(n678), .B(G146), .ZN(G48) );
  NAND2_X1 U738 ( .A1(n679), .A2(n682), .ZN(n680) );
  XNOR2_X1 U739 ( .A(G113), .B(n680), .ZN(G15) );
  NAND2_X1 U740 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U741 ( .A(n683), .B(KEYINPUT114), .ZN(n684) );
  XNOR2_X1 U742 ( .A(G116), .B(n684), .ZN(G18) );
  XNOR2_X1 U743 ( .A(G125), .B(n685), .ZN(n686) );
  XNOR2_X1 U744 ( .A(n686), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U745 ( .A(G134), .B(KEYINPUT115), .Z(n687) );
  XNOR2_X1 U746 ( .A(n688), .B(n687), .ZN(G36) );
  XOR2_X1 U747 ( .A(G140), .B(n689), .Z(G42) );
  INV_X1 U748 ( .A(n690), .ZN(n703) );
  BUF_X2 U749 ( .A(n691), .Z(n700) );
  NAND2_X1 U750 ( .A1(n700), .A2(G469), .ZN(n695) );
  XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n693) );
  NOR2_X1 U752 ( .A1(n703), .A2(n696), .ZN(G54) );
  NAND2_X1 U753 ( .A1(G478), .A2(n700), .ZN(n697) );
  XOR2_X1 U754 ( .A(n699), .B(KEYINPUT123), .Z(n702) );
  NAND2_X1 U755 ( .A1(n700), .A2(G217), .ZN(n701) );
  XNOR2_X1 U756 ( .A(n702), .B(n701), .ZN(n704) );
  NOR2_X1 U757 ( .A1(n704), .A2(n703), .ZN(G66) );
  NAND2_X1 U758 ( .A1(G953), .A2(G224), .ZN(n705) );
  XOR2_X1 U759 ( .A(KEYINPUT61), .B(n705), .Z(n706) );
  NOR2_X1 U760 ( .A1(n707), .A2(n706), .ZN(n710) );
  NOR2_X1 U761 ( .A1(G953), .A2(n708), .ZN(n709) );
  NOR2_X1 U762 ( .A1(n710), .A2(n709), .ZN(n717) );
  XNOR2_X1 U763 ( .A(n345), .B(n711), .ZN(n713) );
  XNOR2_X1 U764 ( .A(n713), .B(n712), .ZN(n715) );
  NAND2_X1 U765 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U766 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U767 ( .A(KEYINPUT124), .B(n718), .ZN(G69) );
  XNOR2_X1 U768 ( .A(n719), .B(n720), .ZN(n724) );
  XNOR2_X1 U769 ( .A(n724), .B(n721), .ZN(n723) );
  NAND2_X1 U770 ( .A1(n723), .A2(n722), .ZN(n729) );
  XNOR2_X1 U771 ( .A(G227), .B(n724), .ZN(n725) );
  NAND2_X1 U772 ( .A1(n725), .A2(G900), .ZN(n726) );
  XOR2_X1 U773 ( .A(KEYINPUT125), .B(n726), .Z(n727) );
  NAND2_X1 U774 ( .A1(G953), .A2(n727), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n729), .A2(n728), .ZN(G72) );
  XNOR2_X1 U776 ( .A(G137), .B(n730), .ZN(n731) );
  XNOR2_X1 U777 ( .A(n731), .B(KEYINPUT127), .ZN(G39) );
  XNOR2_X1 U778 ( .A(G122), .B(KEYINPUT126), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n733), .B(n732), .ZN(G24) );
  XOR2_X1 U780 ( .A(n734), .B(G119), .Z(G21) );
  XOR2_X1 U781 ( .A(n735), .B(G131), .Z(G33) );
  XNOR2_X1 U782 ( .A(G143), .B(n736), .ZN(G45) );
endmodule

