//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n460), .A2(KEYINPUT66), .B1(new_n461), .B2(new_n456), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n462), .B1(KEYINPUT66), .B2(new_n460), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT67), .ZN(G319));
  AND2_X1   g039(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(new_n468), .A3(G137), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(G101), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G125), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n467), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n472), .A2(new_n477), .ZN(G160));
  OAI221_X1 g053(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n467), .C2(G112), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n473), .A2(new_n474), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  INV_X1    g058(.A(new_n467), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n468), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n479), .B(new_n482), .C1(new_n483), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND2_X1  g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n470), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  OAI22_X1  g065(.A1(new_n480), .A2(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(new_n470), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n493), .B(new_n494), .C1(new_n473), .C2(new_n474), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n467), .A2(new_n468), .A3(new_n498), .A4(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n491), .B1(new_n497), .B2(new_n499), .ZN(G164));
  AND2_X1   g075(.A1(G75), .A2(G543), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n501), .B1(new_n504), .B2(G62), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n511), .A2(new_n512), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n507), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n511), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n514), .A2(new_n513), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n510), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n524), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n506), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT69), .B(G52), .Z(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n511), .A2(new_n532), .B1(new_n517), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  INV_X1    g110(.A(G56), .ZN(new_n536));
  INV_X1    g111(.A(G68), .ZN(new_n537));
  INV_X1    g112(.A(G543), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n525), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI221_X1 g116(.A(KEYINPUT70), .B1(new_n537), .B2(new_n538), .C1(new_n525), .C2(new_n536), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(G651), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n517), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n538), .B1(new_n508), .B2(new_n509), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n544), .A2(G81), .B1(G43), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND3_X1  g128(.A1(new_n510), .A2(G53), .A3(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n545), .A2(new_n556), .A3(G53), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n517), .A2(KEYINPUT71), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT71), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n504), .A2(new_n510), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(G91), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n525), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n558), .A2(new_n562), .A3(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n570), .B1(new_n507), .B2(new_n519), .ZN(new_n571));
  INV_X1    g146(.A(G62), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n525), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n573), .B2(new_n501), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n544), .A2(G88), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n545), .A2(G50), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT72), .A4(new_n576), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n571), .A2(new_n577), .ZN(G303));
  NAND3_X1  g153(.A1(new_n559), .A2(G87), .A3(new_n561), .ZN(new_n579));
  INV_X1    g154(.A(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n525), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(new_n545), .B2(G49), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(G288));
  AND3_X1   g158(.A1(KEYINPUT73), .A2(G73), .A3(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(KEYINPUT73), .B1(G73), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n502), .B2(new_n503), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n545), .B2(G48), .ZN(new_n591));
  OAI211_X1 g166(.A(G48), .B(G543), .C1(new_n515), .C2(new_n516), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(KEYINPUT75), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n589), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n559), .A2(G86), .A3(new_n561), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT74), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT74), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n559), .A2(new_n561), .A3(new_n597), .A4(G86), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n594), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G305));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n511), .A2(new_n601), .B1(new_n517), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G60), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n525), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n605), .B1(new_n506), .B2(new_n609), .ZN(G290));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(G301), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n559), .A2(G92), .A3(new_n561), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n525), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n618), .A2(G651), .B1(G54), .B2(new_n545), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT77), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n612), .B1(new_n622), .B2(new_n611), .ZN(G284));
  AOI21_X1  g198(.A(new_n612), .B1(new_n622), .B2(new_n611), .ZN(G321));
  NAND2_X1  g199(.A1(G299), .A2(new_n611), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n611), .B2(G168), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(new_n611), .B2(G168), .ZN(G280));
  XOR2_X1   g202(.A(KEYINPUT78), .B(G559), .Z(new_n628));
  OAI21_X1  g203(.A(new_n622), .B1(G860), .B2(new_n628), .ZN(G148));
  NOR2_X1   g204(.A1(new_n548), .A2(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n622), .A2(new_n628), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT79), .Z(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g209(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT80), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n481), .A2(G135), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT81), .ZN(new_n642));
  INV_X1    g217(.A(new_n485), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n467), .A2(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  AOI22_X1  g221(.A1(new_n643), .A2(G123), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G2096), .ZN(new_n650));
  AOI22_X1  g225(.A1(new_n649), .A2(new_n650), .B1(new_n638), .B2(new_n637), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n640), .B(new_n651), .C1(new_n650), .C2(new_n649), .ZN(G156));
  XOR2_X1   g227(.A(KEYINPUT15), .B(G2435), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT82), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT14), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n659), .B(new_n663), .Z(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G14), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT83), .ZN(new_n672));
  NOR2_X1   g247(.A1(G2072), .A2(G2078), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n444), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n670), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(KEYINPUT17), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n675), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n670), .B(new_n671), .C1(new_n444), .C2(new_n673), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT18), .Z(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n672), .A3(new_n670), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2096), .B(G2100), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1971), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n686), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n686), .B2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT84), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n702), .A2(new_n705), .A3(new_n703), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(G229));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G6), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n599), .B2(new_n710), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n710), .A2(G23), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G288), .B2(G16), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT33), .B(G1976), .Z(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n716), .A2(new_n718), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n710), .A2(G22), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT86), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G166), .B2(new_n710), .ZN(new_n723));
  INV_X1    g298(.A(G1971), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n714), .A2(new_n719), .A3(new_n720), .A4(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n713), .B2(new_n712), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT34), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  MUX2_X1   g305(.A(G24), .B(G290), .S(G16), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1986), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G25), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT85), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n643), .A2(G119), .ZN(new_n736));
  OAI221_X1 g311(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n467), .C2(G107), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n481), .A2(G131), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n735), .B1(new_n739), .B2(G29), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n732), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n729), .A2(new_n730), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(KEYINPUT36), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n729), .A2(new_n746), .A3(new_n730), .A4(new_n743), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT99), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n710), .A2(G20), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT23), .ZN(new_n751));
  INV_X1    g326(.A(G299), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n710), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT98), .B(G1956), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT26), .Z(new_n757));
  INV_X1    g332(.A(G129), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n485), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n481), .A2(G141), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n470), .A2(G105), .A3(G2104), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(new_n733), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n733), .B2(G32), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT31), .B(G11), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT94), .B(G28), .Z(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(KEYINPUT30), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(KEYINPUT30), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(new_n733), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n768), .B1(new_n770), .B2(new_n772), .C1(new_n648), .C2(new_n733), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n767), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n710), .A2(G21), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G168), .B2(new_n710), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT93), .B(G1966), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n710), .A2(G5), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G171), .B2(new_n710), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT95), .B(G1961), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT24), .ZN(new_n783));
  INV_X1    g358(.A(G34), .ZN(new_n784));
  AOI21_X1  g359(.A(G29), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n783), .B2(new_n784), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G160), .B2(new_n733), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n765), .A2(new_n766), .B1(G2084), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n774), .A2(new_n778), .A3(new_n782), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G19), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n548), .B2(G16), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT88), .B(G1341), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G27), .A2(G29), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G164), .B2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT97), .B(G2078), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n787), .A2(G2084), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT96), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n793), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n733), .A2(KEYINPUT28), .A3(G26), .ZN(new_n801));
  AOI21_X1  g376(.A(KEYINPUT28), .B1(new_n733), .B2(G26), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n481), .A2(G140), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT89), .Z(new_n804));
  OR2_X1    g379(.A1(new_n467), .A2(G116), .ZN(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n643), .A2(G128), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  AOI211_X1 g384(.A(new_n801), .B(new_n802), .C1(new_n809), .C2(G29), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT90), .B(G2067), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n733), .A2(G35), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G162), .B2(new_n733), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT29), .B(G2090), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n810), .A2(new_n811), .ZN(new_n818));
  NOR4_X1   g393(.A1(new_n789), .A2(new_n800), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n733), .A2(G33), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n481), .A2(G139), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT91), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(new_n467), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT25), .Z(new_n826));
  NAND3_X1  g401(.A1(new_n822), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT92), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT92), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n822), .A2(new_n829), .A3(new_n824), .A4(new_n826), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n820), .B1(new_n832), .B2(new_n733), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n442), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n710), .A2(G4), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n622), .B2(new_n710), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT87), .B(G1348), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AND4_X1   g413(.A1(new_n755), .A2(new_n819), .A3(new_n834), .A4(new_n838), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n748), .A2(new_n749), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n749), .B1(new_n748), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(G311));
  NAND2_X1  g417(.A1(new_n748), .A2(new_n839), .ZN(G150));
  AOI22_X1  g418(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n506), .ZN(new_n845));
  INV_X1    g420(.A(G55), .ZN(new_n846));
  INV_X1    g421(.A(G93), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n511), .A2(new_n846), .B1(new_n517), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G860), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n622), .A2(G559), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n849), .A2(new_n543), .A3(new_n546), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n849), .B1(new_n543), .B2(new_n546), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n855), .B(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n850), .B1(new_n860), .B2(KEYINPUT39), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n852), .B1(new_n861), .B2(new_n862), .ZN(G145));
  NAND2_X1  g438(.A1(new_n497), .A2(new_n499), .ZN(new_n864));
  INV_X1    g439(.A(new_n491), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n763), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n831), .B2(KEYINPUT101), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n870));
  AOI211_X1 g445(.A(new_n870), .B(new_n763), .C1(new_n828), .C2(new_n830), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n866), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n868), .A2(new_n871), .A3(G164), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n873), .A2(new_n874), .A3(new_n809), .ZN(new_n875));
  INV_X1    g450(.A(new_n809), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n869), .A2(new_n872), .A3(new_n866), .ZN(new_n877));
  OAI21_X1  g452(.A(G164), .B1(new_n868), .B2(new_n871), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI22_X1  g454(.A1(new_n643), .A2(G130), .B1(new_n481), .B2(G142), .ZN(new_n880));
  OAI221_X1 g455(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n467), .C2(G118), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n636), .ZN(new_n883));
  INV_X1    g458(.A(new_n739), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  OAI22_X1  g460(.A1(new_n875), .A2(new_n879), .B1(KEYINPUT102), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n809), .B1(new_n873), .B2(new_n874), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n877), .A2(new_n876), .A3(new_n878), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n885), .A2(KEYINPUT102), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n648), .B(G160), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(G162), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n886), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n885), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n875), .B2(new_n879), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n887), .A2(new_n888), .A3(new_n885), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n892), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n900), .B(new_n901), .ZN(G395));
  XNOR2_X1  g477(.A(new_n631), .B(new_n859), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n620), .A2(G299), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n615), .A2(new_n752), .A3(new_n619), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n908), .A2(KEYINPUT104), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(KEYINPUT41), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n904), .A2(new_n911), .A3(new_n905), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n908), .B(KEYINPUT104), .C1(new_n903), .C2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(G288), .B(KEYINPUT105), .ZN(new_n916));
  XNOR2_X1  g491(.A(G290), .B(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n599), .A2(G166), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n599), .A2(G166), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT106), .B1(new_n918), .B2(new_n919), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n917), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n916), .A2(G290), .ZN(new_n925));
  NAND2_X1  g500(.A1(G290), .A2(new_n916), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n925), .A2(new_n920), .A3(new_n921), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT42), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n909), .A2(new_n915), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n909), .B2(new_n915), .ZN(new_n931));
  OAI21_X1  g506(.A(G868), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(G868), .B2(new_n849), .ZN(G295));
  OAI21_X1  g508(.A(new_n932), .B1(G868), .B2(new_n849), .ZN(G331));
  AND2_X1   g509(.A1(new_n924), .A2(new_n927), .ZN(new_n935));
  NAND2_X1  g510(.A1(G171), .A2(G168), .ZN(new_n936));
  OAI22_X1  g511(.A1(new_n531), .A2(new_n534), .B1(new_n524), .B2(new_n528), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n856), .ZN(new_n940));
  INV_X1    g515(.A(new_n857), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n938), .B1(new_n856), .B2(new_n857), .ZN(new_n943));
  AND4_X1   g518(.A1(new_n904), .A2(new_n942), .A3(new_n905), .A4(new_n943), .ZN(new_n944));
  NOR4_X1   g519(.A1(new_n856), .A2(new_n938), .A3(new_n857), .A4(KEYINPUT107), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n858), .B2(new_n939), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n943), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n944), .B1(new_n948), .B2(new_n913), .ZN(new_n949));
  AOI21_X1  g524(.A(G37), .B1(new_n935), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n928), .B1(new_n949), .B2(KEYINPUT108), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n953));
  AOI211_X1 g528(.A(new_n953), .B(new_n944), .C1(new_n948), .C2(new_n913), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n950), .B(new_n951), .C1(new_n952), .C2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n955), .A2(KEYINPUT44), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n904), .A2(new_n957), .A3(new_n911), .A4(new_n905), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n910), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n912), .A2(KEYINPUT109), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n959), .A2(new_n960), .B1(new_n943), .B2(new_n942), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n945), .A2(new_n947), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n962), .A2(new_n907), .A3(new_n943), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n928), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n950), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT111), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n965), .A2(KEYINPUT111), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n956), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n950), .B1(new_n952), .B2(new_n954), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n964), .A2(new_n951), .A3(new_n950), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT110), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n976));
  AOI211_X1 g551(.A(new_n976), .B(KEYINPUT44), .C1(new_n971), .C2(new_n972), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n969), .B1(new_n975), .B2(new_n977), .ZN(G397));
  INV_X1    g553(.A(KEYINPUT127), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(G164), .B2(G1384), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G40), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n472), .A2(new_n983), .A3(new_n477), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G2067), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n809), .B(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n763), .B(G1996), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n739), .B(new_n741), .Z(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(G290), .B(new_n698), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n985), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n475), .A2(new_n476), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n484), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n995), .A2(G40), .A3(new_n471), .A4(new_n469), .ZN(new_n996));
  NOR2_X1   g571(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n996), .B1(new_n866), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G2084), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n866), .A2(KEYINPUT45), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n984), .A3(new_n981), .ZN(new_n1006));
  INV_X1    g581(.A(G1966), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n998), .A2(KEYINPUT114), .A3(new_n999), .A4(new_n1000), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1003), .A2(new_n1008), .A3(G168), .A4(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n1011));
  AND2_X1   g586(.A1(KEYINPUT121), .A2(G8), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1003), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(G8), .A3(G286), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1011), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT62), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT51), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT62), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(new_n1021), .A3(new_n1015), .A4(new_n1013), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n571), .A2(new_n577), .A3(G8), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT55), .ZN(new_n1024));
  INV_X1    g599(.A(G2090), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n866), .B2(new_n1004), .ZN(new_n1027));
  INV_X1    g602(.A(new_n997), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n984), .B1(G164), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1025), .A2(new_n1030), .B1(new_n1006), .B2(new_n724), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1024), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n866), .A2(new_n984), .A3(new_n1004), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n579), .A2(G1976), .A3(new_n582), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(G8), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT52), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1039), .A2(new_n1034), .A3(G8), .A4(new_n1035), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n592), .A2(KEYINPUT75), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n545), .A2(new_n590), .A3(G48), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n584), .A2(new_n585), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n525), .B2(new_n587), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1042), .A2(new_n1043), .B1(new_n1045), .B2(G651), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n544), .A2(G86), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n696), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1048), .B1(new_n599), .B2(new_n696), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT49), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1034), .A2(G8), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n596), .A2(new_n598), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(new_n696), .A3(new_n1046), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1048), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1051), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1041), .B1(new_n1050), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1006), .A2(new_n724), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n998), .A2(new_n1025), .A3(new_n1000), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1023), .B(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(G8), .A3(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1005), .A2(new_n981), .A3(new_n443), .A4(new_n984), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n998), .A2(new_n1000), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT122), .B(G1961), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1065), .A2(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1066), .A2(G2078), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1005), .A2(new_n981), .A3(new_n984), .A4(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(G301), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  AND4_X1   g647(.A1(new_n1033), .A2(new_n1058), .A3(new_n1064), .A4(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1018), .A2(new_n1022), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT63), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1058), .A2(new_n1033), .A3(new_n1064), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1014), .A2(G8), .A3(G168), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1031), .A2(new_n1024), .A3(new_n1032), .ZN(new_n1079));
  NOR2_X1   g654(.A1(G164), .A2(G1384), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1032), .B1(new_n1080), .B2(new_n984), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1049), .B2(KEYINPUT49), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1053), .A2(KEYINPUT49), .A3(new_n1054), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1037), .B(new_n1040), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1079), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT115), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1061), .A2(new_n1087), .A3(G8), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1024), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1077), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1085), .A2(new_n1089), .A3(KEYINPUT63), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1078), .A2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1051), .B(KEYINPUT112), .ZN(new_n1093));
  NOR2_X1   g668(.A1(G288), .A2(G1976), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1093), .B1(new_n1095), .B2(new_n1053), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1084), .A2(new_n1064), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT113), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1057), .A2(new_n1050), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1041), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1032), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1063), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1100), .A2(new_n1094), .B1(new_n696), .B2(new_n599), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1099), .B(new_n1103), .C1(new_n1104), .C2(new_n1093), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1098), .A2(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1074), .A2(new_n1092), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1005), .A2(new_n981), .A3(new_n984), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(G1956), .B1(new_n998), .B2(new_n1000), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1108), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT118), .B(new_n1110), .C1(new_n1030), .C2(G1956), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n1115));
  XNOR2_X1  g690(.A(G299), .B(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1348), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT117), .B1(new_n1034), .B2(G2067), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT117), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1080), .A2(new_n1122), .A3(new_n986), .A4(new_n984), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1118), .B1(new_n1124), .B2(new_n620), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1116), .B(new_n1110), .C1(new_n1030), .C2(G1956), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1120), .A2(new_n1121), .A3(KEYINPUT60), .A4(new_n1123), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1131));
  INV_X1    g706(.A(new_n620), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1128), .A2(new_n1129), .A3(new_n620), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1124), .A2(KEYINPUT60), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1126), .A2(KEYINPUT61), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1118), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1117), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1126), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n1144));
  INV_X1    g719(.A(G1996), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1005), .A2(new_n981), .A3(new_n1145), .A4(new_n984), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT58), .B(G1341), .Z(new_n1147));
  AOI22_X1  g722(.A1(new_n1146), .A2(KEYINPUT119), .B1(new_n1034), .B2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1005), .A2(new_n981), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(new_n1145), .A4(new_n984), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1144), .B1(new_n1152), .B2(new_n548), .ZN(new_n1153));
  AOI211_X1 g728(.A(KEYINPUT59), .B(new_n547), .C1(new_n1148), .C2(new_n1151), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1139), .B(new_n1143), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1127), .B1(new_n1137), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1157), .A2(new_n1158), .A3(G301), .A4(new_n1071), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1159), .A2(KEYINPUT54), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n472), .B(KEYINPUT123), .Z(new_n1161));
  NOR4_X1   g736(.A1(new_n477), .A2(new_n1066), .A3(new_n983), .A4(G2078), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1161), .A2(new_n1005), .A3(new_n981), .A4(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1157), .A2(new_n1163), .A3(new_n1158), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1164), .A2(new_n1165), .A3(G171), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1165), .B1(new_n1164), .B2(G171), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1160), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g745(.A(KEYINPUT125), .B(new_n1160), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1020), .A2(new_n1015), .A3(new_n1013), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1076), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT54), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1164), .A2(G171), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1175), .B1(new_n1176), .B2(new_n1072), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1173), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1156), .A2(new_n1172), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n993), .B1(new_n1107), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n991), .A2(new_n985), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT48), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n985), .A2(G290), .A3(G1986), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT126), .Z(new_n1185));
  AOI21_X1  g760(.A(new_n1182), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1186), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n985), .B1(new_n987), .B2(new_n763), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT46), .B1(new_n985), .B2(G1996), .ZN(new_n1189));
  OR3_X1    g764(.A1(new_n985), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT47), .Z(new_n1192));
  NAND2_X1  g767(.A1(new_n884), .A2(new_n741), .ZN(new_n1193));
  OAI22_X1  g768(.A1(new_n989), .A2(new_n1193), .B1(G2067), .B2(new_n809), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1194), .A2(new_n984), .A3(new_n982), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1187), .A2(new_n1192), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n979), .B1(new_n1181), .B2(new_n1196), .ZN(new_n1197));
  AND3_X1   g772(.A1(new_n1187), .A2(new_n1192), .A3(new_n1195), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1074), .A2(new_n1092), .A3(new_n1106), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1152), .A2(new_n548), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1152), .A2(new_n1144), .A3(new_n548), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI22_X1  g778(.A1(new_n1118), .A2(new_n1138), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1204));
  OAI211_X1 g779(.A(new_n1203), .B(new_n1204), .C1(new_n1136), .C2(new_n1135), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1178), .B1(new_n1205), .B2(new_n1127), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1199), .B1(new_n1172), .B2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g782(.A(KEYINPUT127), .B(new_n1198), .C1(new_n1207), .C2(new_n993), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1197), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g784(.A(new_n463), .B(new_n683), .C1(new_n667), .C2(new_n668), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1211), .B1(new_n707), .B2(new_n708), .ZN(new_n1212));
  NAND3_X1  g786(.A1(new_n1212), .A2(new_n900), .A3(new_n973), .ZN(G225));
  INV_X1    g787(.A(G225), .ZN(G308));
endmodule


