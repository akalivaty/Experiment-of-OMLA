

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745;

  INV_X1 U372 ( .A(n691), .ZN(n352) );
  INV_X1 U373 ( .A(KEYINPUT64), .ZN(n354) );
  XNOR2_X1 U374 ( .A(n379), .B(KEYINPUT113), .ZN(n738) );
  XNOR2_X1 U375 ( .A(n400), .B(n360), .ZN(n415) );
  AND2_X1 U376 ( .A1(n667), .A2(n547), .ZN(n548) );
  XNOR2_X1 U377 ( .A(n549), .B(KEYINPUT1), .ZN(n670) );
  XNOR2_X1 U378 ( .A(n522), .B(KEYINPUT19), .ZN(n552) );
  BUF_X1 U379 ( .A(G113), .Z(n355) );
  INV_X1 U380 ( .A(n430), .ZN(n432) );
  XNOR2_X1 U381 ( .A(G119), .B(KEYINPUT3), .ZN(n431) );
  INV_X2 U382 ( .A(G953), .ZN(n730) );
  NAND2_X2 U383 ( .A1(n439), .A2(n651), .ZN(n440) );
  AND2_X4 U384 ( .A1(n353), .A2(n352), .ZN(n712) );
  XNOR2_X2 U385 ( .A(n612), .B(n354), .ZN(n353) );
  XNOR2_X2 U386 ( .A(n449), .B(n426), .ZN(n392) );
  NOR2_X1 U387 ( .A1(G953), .A2(G237), .ZN(n492) );
  INV_X1 U388 ( .A(n670), .ZN(n403) );
  NAND2_X1 U389 ( .A1(n589), .A2(n527), .ZN(n669) );
  AND2_X1 U390 ( .A1(n399), .A2(n365), .ZN(n418) );
  NOR2_X1 U391 ( .A1(n661), .A2(n371), .ZN(n562) );
  AND2_X1 U392 ( .A1(n550), .A2(n410), .ZN(n551) );
  NOR2_X1 U393 ( .A1(n648), .A2(n654), .ZN(n561) );
  XNOR2_X2 U394 ( .A(G101), .B(G113), .ZN(n430) );
  XNOR2_X2 U395 ( .A(n458), .B(G472), .ZN(n537) );
  INV_X1 U396 ( .A(KEYINPUT15), .ZN(n434) );
  NAND2_X1 U397 ( .A1(n700), .A2(n610), .ZN(n437) );
  XOR2_X1 U398 ( .A(G116), .B(G107), .Z(n503) );
  XNOR2_X1 U399 ( .A(n429), .B(n455), .ZN(n508) );
  INV_X1 U400 ( .A(G134), .ZN(n455) );
  XOR2_X1 U401 ( .A(G122), .B(G104), .Z(n487) );
  NOR2_X1 U402 ( .A1(n376), .A2(n373), .ZN(n372) );
  INV_X1 U403 ( .A(KEYINPUT46), .ZN(n374) );
  XNOR2_X1 U404 ( .A(G143), .B(G128), .ZN(n429) );
  XOR2_X1 U405 ( .A(G146), .B(G125), .Z(n472) );
  XNOR2_X1 U406 ( .A(KEYINPUT67), .B(n529), .ZN(n547) );
  XNOR2_X1 U407 ( .A(n409), .B(n408), .ZN(n407) );
  XNOR2_X1 U408 ( .A(G128), .B(KEYINPUT94), .ZN(n409) );
  XNOR2_X1 U409 ( .A(G119), .B(G110), .ZN(n408) );
  XNOR2_X1 U410 ( .A(n406), .B(KEYINPUT23), .ZN(n405) );
  XNOR2_X1 U411 ( .A(KEYINPUT24), .B(KEYINPUT78), .ZN(n406) );
  INV_X1 U412 ( .A(KEYINPUT103), .ZN(n504) );
  XOR2_X1 U413 ( .A(G131), .B(G140), .Z(n494) );
  XNOR2_X1 U414 ( .A(n355), .B(G143), .ZN(n490) );
  XNOR2_X1 U415 ( .A(KEYINPUT101), .B(KEYINPUT11), .ZN(n488) );
  NOR2_X1 U416 ( .A1(n608), .A2(n424), .ZN(n423) );
  NAND2_X1 U417 ( .A1(n417), .A2(KEYINPUT79), .ZN(n416) );
  XNOR2_X1 U418 ( .A(n387), .B(n386), .ZN(n390) );
  XNOR2_X1 U419 ( .A(KEYINPUT71), .B(KEYINPUT17), .ZN(n387) );
  NAND2_X1 U420 ( .A1(n730), .A2(G224), .ZN(n386) );
  INV_X1 U421 ( .A(n429), .ZN(n391) );
  INV_X1 U422 ( .A(n472), .ZN(n412) );
  XNOR2_X1 U423 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n427) );
  XNOR2_X1 U424 ( .A(n558), .B(n557), .ZN(n573) );
  XNOR2_X1 U425 ( .A(n512), .B(n511), .ZN(n564) );
  XNOR2_X1 U426 ( .A(n398), .B(n397), .ZN(n565) );
  XNOR2_X1 U427 ( .A(n499), .B(G475), .ZN(n397) );
  NOR2_X1 U428 ( .A1(n626), .A2(G902), .ZN(n398) );
  NOR2_X1 U429 ( .A1(n572), .A2(n563), .ZN(n377) );
  INV_X1 U430 ( .A(KEYINPUT44), .ZN(n413) );
  AND2_X1 U431 ( .A1(n525), .A2(G953), .ZN(n385) );
  INV_X1 U432 ( .A(KEYINPUT108), .ZN(n384) );
  XOR2_X1 U433 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n451) );
  XOR2_X1 U434 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n489) );
  NOR2_X1 U435 ( .A1(n422), .A2(KEYINPUT79), .ZN(n421) );
  XNOR2_X1 U436 ( .A(n508), .B(n456), .ZN(n728) );
  XNOR2_X1 U437 ( .A(KEYINPUT4), .B(G131), .ZN(n456) );
  XNOR2_X1 U438 ( .A(n380), .B(n359), .ZN(n441) );
  XNOR2_X1 U439 ( .A(KEYINPUT14), .B(KEYINPUT91), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n396), .B(n361), .ZN(n617) );
  NAND2_X1 U441 ( .A1(n378), .A2(n372), .ZN(n396) );
  OR2_X1 U442 ( .A1(G237), .A2(G902), .ZN(n438) );
  XNOR2_X1 U443 ( .A(n484), .B(n483), .ZN(n658) );
  NAND2_X1 U444 ( .A1(n403), .A2(n402), .ZN(n484) );
  NOR2_X1 U445 ( .A1(n591), .A2(n669), .ZN(n402) );
  XNOR2_X1 U446 ( .A(n381), .B(KEYINPUT73), .ZN(n540) );
  NAND2_X1 U447 ( .A1(n383), .A2(n382), .ZN(n381) );
  INV_X1 U448 ( .A(n526), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n383) );
  INV_X1 U450 ( .A(G902), .ZN(n510) );
  INV_X1 U451 ( .A(n669), .ZN(n594) );
  XNOR2_X1 U452 ( .A(n728), .B(G146), .ZN(n466) );
  XNOR2_X1 U453 ( .A(G110), .B(G107), .ZN(n461) );
  XNOR2_X1 U454 ( .A(G104), .B(G101), .ZN(n462) );
  AND2_X1 U455 ( .A1(n547), .A2(n530), .ZN(n531) );
  BUF_X1 U456 ( .A(n537), .Z(n667) );
  XNOR2_X1 U457 ( .A(n407), .B(n405), .ZN(n476) );
  XNOR2_X1 U458 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U459 ( .A(n498), .B(n497), .ZN(n626) );
  NAND2_X1 U460 ( .A1(n418), .A2(n416), .ZN(n420) );
  XNOR2_X1 U461 ( .A(n389), .B(n411), .ZN(n388) );
  XNOR2_X1 U462 ( .A(n428), .B(n412), .ZN(n411) );
  XNOR2_X1 U463 ( .A(n391), .B(n390), .ZN(n389) );
  XOR2_X1 U464 ( .A(KEYINPUT40), .B(n559), .Z(n740) );
  XOR2_X1 U465 ( .A(n472), .B(KEYINPUT10), .Z(n356) );
  AND2_X1 U466 ( .A1(n640), .A2(n531), .ZN(n357) );
  XNOR2_X1 U467 ( .A(n468), .B(n467), .ZN(n549) );
  INV_X1 U468 ( .A(n549), .ZN(n410) );
  OR2_X1 U469 ( .A1(n571), .A2(n570), .ZN(n358) );
  AND2_X1 U470 ( .A1(n542), .A2(n541), .ZN(n556) );
  AND2_X1 U471 ( .A1(G234), .A2(G237), .ZN(n359) );
  XOR2_X1 U472 ( .A(n515), .B(KEYINPUT72), .Z(n360) );
  XOR2_X1 U473 ( .A(KEYINPUT66), .B(KEYINPUT48), .Z(n361) );
  XOR2_X1 U474 ( .A(n626), .B(n625), .Z(n362) );
  XOR2_X1 U475 ( .A(n621), .B(n620), .Z(n363) );
  XNOR2_X1 U476 ( .A(n700), .B(n699), .ZN(n364) );
  NOR2_X1 U477 ( .A1(n423), .A2(n611), .ZN(n365) );
  INV_X1 U478 ( .A(KEYINPUT79), .ZN(n424) );
  NOR2_X1 U479 ( .A1(n730), .A2(G952), .ZN(n716) );
  INV_X1 U480 ( .A(n716), .ZN(n366) );
  AND2_X2 U481 ( .A1(n367), .A2(n366), .ZN(n624) );
  XNOR2_X1 U482 ( .A(n622), .B(n363), .ZN(n367) );
  AND2_X2 U483 ( .A1(n368), .A2(n366), .ZN(n628) );
  XNOR2_X1 U484 ( .A(n627), .B(n362), .ZN(n368) );
  AND2_X2 U485 ( .A1(n369), .A2(n366), .ZN(n702) );
  XNOR2_X1 U486 ( .A(n701), .B(n364), .ZN(n369) );
  NAND2_X1 U487 ( .A1(n370), .A2(n425), .ZN(n419) );
  NAND2_X1 U488 ( .A1(n617), .A2(n580), .ZN(n370) );
  NOR2_X1 U489 ( .A1(n720), .A2(n370), .ZN(n689) );
  XNOR2_X1 U490 ( .A(n370), .B(n732), .ZN(n731) );
  INV_X1 U491 ( .A(n551), .ZN(n371) );
  XNOR2_X1 U492 ( .A(n375), .B(n374), .ZN(n373) );
  NOR2_X1 U493 ( .A1(n743), .A2(n740), .ZN(n375) );
  NAND2_X1 U494 ( .A1(n377), .A2(n358), .ZN(n376) );
  INV_X1 U495 ( .A(n738), .ZN(n378) );
  NAND2_X1 U496 ( .A1(n404), .A2(n535), .ZN(n379) );
  XNOR2_X2 U497 ( .A(n717), .B(n388), .ZN(n700) );
  XNOR2_X2 U498 ( .A(n392), .B(n433), .ZN(n717) );
  XNOR2_X2 U499 ( .A(n432), .B(n431), .ZN(n449) );
  XNOR2_X2 U500 ( .A(n393), .B(n607), .ZN(n613) );
  NAND2_X1 U501 ( .A1(n394), .A2(n605), .ZN(n393) );
  XNOR2_X1 U502 ( .A(n395), .B(n413), .ZN(n394) );
  NAND2_X1 U503 ( .A1(n414), .A2(n415), .ZN(n395) );
  NAND2_X1 U504 ( .A1(n613), .A2(n421), .ZN(n399) );
  INV_X1 U505 ( .A(n415), .ZN(n587) );
  NAND2_X1 U506 ( .A1(n401), .A2(n545), .ZN(n400) );
  XNOR2_X1 U507 ( .A(n486), .B(n485), .ZN(n401) );
  XNOR2_X1 U508 ( .A(n534), .B(KEYINPUT36), .ZN(n404) );
  XNOR2_X2 U509 ( .A(n478), .B(n479), .ZN(n589) );
  NAND2_X1 U510 ( .A1(n410), .A2(n594), .ZN(n599) );
  NAND2_X1 U511 ( .A1(n573), .A2(n640), .ZN(n559) );
  NOR2_X1 U512 ( .A1(n744), .A2(n586), .ZN(n414) );
  INV_X1 U513 ( .A(n613), .ZN(n417) );
  NAND2_X1 U514 ( .A1(n420), .A2(n419), .ZN(n612) );
  INV_X1 U515 ( .A(n608), .ZN(n422) );
  INV_X1 U516 ( .A(n611), .ZN(n425) );
  XNOR2_X1 U517 ( .A(G110), .B(KEYINPUT16), .ZN(n426) );
  INV_X1 U518 ( .A(KEYINPUT34), .ZN(n485) );
  XNOR2_X1 U519 ( .A(n507), .B(n506), .ZN(n509) );
  XNOR2_X1 U520 ( .A(n427), .B(KEYINPUT90), .ZN(n428) );
  XNOR2_X1 U521 ( .A(n487), .B(n503), .ZN(n433) );
  XNOR2_X1 U522 ( .A(G902), .B(KEYINPUT89), .ZN(n435) );
  XNOR2_X1 U523 ( .A(n435), .B(n434), .ZN(n610) );
  NAND2_X1 U524 ( .A1(n438), .A2(G210), .ZN(n436) );
  XNOR2_X2 U525 ( .A(n437), .B(n436), .ZN(n536) );
  INV_X1 U526 ( .A(n536), .ZN(n439) );
  NAND2_X1 U527 ( .A1(G214), .A2(n438), .ZN(n651) );
  XNOR2_X2 U528 ( .A(n440), .B(KEYINPUT84), .ZN(n522) );
  NAND2_X1 U529 ( .A1(G952), .A2(n441), .ZN(n683) );
  NOR2_X1 U530 ( .A1(G953), .A2(n683), .ZN(n526) );
  NAND2_X1 U531 ( .A1(G902), .A2(n441), .ZN(n524) );
  XOR2_X1 U532 ( .A(G898), .B(KEYINPUT92), .Z(n723) );
  NAND2_X1 U533 ( .A1(G953), .A2(n723), .ZN(n718) );
  NOR2_X1 U534 ( .A1(n524), .A2(n718), .ZN(n442) );
  NOR2_X1 U535 ( .A1(n526), .A2(n442), .ZN(n443) );
  XNOR2_X1 U536 ( .A(KEYINPUT93), .B(n443), .ZN(n444) );
  NAND2_X1 U537 ( .A1(n552), .A2(n444), .ZN(n447) );
  INV_X1 U538 ( .A(KEYINPUT86), .ZN(n445) );
  XNOR2_X1 U539 ( .A(n445), .B(KEYINPUT0), .ZN(n446) );
  XNOR2_X2 U540 ( .A(n447), .B(n446), .ZN(n518) );
  BUF_X2 U541 ( .A(n518), .Z(n601) );
  XNOR2_X1 U542 ( .A(G116), .B(KEYINPUT5), .ZN(n448) );
  XNOR2_X1 U543 ( .A(n449), .B(n448), .ZN(n454) );
  NAND2_X1 U544 ( .A1(n492), .A2(G210), .ZN(n450) );
  XNOR2_X1 U545 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U546 ( .A(n452), .B(G137), .Z(n453) );
  XNOR2_X1 U547 ( .A(n454), .B(n453), .ZN(n457) );
  XNOR2_X1 U548 ( .A(n457), .B(n466), .ZN(n621) );
  NAND2_X1 U549 ( .A1(n621), .A2(n510), .ZN(n458) );
  XNOR2_X1 U550 ( .A(n537), .B(KEYINPUT6), .ZN(n591) );
  NAND2_X1 U551 ( .A1(n730), .A2(G227), .ZN(n459) );
  XNOR2_X1 U552 ( .A(n459), .B(KEYINPUT70), .ZN(n460) );
  XNOR2_X1 U553 ( .A(G140), .B(G137), .ZN(n473) );
  XNOR2_X1 U554 ( .A(n460), .B(n473), .ZN(n464) );
  XNOR2_X1 U555 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U556 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U557 ( .A(n466), .B(n465), .ZN(n705) );
  OR2_X1 U558 ( .A1(n705), .A2(G902), .ZN(n468) );
  INV_X1 U559 ( .A(G469), .ZN(n467) );
  XOR2_X1 U560 ( .A(KEYINPUT95), .B(KEYINPUT25), .Z(n471) );
  NAND2_X1 U561 ( .A1(n610), .A2(G234), .ZN(n469) );
  XNOR2_X1 U562 ( .A(n469), .B(KEYINPUT20), .ZN(n480) );
  NAND2_X1 U563 ( .A1(G217), .A2(n480), .ZN(n470) );
  XNOR2_X1 U564 ( .A(n471), .B(n470), .ZN(n479) );
  XNOR2_X1 U565 ( .A(n356), .B(n473), .ZN(n729) );
  NAND2_X1 U566 ( .A1(G234), .A2(n730), .ZN(n474) );
  XOR2_X1 U567 ( .A(KEYINPUT8), .B(n474), .Z(n500) );
  NAND2_X1 U568 ( .A1(G221), .A2(n500), .ZN(n475) );
  XNOR2_X1 U569 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U570 ( .A(n729), .B(n477), .ZN(n713) );
  NOR2_X1 U571 ( .A1(n713), .A2(G902), .ZN(n478) );
  NAND2_X1 U572 ( .A1(G221), .A2(n480), .ZN(n482) );
  XOR2_X1 U573 ( .A(KEYINPUT21), .B(KEYINPUT96), .Z(n481) );
  XNOR2_X1 U574 ( .A(n482), .B(n481), .ZN(n527) );
  XNOR2_X1 U575 ( .A(KEYINPUT68), .B(KEYINPUT33), .ZN(n483) );
  NAND2_X1 U576 ( .A1(n601), .A2(n658), .ZN(n486) );
  XNOR2_X1 U577 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n499) );
  XOR2_X1 U578 ( .A(n356), .B(n487), .Z(n498) );
  XNOR2_X1 U579 ( .A(n489), .B(n488), .ZN(n491) );
  XNOR2_X1 U580 ( .A(n491), .B(n490), .ZN(n496) );
  NAND2_X1 U581 ( .A1(G214), .A2(n492), .ZN(n493) );
  XNOR2_X1 U582 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U583 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U584 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n502) );
  NAND2_X1 U585 ( .A1(G217), .A2(n500), .ZN(n501) );
  XNOR2_X1 U586 ( .A(n502), .B(n501), .ZN(n507) );
  XNOR2_X1 U587 ( .A(G122), .B(n503), .ZN(n505) );
  XNOR2_X1 U588 ( .A(n509), .B(n508), .ZN(n710) );
  NAND2_X1 U589 ( .A1(n710), .A2(n510), .ZN(n512) );
  XOR2_X1 U590 ( .A(KEYINPUT104), .B(G478), .Z(n511) );
  INV_X1 U591 ( .A(n564), .ZN(n513) );
  NAND2_X1 U592 ( .A1(n565), .A2(n513), .ZN(n514) );
  XNOR2_X1 U593 ( .A(n514), .B(KEYINPUT107), .ZN(n545) );
  XNOR2_X1 U594 ( .A(KEYINPUT82), .B(KEYINPUT35), .ZN(n515) );
  XOR2_X1 U595 ( .A(G122), .B(n587), .Z(G24) );
  INV_X1 U596 ( .A(n527), .ZN(n662) );
  INV_X1 U597 ( .A(n565), .ZN(n516) );
  NAND2_X1 U598 ( .A1(n564), .A2(n516), .ZN(n654) );
  NOR2_X1 U599 ( .A1(n662), .A2(n654), .ZN(n517) );
  NAND2_X1 U600 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U601 ( .A(n519), .B(KEYINPUT22), .ZN(n584) );
  BUF_X1 U602 ( .A(n584), .Z(n588) );
  NOR2_X1 U603 ( .A1(n667), .A2(n589), .ZN(n520) );
  NAND2_X1 U604 ( .A1(n670), .A2(n520), .ZN(n521) );
  NOR2_X1 U605 ( .A1(n588), .A2(n521), .ZN(n586) );
  XOR2_X1 U606 ( .A(G110), .B(n586), .Z(G12) );
  BUF_X1 U607 ( .A(n522), .Z(n533) );
  NAND2_X1 U608 ( .A1(n565), .A2(n564), .ZN(n523) );
  XNOR2_X2 U609 ( .A(n523), .B(KEYINPUT105), .ZN(n640) );
  NOR2_X1 U610 ( .A1(G900), .A2(n524), .ZN(n525) );
  NOR2_X1 U611 ( .A1(n540), .A2(n589), .ZN(n528) );
  NAND2_X1 U612 ( .A1(n528), .A2(n527), .ZN(n529) );
  INV_X1 U613 ( .A(n591), .ZN(n530) );
  XNOR2_X1 U614 ( .A(n357), .B(KEYINPUT109), .ZN(n576) );
  XNOR2_X1 U615 ( .A(n576), .B(KEYINPUT112), .ZN(n532) );
  NOR2_X1 U616 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U617 ( .A(n670), .B(KEYINPUT88), .ZN(n582) );
  INV_X1 U618 ( .A(n582), .ZN(n535) );
  BUF_X2 U619 ( .A(n536), .Z(n578) );
  NAND2_X1 U620 ( .A1(n537), .A2(n651), .ZN(n538) );
  XNOR2_X1 U621 ( .A(KEYINPUT30), .B(n538), .ZN(n539) );
  NOR2_X1 U622 ( .A1(n540), .A2(n539), .ZN(n542) );
  INV_X1 U623 ( .A(n599), .ZN(n541) );
  INV_X1 U624 ( .A(n556), .ZN(n543) );
  NOR2_X1 U625 ( .A1(n578), .A2(n543), .ZN(n544) );
  NAND2_X1 U626 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U627 ( .A(KEYINPUT110), .B(n546), .ZN(n742) );
  XNOR2_X1 U628 ( .A(KEYINPUT28), .B(n548), .ZN(n550) );
  AND2_X1 U629 ( .A1(n552), .A2(n551), .ZN(n638) );
  INV_X1 U630 ( .A(n638), .ZN(n553) );
  NAND2_X1 U631 ( .A1(KEYINPUT47), .A2(n553), .ZN(n554) );
  NAND2_X1 U632 ( .A1(KEYINPUT77), .A2(n554), .ZN(n555) );
  NAND2_X1 U633 ( .A1(n742), .A2(n555), .ZN(n563) );
  XNOR2_X2 U634 ( .A(n578), .B(KEYINPUT38), .ZN(n652) );
  NAND2_X1 U635 ( .A1(n556), .A2(n652), .ZN(n558) );
  XOR2_X1 U636 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n557) );
  NAND2_X1 U637 ( .A1(n652), .A2(n651), .ZN(n560) );
  XOR2_X1 U638 ( .A(KEYINPUT111), .B(n560), .Z(n648) );
  XNOR2_X1 U639 ( .A(n561), .B(KEYINPUT41), .ZN(n661) );
  XNOR2_X1 U640 ( .A(n562), .B(KEYINPUT42), .ZN(n743) );
  NOR2_X1 U641 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U642 ( .A(n566), .B(KEYINPUT106), .ZN(n644) );
  NOR2_X1 U643 ( .A1(n644), .A2(n640), .ZN(n649) );
  NOR2_X1 U644 ( .A1(KEYINPUT47), .A2(n649), .ZN(n567) );
  NAND2_X1 U645 ( .A1(n638), .A2(n567), .ZN(n568) );
  XNOR2_X1 U646 ( .A(KEYINPUT69), .B(n568), .ZN(n572) );
  INV_X1 U647 ( .A(KEYINPUT47), .ZN(n571) );
  NOR2_X1 U648 ( .A1(n638), .A2(KEYINPUT77), .ZN(n569) );
  NOR2_X1 U649 ( .A1(n649), .A2(n569), .ZN(n570) );
  NAND2_X1 U650 ( .A1(n573), .A2(n644), .ZN(n574) );
  XNOR2_X1 U651 ( .A(n574), .B(KEYINPUT114), .ZN(n741) );
  NAND2_X1 U652 ( .A1(n670), .A2(n651), .ZN(n575) );
  OR2_X1 U653 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U654 ( .A(n577), .B(KEYINPUT43), .ZN(n579) );
  NAND2_X1 U655 ( .A1(n579), .A2(n578), .ZN(n647) );
  AND2_X1 U656 ( .A1(n741), .A2(n647), .ZN(n580) );
  INV_X1 U657 ( .A(n589), .ZN(n663) );
  NAND2_X1 U658 ( .A1(n591), .A2(n663), .ZN(n581) );
  OR2_X1 U659 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U660 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U661 ( .A(n585), .B(KEYINPUT32), .ZN(n744) );
  INV_X1 U662 ( .A(n588), .ZN(n593) );
  AND2_X1 U663 ( .A1(n670), .A2(n589), .ZN(n590) );
  AND2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n629) );
  NAND2_X1 U666 ( .A1(n667), .A2(n594), .ZN(n595) );
  OR2_X1 U667 ( .A1(n670), .A2(n595), .ZN(n674) );
  INV_X1 U668 ( .A(n674), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n601), .A2(n596), .ZN(n598) );
  XOR2_X1 U670 ( .A(KEYINPUT99), .B(KEYINPUT31), .Z(n597) );
  XNOR2_X1 U671 ( .A(n598), .B(n597), .ZN(n643) );
  NOR2_X1 U672 ( .A1(n667), .A2(n599), .ZN(n600) );
  AND2_X1 U673 ( .A1(n601), .A2(n600), .ZN(n631) );
  OR2_X1 U674 ( .A1(n643), .A2(n631), .ZN(n603) );
  INV_X1 U675 ( .A(n649), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U677 ( .A1(n629), .A2(n604), .ZN(n605) );
  INV_X1 U678 ( .A(KEYINPUT81), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT45), .ZN(n607) );
  INV_X1 U680 ( .A(n610), .ZN(n608) );
  INV_X1 U681 ( .A(KEYINPUT2), .ZN(n609) );
  NOR2_X1 U682 ( .A1(n610), .A2(n609), .ZN(n611) );
  BUF_X1 U683 ( .A(n613), .Z(n687) );
  NAND2_X1 U684 ( .A1(n741), .A2(KEYINPUT2), .ZN(n614) );
  XOR2_X1 U685 ( .A(KEYINPUT74), .B(n614), .Z(n615) );
  AND2_X1 U686 ( .A1(n615), .A2(n647), .ZN(n616) );
  AND2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n618) );
  AND2_X1 U688 ( .A1(n687), .A2(n618), .ZN(n691) );
  NAND2_X1 U689 ( .A1(n712), .A2(G472), .ZN(n622) );
  XNOR2_X1 U690 ( .A(KEYINPUT87), .B(KEYINPUT62), .ZN(n620) );
  XNOR2_X1 U691 ( .A(KEYINPUT115), .B(KEYINPUT63), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n624), .B(n623), .ZN(G57) );
  NAND2_X1 U693 ( .A1(n712), .A2(G475), .ZN(n627) );
  XNOR2_X1 U694 ( .A(KEYINPUT65), .B(KEYINPUT59), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n628), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U696 ( .A(G101), .B(n629), .ZN(G3) );
  NAND2_X1 U697 ( .A1(n631), .A2(n640), .ZN(n630) );
  XNOR2_X1 U698 ( .A(n630), .B(G104), .ZN(G6) );
  XOR2_X1 U699 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n633) );
  NAND2_X1 U700 ( .A1(n631), .A2(n644), .ZN(n632) );
  XNOR2_X1 U701 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U702 ( .A(G107), .B(n634), .ZN(G9) );
  XOR2_X1 U703 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n636) );
  NAND2_X1 U704 ( .A1(n638), .A2(n644), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U706 ( .A(G128), .B(n637), .ZN(G30) );
  NAND2_X1 U707 ( .A1(n638), .A2(n640), .ZN(n639) );
  XNOR2_X1 U708 ( .A(n639), .B(G146), .ZN(G48) );
  XOR2_X1 U709 ( .A(n355), .B(KEYINPUT117), .Z(n642) );
  NAND2_X1 U710 ( .A1(n643), .A2(n640), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n642), .B(n641), .ZN(G15) );
  NAND2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U713 ( .A(n645), .B(KEYINPUT118), .ZN(n646) );
  XNOR2_X1 U714 ( .A(G116), .B(n646), .ZN(G18) );
  XNOR2_X1 U715 ( .A(G140), .B(n647), .ZN(G42) );
  NOR2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U717 ( .A(KEYINPUT123), .B(n650), .Z(n657) );
  NOR2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U719 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U720 ( .A(KEYINPUT122), .B(n655), .ZN(n656) );
  NOR2_X1 U721 ( .A1(n657), .A2(n656), .ZN(n659) );
  INV_X1 U722 ( .A(n658), .ZN(n684) );
  NOR2_X1 U723 ( .A1(n659), .A2(n684), .ZN(n660) );
  XNOR2_X1 U724 ( .A(n660), .B(KEYINPUT124), .ZN(n680) );
  XOR2_X1 U725 ( .A(KEYINPUT121), .B(KEYINPUT51), .Z(n677) );
  XOR2_X1 U726 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n665) );
  NAND2_X1 U727 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U728 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X1 U729 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U730 ( .A(KEYINPUT120), .B(n668), .ZN(n673) );
  NAND2_X1 U731 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U732 ( .A(n671), .B(KEYINPUT50), .ZN(n672) );
  NAND2_X1 U733 ( .A1(n673), .A2(n672), .ZN(n675) );
  NAND2_X1 U734 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U735 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X1 U736 ( .A1(n661), .A2(n678), .ZN(n679) );
  NOR2_X1 U737 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U738 ( .A(n681), .B(KEYINPUT52), .ZN(n682) );
  NOR2_X1 U739 ( .A1(n683), .A2(n682), .ZN(n686) );
  NOR2_X1 U740 ( .A1(n661), .A2(n684), .ZN(n685) );
  NOR2_X1 U741 ( .A1(n686), .A2(n685), .ZN(n694) );
  INV_X1 U742 ( .A(n687), .ZN(n720) );
  XNOR2_X1 U743 ( .A(KEYINPUT76), .B(KEYINPUT2), .ZN(n688) );
  NOR2_X1 U744 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U745 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U746 ( .A(KEYINPUT80), .B(n692), .Z(n693) );
  NAND2_X1 U747 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U748 ( .A1(n695), .A2(G953), .ZN(n696) );
  XNOR2_X1 U749 ( .A(n696), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U750 ( .A1(n712), .A2(G210), .ZN(n701) );
  XOR2_X1 U751 ( .A(KEYINPUT85), .B(KEYINPUT75), .Z(n698) );
  XNOR2_X1 U752 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n697) );
  XNOR2_X1 U753 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U754 ( .A(n702), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U755 ( .A1(n712), .A2(G469), .ZN(n707) );
  XNOR2_X1 U756 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n703), .B(KEYINPUT57), .ZN(n704) );
  XNOR2_X1 U758 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U759 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U760 ( .A1(n716), .A2(n708), .ZN(G54) );
  NAND2_X1 U761 ( .A1(n712), .A2(G478), .ZN(n709) );
  XOR2_X1 U762 ( .A(n710), .B(n709), .Z(n711) );
  NOR2_X1 U763 ( .A1(n716), .A2(n711), .ZN(G63) );
  NAND2_X1 U764 ( .A1(n712), .A2(G217), .ZN(n714) );
  XNOR2_X1 U765 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U766 ( .A1(n716), .A2(n715), .ZN(G66) );
  XNOR2_X1 U767 ( .A(n717), .B(KEYINPUT126), .ZN(n719) );
  NAND2_X1 U768 ( .A1(n719), .A2(n718), .ZN(n727) );
  NOR2_X1 U769 ( .A1(n720), .A2(G953), .ZN(n725) );
  NAND2_X1 U770 ( .A1(G953), .A2(G224), .ZN(n721) );
  XOR2_X1 U771 ( .A(KEYINPUT61), .B(n721), .Z(n722) );
  NOR2_X1 U772 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U773 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U774 ( .A(n727), .B(n726), .ZN(G69) );
  XNOR2_X1 U775 ( .A(n729), .B(n728), .ZN(n732) );
  NAND2_X1 U776 ( .A1(n731), .A2(n730), .ZN(n737) );
  XNOR2_X1 U777 ( .A(n732), .B(G227), .ZN(n733) );
  NAND2_X1 U778 ( .A1(n733), .A2(G900), .ZN(n734) );
  XOR2_X1 U779 ( .A(KEYINPUT127), .B(n734), .Z(n735) );
  NAND2_X1 U780 ( .A1(G953), .A2(n735), .ZN(n736) );
  NAND2_X1 U781 ( .A1(n737), .A2(n736), .ZN(G72) );
  XNOR2_X1 U782 ( .A(G125), .B(n738), .ZN(n739) );
  XNOR2_X1 U783 ( .A(n739), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U784 ( .A(G131), .B(n740), .Z(G33) );
  XNOR2_X1 U785 ( .A(G134), .B(n741), .ZN(G36) );
  XNOR2_X1 U786 ( .A(G143), .B(n742), .ZN(G45) );
  XOR2_X1 U787 ( .A(n743), .B(G137), .Z(G39) );
  BUF_X1 U788 ( .A(n744), .Z(n745) );
  XOR2_X1 U789 ( .A(G119), .B(n745), .Z(G21) );
endmodule

