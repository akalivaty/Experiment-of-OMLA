//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  OAI211_X1 g005(.A(new_n187), .B(KEYINPUT11), .C1(new_n188), .C2(G137), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT70), .B1(new_n193), .B2(G134), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT70), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(new_n188), .A3(G137), .ZN(new_n196));
  AOI22_X1  g010(.A1(new_n191), .A2(new_n192), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(new_n196), .ZN(new_n200));
  INV_X1    g014(.A(new_n192), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n193), .A2(G134), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT11), .B1(new_n202), .B2(new_n187), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n198), .B(new_n200), .C1(new_n201), .C2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT71), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n197), .A2(KEYINPUT71), .A3(new_n198), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n199), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT10), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT66), .A2(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT66), .A2(G146), .ZN(new_n211));
  OAI21_X1  g025(.A(G143), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT65), .A2(G143), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT65), .A2(G143), .ZN(new_n214));
  OAI21_X1  g028(.A(G146), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT65), .A2(G143), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n217), .B1(new_n223), .B2(KEYINPUT1), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT87), .B1(new_n216), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n212), .A2(new_n215), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT87), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n213), .A2(new_n214), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(new_n221), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n226), .B(new_n227), .C1(new_n230), .C2(new_n217), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n212), .A2(new_n215), .A3(new_n228), .A4(G128), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n225), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G104), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT3), .B1(new_n234), .B2(G107), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n236));
  INV_X1    g050(.A(G107), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(G104), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(G107), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n235), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G101), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n239), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n234), .A2(G107), .ZN(new_n244));
  OAI21_X1  g058(.A(G101), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n233), .A2(KEYINPUT88), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT88), .B1(new_n233), .B2(new_n246), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n209), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT86), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n240), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n235), .A2(new_n238), .A3(new_n239), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT86), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n253), .A3(G101), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT4), .A3(new_n242), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT0), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(new_n217), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n212), .A2(new_n215), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n212), .A2(new_n215), .A3(KEYINPUT67), .A4(new_n257), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OR2_X1    g076(.A1(KEYINPUT66), .A2(G146), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT66), .A2(G146), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n219), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n257), .B1(new_n265), .B2(new_n223), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n256), .A2(new_n217), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n251), .A2(new_n253), .A3(new_n269), .A4(G101), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n255), .A2(new_n262), .A3(new_n268), .A4(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT73), .B(G128), .Z(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(KEYINPUT1), .B2(new_n212), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n265), .A2(new_n223), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n232), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n246), .A2(new_n275), .A3(KEYINPUT10), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n208), .B1(new_n249), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n271), .A2(new_n276), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n233), .A2(new_n246), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT88), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n233), .A2(KEYINPUT88), .A3(new_n246), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n280), .B1(new_n285), .B2(new_n209), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT89), .B1(new_n286), .B2(new_n208), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n249), .A2(new_n277), .A3(KEYINPUT89), .A4(new_n208), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n279), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT91), .ZN(new_n291));
  OR2_X1    g105(.A1(KEYINPUT78), .A2(G953), .ZN(new_n292));
  NAND2_X1  g106(.A1(KEYINPUT78), .A2(G953), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G227), .ZN(new_n295));
  XNOR2_X1  g109(.A(G110), .B(G140), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n290), .A2(new_n291), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n249), .A2(new_n208), .A3(new_n277), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT89), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n278), .B1(new_n302), .B2(new_n288), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT91), .B1(new_n303), .B2(new_n297), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n246), .A2(new_n275), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n306), .B1(new_n283), .B2(new_n284), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(new_n208), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT12), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n302), .A2(new_n288), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(new_n297), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n299), .A2(new_n304), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G469), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n310), .A2(new_n297), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT90), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT90), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n310), .A2(new_n318), .A3(new_n297), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n279), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n297), .B1(new_n309), .B2(new_n310), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(G469), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(G469), .A2(G902), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n315), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT98), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT73), .B(G128), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(new_n219), .ZN(new_n328));
  OAI21_X1  g142(.A(G134), .B1(new_n328), .B2(KEYINPUT13), .ZN(new_n329));
  OAI22_X1  g143(.A1(new_n229), .A2(new_n217), .B1(new_n327), .B2(new_n219), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(KEYINPUT75), .A2(G116), .ZN(new_n332));
  NOR2_X1   g146(.A1(KEYINPUT75), .A2(G116), .ZN(new_n333));
  OAI21_X1  g147(.A(G122), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G116), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(G122), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(G107), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n330), .B(G134), .ZN(new_n339));
  OAI211_X1 g153(.A(KEYINPUT14), .B(G122), .C1(new_n332), .C2(new_n333), .ZN(new_n340));
  OAI211_X1 g154(.A(G107), .B(new_n340), .C1(new_n336), .C2(KEYINPUT14), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n339), .B(new_n341), .C1(G107), .C2(new_n336), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g157(.A(KEYINPUT9), .B(G234), .Z(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G217), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n345), .A2(new_n346), .A3(G953), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n338), .A2(new_n342), .A3(new_n347), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G478), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n352), .A2(KEYINPUT15), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n314), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n353), .B1(new_n351), .B2(new_n314), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G237), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n294), .A2(G214), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n229), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n294), .A2(new_n219), .A3(G214), .A4(new_n358), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n360), .A2(KEYINPUT17), .A3(G131), .A4(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT16), .ZN(new_n363));
  INV_X1    g177(.A(G140), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(G125), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n365), .A2(KEYINPUT82), .ZN(new_n366));
  XNOR2_X1  g180(.A(G125), .B(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT16), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(KEYINPUT82), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n221), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n366), .A2(new_n368), .A3(G146), .A4(new_n369), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n362), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT95), .ZN(new_n374));
  AOI21_X1  g188(.A(G131), .B1(new_n360), .B2(new_n361), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT17), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n360), .A2(G131), .A3(new_n361), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT95), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n362), .A2(new_n380), .A3(new_n371), .A4(new_n372), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n374), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n360), .A2(new_n361), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT18), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n360), .A2(KEYINPUT18), .A3(G131), .A4(new_n361), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n367), .B1(new_n211), .B2(new_n210), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n221), .B2(new_n367), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n376), .A2(new_n385), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(G113), .B(G122), .Z(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT94), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(new_n234), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n382), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n392), .B1(new_n382), .B2(new_n389), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n314), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G475), .ZN(new_n397));
  INV_X1    g211(.A(new_n378), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT19), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n367), .B(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n210), .A2(new_n211), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n372), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI22_X1  g216(.A1(new_n398), .A2(new_n375), .B1(new_n402), .B2(KEYINPUT93), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n402), .A2(KEYINPUT93), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n389), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n392), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(G475), .B1(new_n393), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n314), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n408), .B2(new_n314), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n357), .B(new_n397), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT21), .B(G898), .Z(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT96), .ZN(new_n415));
  AOI211_X1 g229(.A(new_n314), .B(new_n294), .C1(G234), .C2(G237), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G952), .ZN(new_n418));
  AOI211_X1 g232(.A(G953), .B(new_n418), .C1(G234), .C2(G237), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n420), .B(KEYINPUT97), .Z(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n326), .B1(new_n413), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n412), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n424), .A2(new_n410), .B1(G475), .B2(new_n396), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n425), .A2(KEYINPUT98), .A3(new_n421), .A4(new_n357), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G221), .B1(new_n345), .B2(G902), .ZN(new_n429));
  OAI21_X1  g243(.A(G214), .B1(G237), .B2(G902), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n262), .A2(new_n268), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G125), .ZN(new_n433));
  INV_X1    g247(.A(G125), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n275), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G224), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(G953), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n436), .B(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT2), .ZN(new_n441));
  INV_X1    g255(.A(G113), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT74), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT74), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(KEYINPUT2), .B2(G113), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G119), .B1(new_n332), .B2(new_n333), .ZN(new_n447));
  NAND2_X1  g261(.A1(KEYINPUT2), .A2(G113), .ZN(new_n448));
  INV_X1    g262(.A(G119), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G116), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n446), .A2(new_n447), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT5), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n449), .A3(G116), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT92), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n447), .A2(new_n450), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n454), .B(G113), .C1(new_n452), .C2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n246), .A2(new_n451), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n255), .A2(new_n270), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n446), .A2(new_n448), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n455), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n460), .A2(new_n451), .A3(KEYINPUT76), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT76), .B1(new_n460), .B2(new_n451), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n457), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n465));
  XOR2_X1   g279(.A(G110), .B(G122), .Z(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n466), .ZN(new_n468));
  INV_X1    g282(.A(new_n466), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n457), .B(new_n469), .C1(new_n458), .C2(new_n463), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(KEYINPUT6), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n440), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n456), .A2(new_n451), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n473), .B(new_n246), .Z(new_n474));
  XOR2_X1   g288(.A(new_n466), .B(KEYINPUT8), .Z(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n436), .A2(KEYINPUT7), .A3(new_n439), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n439), .A2(KEYINPUT7), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n433), .A2(new_n435), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n476), .A2(new_n477), .A3(new_n479), .A4(new_n470), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n472), .A2(new_n314), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G210), .B1(G237), .B2(G902), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n472), .A2(new_n314), .A3(new_n482), .A4(new_n480), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n431), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n325), .A2(new_n428), .A3(new_n429), .A4(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT28), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n193), .A2(G134), .ZN(new_n489));
  INV_X1    g303(.A(new_n202), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n490), .B2(KEYINPUT72), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(KEYINPUT72), .B2(new_n490), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G131), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n204), .A2(new_n205), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT71), .B1(new_n197), .B2(new_n198), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n275), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT77), .ZN(new_n497));
  OAI22_X1  g311(.A1(new_n494), .A2(new_n495), .B1(new_n198), .B2(new_n197), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n432), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n206), .A2(new_n207), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT77), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n275), .A4(new_n493), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n463), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n497), .A2(new_n499), .A3(new_n463), .A4(new_n502), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n488), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n262), .A2(new_n268), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n496), .B(new_n463), .C1(new_n208), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n488), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT79), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(KEYINPUT79), .A3(new_n488), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT29), .B1(new_n507), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n506), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT68), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n262), .A2(KEYINPUT68), .A3(new_n268), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n498), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n463), .B1(new_n520), .B2(new_n496), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT28), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT29), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n522), .A2(new_n523), .A3(new_n512), .A4(new_n513), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(G101), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n294), .A2(G210), .A3(new_n358), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n515), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT30), .A4(new_n502), .ZN(new_n530));
  INV_X1    g344(.A(new_n496), .ZN(new_n531));
  AOI221_X4 g345(.A(new_n517), .B1(new_n266), .B2(new_n267), .C1(new_n260), .C2(new_n261), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT68), .B1(new_n262), .B2(new_n268), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n531), .B1(new_n534), .B2(new_n498), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n504), .B(new_n530), .C1(new_n535), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n528), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n506), .A3(new_n539), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n540), .A2(KEYINPUT29), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n529), .A2(new_n314), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G472), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT81), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n506), .A3(new_n528), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT31), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n520), .A2(new_n496), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n504), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n488), .B1(new_n549), .B2(new_n506), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n539), .B1(new_n550), .B2(new_n514), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT31), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n538), .A2(new_n552), .A3(new_n506), .A4(new_n528), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n547), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G472), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n314), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT80), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT32), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT32), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n554), .A2(new_n560), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n542), .A2(KEYINPUT81), .A3(G472), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n545), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n294), .A2(G221), .A3(G234), .ZN(new_n565));
  XOR2_X1   g379(.A(new_n565), .B(KEYINPUT22), .Z(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G137), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n449), .A2(G128), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(new_n327), .B2(new_n449), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT24), .B(G110), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(KEYINPUT23), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT23), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n449), .B2(G128), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n571), .B1(new_n575), .B2(G110), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n372), .A3(new_n387), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT84), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(G110), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n371), .A2(new_n372), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n580), .B(new_n581), .C1(new_n569), .C2(new_n570), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT83), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n567), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n577), .B(KEYINPUT84), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT83), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n582), .B(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n567), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT25), .B1(new_n590), .B2(G902), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n346), .B1(G234), .B2(new_n314), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT25), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n584), .A2(new_n589), .A3(new_n593), .A4(new_n314), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT85), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n592), .A2(G902), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n584), .A2(KEYINPUT85), .A3(new_n589), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n564), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n487), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(new_n241), .ZN(G3));
  NAND3_X1  g418(.A1(new_n325), .A2(new_n601), .A3(new_n429), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n554), .A2(new_n314), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G472), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n607), .A2(KEYINPUT99), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(KEYINPUT99), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n558), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n611), .B(KEYINPUT100), .Z(new_n612));
  NAND2_X1  g426(.A1(new_n486), .A2(new_n421), .ZN(new_n613));
  INV_X1    g427(.A(new_n425), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n351), .B(KEYINPUT33), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n615), .A2(KEYINPUT101), .A3(G478), .A4(new_n314), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n351), .A2(KEYINPUT33), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n349), .B2(new_n350), .ZN(new_n619));
  OAI211_X1 g433(.A(G478), .B(new_n314), .C1(new_n617), .C2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n351), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n352), .B1(new_n623), .B2(G902), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n616), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n614), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n613), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n612), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT34), .B(G104), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT102), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n628), .B(new_n630), .ZN(G6));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n410), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n411), .A2(new_n412), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n633), .B1(new_n634), .B2(new_n632), .ZN(new_n635));
  INV_X1    g449(.A(new_n357), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n397), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n613), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n612), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n567), .A2(KEYINPUT36), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT104), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n585), .A2(new_n587), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n598), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n595), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n608), .A2(new_n558), .A3(new_n609), .A4(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n487), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT37), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G110), .ZN(G12));
  INV_X1    g466(.A(G900), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n419), .B1(new_n416), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n396), .B2(G475), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n635), .A2(KEYINPUT105), .A3(new_n636), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n424), .A2(new_n632), .A3(new_n410), .ZN(new_n657));
  INV_X1    g471(.A(new_n633), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n657), .A2(new_n658), .A3(new_n636), .A4(new_n655), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n325), .A2(new_n662), .A3(new_n429), .ZN(new_n663));
  INV_X1    g477(.A(new_n648), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n542), .A2(KEYINPUT81), .A3(G472), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT81), .B1(new_n542), .B2(G472), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n664), .B1(new_n667), .B2(new_n562), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n663), .A2(new_n668), .A3(KEYINPUT106), .A4(new_n486), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n564), .A2(new_n486), .A3(new_n648), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n325), .A2(new_n662), .A3(new_n429), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  XNOR2_X1  g489(.A(new_n654), .B(KEYINPUT39), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n325), .A2(new_n429), .A3(new_n677), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n425), .A2(new_n357), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n678), .B2(KEYINPUT40), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n484), .A2(new_n485), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT38), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n538), .A2(new_n506), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n528), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n505), .A2(new_n506), .A3(new_n539), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n314), .A3(new_n687), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n559), .A2(new_n561), .B1(G472), .B2(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n689), .A2(new_n431), .A3(new_n648), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n679), .A2(new_n682), .A3(new_n684), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n229), .ZN(G45));
  INV_X1    g506(.A(new_n671), .ZN(new_n693));
  INV_X1    g507(.A(new_n626), .ZN(new_n694));
  INV_X1    g508(.A(new_n654), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n325), .A2(new_n429), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  INV_X1    g513(.A(new_n602), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n313), .B1(new_n312), .B2(new_n314), .ZN(new_n702));
  INV_X1    g516(.A(new_n429), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n700), .A2(new_n627), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT107), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT41), .B(G113), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NAND4_X1  g522(.A1(new_n704), .A2(new_n601), .A3(new_n564), .A4(new_n639), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  NAND4_X1  g524(.A1(new_n668), .A2(new_n486), .A3(new_n428), .A4(new_n704), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  OAI21_X1  g526(.A(new_n539), .B1(new_n507), .B2(new_n514), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n547), .A2(new_n713), .A3(new_n553), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n557), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n714), .A2(KEYINPUT108), .A3(new_n557), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n601), .A2(new_n607), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n613), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n704), .A3(new_n680), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NAND2_X1  g536(.A1(new_n312), .A2(new_n314), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G469), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(new_n429), .A3(new_n315), .A4(new_n486), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n626), .A2(new_n654), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n717), .A2(new_n718), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n607), .A3(new_n648), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  NAND3_X1  g547(.A1(new_n484), .A2(new_n430), .A3(new_n485), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n734), .B(KEYINPUT109), .Z(new_n735));
  AND3_X1   g549(.A1(new_n564), .A2(new_n735), .A3(new_n601), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT42), .B1(new_n736), .B2(new_n697), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n564), .A2(new_n735), .A3(new_n601), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n738), .A2(new_n696), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n198), .ZN(G33));
  NOR2_X1   g556(.A1(new_n738), .A2(new_n672), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n188), .ZN(G36));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n318), .B1(new_n310), .B2(new_n297), .ZN(new_n746));
  AOI211_X1 g560(.A(KEYINPUT90), .B(new_n298), .C1(new_n302), .C2(new_n288), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n746), .A2(new_n747), .A3(new_n278), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n745), .B1(new_n748), .B2(new_n321), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n320), .A2(KEYINPUT45), .A3(new_n322), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(G469), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT46), .B1(new_n751), .B2(new_n324), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI211_X1 g568(.A(KEYINPUT110), .B(KEYINPUT46), .C1(new_n751), .C2(new_n324), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n751), .A2(KEYINPUT46), .A3(new_n324), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n315), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n703), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(KEYINPUT111), .ZN(new_n761));
  INV_X1    g575(.A(new_n625), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n761), .B1(new_n762), .B2(new_n614), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n614), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n760), .A2(KEYINPUT111), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n763), .B1(new_n766), .B2(new_n761), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n610), .A3(new_n648), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n769), .A2(KEYINPUT44), .ZN(new_n770));
  INV_X1    g584(.A(new_n735), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n769), .B2(KEYINPUT44), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n759), .A2(new_n770), .A3(new_n677), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT112), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n193), .ZN(G39));
  OR3_X1    g589(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n776));
  XNOR2_X1  g590(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n429), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n777), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(new_n758), .B2(new_n703), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n771), .A2(new_n564), .A3(new_n727), .A4(new_n601), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n701), .A2(new_n702), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n429), .A3(new_n486), .A4(new_n726), .ZN(new_n786));
  OAI22_X1  g600(.A1(new_n786), .A2(new_n730), .B1(new_n671), .B2(new_n696), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n673), .B2(new_n669), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n325), .A2(new_n429), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n689), .A2(new_n648), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n680), .A2(new_n486), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n790), .A2(new_n695), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT52), .B1(new_n788), .B2(new_n793), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n693), .A2(new_n697), .B1(new_n728), .B2(new_n731), .ZN(new_n795));
  AND4_X1   g609(.A1(KEYINPUT52), .A2(new_n674), .A3(new_n795), .A4(new_n793), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n709), .A2(new_n721), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(KEYINPUT114), .A3(new_n705), .A4(new_n711), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n704), .A2(new_n601), .A3(new_n564), .ZN(new_n801));
  INV_X1    g615(.A(new_n627), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n704), .A2(new_n428), .ZN(new_n803));
  OAI22_X1  g617(.A1(new_n801), .A2(new_n802), .B1(new_n803), .B2(new_n671), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n709), .A2(new_n721), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n800), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n799), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n726), .A2(new_n729), .A3(new_n607), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n545), .A2(new_n562), .A3(new_n563), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n635), .A2(new_n357), .A3(new_n655), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n635), .A2(KEYINPUT116), .A3(new_n357), .A4(new_n655), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n808), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n790), .A3(new_n648), .A4(new_n735), .ZN(new_n816));
  INV_X1    g630(.A(new_n743), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n816), .B(new_n817), .C1(new_n737), .C2(new_n740), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n626), .B1(new_n357), .B2(new_n614), .ZN(new_n820));
  INV_X1    g634(.A(new_n613), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n605), .A2(new_n610), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n487), .ZN(new_n825));
  INV_X1    g639(.A(new_n649), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n825), .B1(new_n700), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n827), .A3(KEYINPUT115), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n487), .B1(new_n602), .B2(new_n649), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n829), .B1(new_n830), .B2(new_n823), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n807), .A2(new_n819), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n784), .B1(new_n797), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n807), .A2(new_n832), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n788), .A2(KEYINPUT52), .A3(new_n793), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n674), .A2(new_n795), .A3(new_n793), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n835), .A2(KEYINPUT53), .A3(new_n840), .A4(new_n819), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n834), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n816), .A2(KEYINPUT53), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n741), .A2(new_n743), .A3(new_n805), .A4(new_n804), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n840), .A2(new_n832), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n834), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n767), .A2(new_n419), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n719), .ZN(new_n850));
  INV_X1    g664(.A(new_n684), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n704), .A2(new_n431), .A3(new_n851), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n852), .A2(KEYINPUT117), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(KEYINPUT117), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT50), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n704), .A2(new_n735), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n849), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n689), .A2(new_n419), .ZN(new_n863));
  INV_X1    g677(.A(new_n601), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n614), .A2(new_n625), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n862), .A2(new_n731), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n857), .A2(new_n868), .A3(new_n858), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n860), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n778), .A2(new_n780), .B1(new_n703), .B2(new_n785), .ZN(new_n871));
  INV_X1    g685(.A(new_n850), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n871), .A2(new_n771), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n843), .B(new_n848), .C1(KEYINPUT51), .C2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n873), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(KEYINPUT51), .A3(new_n859), .A4(new_n867), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n862), .A2(new_n700), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT48), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n418), .A2(G953), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n872), .B2(new_n725), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n694), .B2(new_n865), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n877), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  OAI22_X1  g697(.A1(new_n875), .A2(new_n883), .B1(G952), .B2(G953), .ZN(new_n884));
  INV_X1    g698(.A(new_n785), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n430), .B(new_n764), .C1(new_n885), .C2(KEYINPUT49), .ZN(new_n886));
  AOI211_X1 g700(.A(new_n864), .B(new_n886), .C1(KEYINPUT49), .C2(new_n885), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n429), .A3(new_n851), .A4(new_n689), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n884), .A2(new_n888), .ZN(G75));
  NOR2_X1   g703(.A1(new_n294), .A2(G952), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT119), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n834), .A2(new_n847), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(G210), .A3(G902), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n471), .A2(new_n467), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n440), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT55), .Z(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n898), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n893), .A2(new_n894), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n891), .B1(new_n899), .B2(new_n901), .ZN(G51));
  XOR2_X1   g716(.A(new_n324), .B(KEYINPUT57), .Z(new_n903));
  AND3_X1   g717(.A1(new_n834), .A2(new_n844), .A3(new_n847), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n844), .B1(new_n834), .B2(new_n847), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n312), .B(KEYINPUT120), .Z(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n892), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n909), .A2(new_n314), .A3(new_n751), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n890), .B1(new_n908), .B2(new_n910), .ZN(G54));
  NAND3_X1  g725(.A1(new_n892), .A2(KEYINPUT58), .A3(G902), .ZN(new_n912));
  INV_X1    g726(.A(G475), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n393), .A2(new_n407), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n890), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n912), .B2(new_n913), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G60));
  INV_X1    g733(.A(new_n615), .ZN(new_n920));
  NAND2_X1  g734(.A1(G478), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT59), .Z(new_n922));
  NOR2_X1   g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n904), .B2(new_n905), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT121), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n926), .B(new_n923), .C1(new_n904), .C2(new_n905), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n891), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n922), .B1(new_n843), .B2(new_n848), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(new_n615), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n928), .A2(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(new_n597), .A2(new_n599), .ZN(new_n933));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT122), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT60), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n933), .B1(new_n909), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n892), .A2(new_n646), .A3(new_n936), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n938), .A2(new_n929), .A3(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n938), .A2(KEYINPUT61), .A3(new_n929), .A4(new_n939), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(G66));
  OAI21_X1  g758(.A(G953), .B1(new_n415), .B2(new_n437), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n807), .B2(new_n832), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n807), .A2(new_n946), .A3(new_n832), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n294), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(G898), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n896), .B1(new_n953), .B2(new_n951), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n952), .B(new_n954), .Z(G69));
  NAND3_X1  g769(.A1(new_n691), .A2(new_n674), .A3(new_n795), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n788), .A2(KEYINPUT62), .A3(new_n691), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n736), .A2(new_n790), .A3(new_n677), .A4(new_n820), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n960), .A2(new_n782), .A3(new_n773), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n294), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n530), .B1(new_n535), .B2(new_n537), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(new_n400), .Z(new_n965));
  AOI21_X1  g779(.A(KEYINPUT124), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n967));
  INV_X1    g781(.A(new_n965), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n967), .B(new_n968), .C1(new_n962), .C2(new_n294), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n294), .B1(G227), .B2(G900), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n674), .A2(new_n795), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n817), .B1(new_n737), .B2(new_n740), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n759), .A2(new_n700), .A3(new_n677), .A4(new_n792), .ZN(new_n975));
  AND4_X1   g789(.A1(new_n773), .A2(new_n782), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n965), .B1(new_n976), .B2(new_n294), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n653), .B2(new_n294), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n970), .A2(new_n971), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n971), .B1(new_n970), .B2(new_n978), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(G72));
  XNOR2_X1  g795(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n555), .A2(new_n314), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n982), .B(new_n983), .Z(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n976), .B2(new_n950), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n917), .B1(new_n986), .B2(new_n540), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g803(.A(KEYINPUT127), .B(new_n917), .C1(new_n986), .C2(new_n540), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n842), .A2(new_n540), .A3(new_n686), .A4(new_n984), .ZN(new_n992));
  INV_X1    g806(.A(new_n949), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n993), .A2(new_n947), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n984), .B1(new_n994), .B2(new_n962), .ZN(new_n995));
  INV_X1    g809(.A(new_n686), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n995), .A2(KEYINPUT126), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(KEYINPUT126), .B1(new_n995), .B2(new_n996), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n992), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n991), .A2(new_n999), .ZN(G57));
endmodule


