//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G125), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n188), .A2(KEYINPUT16), .A3(G140), .ZN(new_n189));
  XNOR2_X1  g003(.A(G125), .B(G140), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(KEYINPUT16), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n191), .A2(G146), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT92), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n194), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT92), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(new_n192), .ZN(new_n198));
  INV_X1    g012(.A(G237), .ZN(new_n199));
  INV_X1    g013(.A(G953), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G214), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  XNOR2_X1  g016(.A(new_n201), .B(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n201), .B(G143), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n203), .A2(KEYINPUT17), .A3(G131), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n195), .A2(new_n198), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G113), .B(G122), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT18), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n205), .B1(new_n215), .B2(new_n206), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n203), .A2(KEYINPUT18), .A3(G131), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n190), .B(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n211), .A2(new_n214), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n214), .B1(new_n211), .B2(new_n220), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n187), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G475), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT20), .ZN(new_n225));
  NOR2_X1   g039(.A1(G475), .A2(G902), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT89), .ZN(new_n227));
  INV_X1    g041(.A(G140), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G125), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n188), .A2(G140), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT90), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n227), .B(KEYINPUT19), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT89), .B1(new_n190), .B2(KEYINPUT90), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT19), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(new_n190), .B2(KEYINPUT89), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n233), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n192), .B1(new_n237), .B2(G146), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT91), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n204), .A2(new_n207), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n241), .B(new_n192), .C1(new_n237), .C2(G146), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n214), .B1(new_n243), .B2(new_n220), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n225), .B(new_n226), .C1(new_n244), .C2(new_n221), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n211), .A2(new_n214), .A3(new_n220), .ZN(new_n247));
  INV_X1    g061(.A(new_n220), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n238), .A2(KEYINPUT91), .B1(new_n204), .B2(new_n207), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(new_n242), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n247), .B1(new_n250), .B2(new_n214), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n225), .B1(new_n251), .B2(new_n226), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n224), .B1(new_n246), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT15), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G478), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT9), .B(G234), .ZN(new_n256));
  INV_X1    g070(.A(G217), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n256), .A2(new_n257), .A3(G953), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT96), .ZN(new_n259));
  OR2_X1    g073(.A1(KEYINPUT76), .A2(G107), .ZN(new_n260));
  INV_X1    g074(.A(G116), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G122), .ZN(new_n262));
  INV_X1    g076(.A(G122), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G116), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT76), .A2(G107), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n260), .A2(new_n262), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n202), .A2(G128), .ZN(new_n267));
  INV_X1    g081(.A(G128), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G143), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n267), .B2(new_n269), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n266), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n261), .A2(KEYINPUT14), .A3(G122), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G107), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n262), .A2(new_n264), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT14), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT95), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n268), .A2(G143), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n202), .A2(G128), .ZN(new_n281));
  OAI21_X1  g095(.A(G134), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n262), .A2(new_n264), .ZN(new_n285));
  OAI211_X1 g099(.A(G107), .B(new_n274), .C1(new_n285), .C2(KEYINPUT14), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT95), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n284), .A2(new_n286), .A3(new_n287), .A4(new_n266), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n279), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT76), .B(G107), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n262), .A2(new_n264), .B1(new_n260), .B2(new_n265), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n283), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT13), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n268), .B2(G143), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT93), .B1(new_n295), .B2(new_n280), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT93), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n297), .B(new_n267), .C1(new_n281), .C2(new_n294), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT94), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n280), .A2(new_n299), .A3(KEYINPUT13), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT94), .B1(new_n267), .B2(new_n294), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n296), .A2(new_n298), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n293), .B1(G134), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n259), .B1(new_n289), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(G134), .ZN(new_n305));
  INV_X1    g119(.A(new_n292), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n271), .B1(new_n306), .B2(new_n266), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n308), .A2(KEYINPUT96), .A3(new_n279), .A4(new_n288), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n258), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n258), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n279), .A3(new_n288), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(new_n259), .ZN(new_n313));
  OAI211_X1 g127(.A(KEYINPUT98), .B(new_n187), .C1(new_n310), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT97), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g130(.A(KEYINPUT97), .B(new_n187), .C1(new_n310), .C2(new_n313), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n255), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G952), .ZN(new_n319));
  AOI211_X1 g133(.A(G953), .B(new_n319), .C1(G234), .C2(G237), .ZN(new_n320));
  AOI211_X1 g134(.A(new_n187), .B(new_n200), .C1(G234), .C2(G237), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT21), .B(G898), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n314), .A2(new_n315), .B1(new_n254), .B2(G478), .ZN(new_n324));
  NOR4_X1   g138(.A1(new_n253), .A2(new_n318), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G221), .ZN(new_n326));
  INV_X1    g140(.A(new_n256), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(new_n187), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G110), .B(G140), .ZN(new_n330));
  INV_X1    g144(.A(G227), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G953), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT12), .ZN(new_n335));
  INV_X1    g149(.A(G107), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G104), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n213), .A2(KEYINPUT75), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n336), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g154(.A1(KEYINPUT76), .A2(G107), .ZN(new_n341));
  NOR2_X1   g155(.A1(KEYINPUT76), .A2(G107), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n213), .A2(KEYINPUT3), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n340), .A2(KEYINPUT3), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n213), .A2(KEYINPUT75), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n337), .A2(G104), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(G107), .ZN(new_n348));
  INV_X1    g162(.A(G101), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n213), .B1(new_n341), .B2(new_n342), .ZN(new_n354));
  AOI211_X1 g168(.A(new_n353), .B(new_n349), .C1(new_n340), .C2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT75), .B(G104), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n354), .B1(new_n356), .B2(G107), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT77), .B1(new_n357), .B2(G101), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n352), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n218), .A2(G143), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n202), .A2(G146), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT1), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .A4(G128), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n202), .A2(G146), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT64), .B1(new_n218), .B2(G143), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT64), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n202), .A3(G146), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n364), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n268), .B1(new_n360), .B2(KEYINPUT1), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(G104), .B1(new_n260), .B2(new_n265), .ZN(new_n372));
  AOI21_X1  g186(.A(G107), .B1(new_n346), .B2(new_n347), .ZN(new_n373));
  OAI21_X1  g187(.A(G101), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n353), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n357), .A2(KEYINPUT77), .A3(G101), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G143), .B(G146), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(G128), .B1(new_n364), .B2(new_n362), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n345), .A2(new_n351), .B1(new_n363), .B2(new_n381), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n359), .A2(new_n371), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT11), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n270), .B2(G137), .ZN(new_n385));
  INV_X1    g199(.A(G137), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT11), .A3(G134), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n270), .A2(G137), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G131), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n385), .A2(new_n387), .A3(new_n206), .A4(new_n388), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n335), .B1(new_n383), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n377), .A2(new_n382), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n375), .A2(new_n376), .B1(new_n345), .B2(new_n351), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n395), .B1(new_n396), .B2(new_n370), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(KEYINPUT12), .A3(new_n392), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT0), .A4(G128), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT65), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n378), .A2(KEYINPUT65), .A3(KEYINPUT0), .A4(G128), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n366), .B1(new_n202), .B2(G146), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n218), .A2(KEYINPUT64), .A3(G143), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n360), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(KEYINPUT0), .B(G128), .Z(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n345), .B2(new_n351), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n344), .A2(new_n260), .A3(new_n265), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n413), .B(new_n348), .C1(new_n373), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G101), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n410), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(new_n411), .A3(G101), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n370), .A2(KEYINPUT10), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n417), .A2(new_n418), .B1(new_n396), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT78), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT10), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n421), .B1(new_n395), .B2(new_n422), .ZN(new_n423));
  AOI211_X1 g237(.A(KEYINPUT78), .B(KEYINPUT10), .C1(new_n377), .C2(new_n382), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n420), .B(new_n393), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n334), .B1(new_n399), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n392), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n402), .A2(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n415), .A2(G101), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n413), .B1(new_n373), .B2(new_n414), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT4), .B1(new_n432), .B2(new_n350), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n430), .B(new_n418), .C1(new_n431), .C2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n377), .A2(new_n352), .A3(new_n419), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n363), .B1(new_n369), .B2(new_n378), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n432), .B2(new_n350), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n375), .B2(new_n376), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT78), .B1(new_n439), .B2(KEYINPUT10), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n395), .A2(new_n421), .A3(new_n422), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n436), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n333), .B1(new_n442), .B2(new_n393), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n429), .B1(new_n443), .B2(KEYINPUT79), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n425), .A2(new_n334), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT79), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n427), .B(G469), .C1(new_n444), .C2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G469), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n334), .B1(new_n429), .B2(new_n425), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n399), .A2(new_n425), .A3(new_n334), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n449), .B(new_n187), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n449), .A2(new_n187), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n448), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n325), .A2(new_n329), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT70), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n268), .B2(G119), .ZN(new_n458));
  INV_X1    g272(.A(G119), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT70), .A3(G128), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n268), .A2(G119), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT24), .B(G110), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT23), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n459), .A2(G128), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n268), .A2(KEYINPUT23), .A3(G119), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G110), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n192), .B2(new_n196), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n462), .A2(new_n463), .ZN(new_n474));
  INV_X1    g288(.A(G110), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n466), .A2(new_n468), .A3(new_n475), .A4(new_n467), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT71), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT71), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n474), .A2(new_n479), .A3(new_n476), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n231), .A2(G146), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n191), .B2(G146), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT72), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n474), .A2(new_n479), .A3(new_n476), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n479), .B1(new_n474), .B2(new_n476), .ZN(new_n486));
  OAI211_X1 g300(.A(KEYINPUT72), .B(new_n483), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n473), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT22), .B(G137), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n200), .A2(G221), .A3(G234), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT72), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n487), .ZN(new_n497));
  INV_X1    g311(.A(new_n492), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n473), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n187), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n493), .A2(KEYINPUT25), .A3(new_n187), .A4(new_n499), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n502), .A2(KEYINPUT73), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n257), .B1(G234), .B2(new_n187), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n502), .B2(KEYINPUT73), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n498), .B1(new_n497), .B2(new_n473), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n472), .B(new_n492), .C1(new_n496), .C2(new_n487), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT74), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT74), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n507), .B2(new_n508), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n505), .A2(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI22_X1  g329(.A1(new_n504), .A2(new_n506), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n392), .A2(new_n404), .A3(new_n409), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT67), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n430), .A2(KEYINPUT67), .A3(new_n392), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n270), .A2(G137), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n386), .A2(G134), .ZN(new_n523));
  OAI21_X1  g337(.A(G131), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n391), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n525), .A2(new_n370), .A3(KEYINPUT68), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT68), .B1(new_n525), .B2(new_n370), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n521), .A2(KEYINPUT30), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n459), .A2(G116), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n261), .A2(G119), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT2), .B(G113), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n532), .A2(new_n534), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n525), .A2(new_n370), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT66), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT66), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n525), .A2(new_n370), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n517), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n529), .A2(new_n538), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n538), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n521), .A2(new_n547), .A3(new_n528), .ZN(new_n548));
  XOR2_X1   g362(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n549));
  NAND3_X1  g363(.A1(new_n199), .A2(new_n200), .A3(G210), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT26), .B(G101), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n546), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n546), .A2(KEYINPUT31), .A3(new_n548), .A4(new_n553), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n538), .B1(new_n370), .B2(new_n525), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT28), .B1(new_n559), .B2(new_n517), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n543), .A2(new_n538), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n548), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT28), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n553), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n558), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT32), .ZN(new_n569));
  NOR2_X1   g383(.A1(G472), .A2(G902), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n556), .A2(new_n557), .B1(new_n565), .B2(new_n566), .ZN(new_n572));
  INV_X1    g386(.A(new_n570), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT32), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n546), .A2(new_n548), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n566), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT29), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n577), .B(new_n578), .C1(new_n565), .C2(new_n566), .ZN(new_n579));
  AND4_X1   g393(.A1(KEYINPUT67), .A2(new_n392), .A3(new_n404), .A4(new_n409), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT67), .B1(new_n430), .B2(new_n392), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n527), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n525), .A2(new_n370), .A3(KEYINPUT68), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n538), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n564), .B1(new_n586), .B2(new_n548), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(new_n560), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n566), .A2(new_n578), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n579), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n516), .B1(new_n575), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(G214), .B1(G237), .B2(G902), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n538), .B(new_n418), .C1(new_n431), .C2(new_n433), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n533), .A2(KEYINPUT5), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n530), .A2(KEYINPUT5), .ZN(new_n598));
  INV_X1    g412(.A(G113), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n597), .A2(new_n600), .B1(new_n533), .B2(new_n535), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n352), .B(new_n601), .C1(new_n355), .C2(new_n358), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT80), .B1(new_n596), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n596), .A2(KEYINPUT80), .A3(new_n602), .ZN(new_n605));
  XNOR2_X1  g419(.A(G110), .B(G122), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n606), .B(KEYINPUT81), .Z(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n604), .A2(KEYINPUT6), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT6), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n596), .A2(new_n602), .A3(new_n607), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT82), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n596), .A2(KEYINPUT82), .A3(new_n602), .A4(new_n607), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n596), .A2(KEYINPUT80), .A3(new_n602), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n616), .A2(new_n603), .A3(new_n607), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n609), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n410), .A2(G125), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT83), .ZN(new_n620));
  OR3_X1    g434(.A1(new_n430), .A2(KEYINPUT83), .A3(new_n188), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n371), .A2(new_n188), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT84), .B(G224), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(G953), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT85), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT86), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n623), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n618), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n619), .A2(new_n622), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT7), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n630), .B1(new_n631), .B2(new_n626), .ZN(new_n632));
  INV_X1    g446(.A(new_n601), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n359), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n634), .A2(new_n602), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n607), .B(KEYINPUT8), .Z(new_n636));
  OAI21_X1  g450(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT87), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n631), .B1(new_n626), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n638), .B2(new_n626), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n623), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n613), .A2(new_n614), .ZN(new_n643));
  AOI21_X1  g457(.A(G902), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n629), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(G210), .B1(G237), .B2(G902), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT88), .Z(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n629), .A2(new_n644), .A3(new_n646), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n595), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n456), .A2(new_n593), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G101), .ZN(G3));
  AOI21_X1  g466(.A(new_n646), .B1(new_n629), .B2(new_n644), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n595), .B1(new_n654), .B2(new_n649), .ZN(new_n655));
  INV_X1    g469(.A(new_n323), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n312), .A2(new_n657), .A3(new_n258), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n258), .B1(new_n312), .B2(new_n657), .ZN(new_n660));
  OAI21_X1  g474(.A(KEYINPUT33), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT33), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(new_n310), .B2(new_n313), .ZN(new_n663));
  INV_X1    g477(.A(G478), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(G902), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n661), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n187), .B1(new_n310), .B2(new_n313), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n667), .A2(KEYINPUT100), .A3(new_n664), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT100), .B1(new_n667), .B2(new_n664), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n253), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n655), .A2(new_n656), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n452), .A2(new_n454), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n440), .A2(new_n441), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n393), .B1(new_n676), .B2(new_n420), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n445), .B2(new_n446), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n443), .A2(KEYINPUT79), .ZN(new_n679));
  AOI211_X1 g493(.A(new_n449), .B(new_n426), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n329), .B1(new_n675), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n572), .B2(G902), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n572), .B2(new_n573), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n681), .A2(new_n683), .A3(new_n516), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n674), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT34), .B(G104), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G6));
  INV_X1    g501(.A(new_n318), .ZN(new_n688));
  INV_X1    g502(.A(new_n324), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n253), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n655), .A2(new_n656), .A3(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n684), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT101), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT35), .B(G107), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G9));
  NOR2_X1   g510(.A1(new_n492), .A2(KEYINPUT36), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n489), .A2(KEYINPUT102), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n497), .B2(new_n473), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n698), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n699), .A2(new_n701), .A3(new_n698), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n514), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n504), .B2(new_n506), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT103), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n708), .B(new_n705), .C1(new_n504), .C2(new_n506), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n683), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n456), .A2(new_n710), .A3(new_n650), .A4(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT37), .B(G110), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G12));
  INV_X1    g528(.A(G900), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n320), .B1(new_n321), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n690), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n707), .B2(new_n709), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n569), .B1(new_n568), .B2(new_n570), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n572), .A2(KEYINPUT32), .A3(new_n573), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n592), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n629), .A2(new_n646), .A3(new_n644), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n594), .B1(new_n723), .B2(new_n653), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n681), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n719), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G128), .ZN(G30));
  AND3_X1   g541(.A1(new_n521), .A2(new_n547), .A3(new_n528), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n547), .B1(new_n521), .B2(new_n528), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n566), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n554), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n731), .B2(G902), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n575), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT40), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT105), .B(KEYINPUT39), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n716), .B(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n455), .A2(new_n329), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n733), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(new_n734), .B2(new_n737), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n648), .A2(new_n649), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n710), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n253), .B1(new_n318), .B2(new_n324), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n594), .A3(new_n743), .A4(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n739), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n202), .ZN(G45));
  NAND3_X1  g562(.A1(new_n670), .A2(new_n253), .A3(new_n717), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n725), .A2(new_n722), .A3(new_n710), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G146), .ZN(G48));
  AOI21_X1  g566(.A(new_n515), .B1(new_n510), .B2(new_n512), .ZN(new_n753));
  INV_X1    g567(.A(new_n505), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT25), .B1(new_n509), .B2(new_n187), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT73), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n502), .A2(KEYINPUT73), .A3(new_n503), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n753), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n187), .B1(new_n450), .B2(new_n451), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(G469), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n761), .A2(new_n329), .A3(new_n452), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n722), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n673), .ZN(new_n764));
  XOR2_X1   g578(.A(KEYINPUT41), .B(G113), .Z(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G15));
  NOR2_X1   g580(.A1(new_n763), .A2(new_n691), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n261), .ZN(G18));
  NAND2_X1  g582(.A1(new_n710), .A2(new_n722), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n655), .A2(new_n325), .A3(new_n762), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n459), .ZN(G21));
  NAND2_X1  g586(.A1(new_n568), .A2(new_n187), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT106), .B1(new_n587), .B2(new_n560), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT28), .B1(new_n728), .B2(new_n729), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT106), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n561), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(new_n777), .A3(new_n566), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n558), .ZN(new_n779));
  AOI22_X1  g593(.A1(new_n773), .A2(G472), .B1(new_n570), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n762), .A2(new_n780), .A3(new_n759), .A4(new_n656), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n655), .A2(new_n745), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n263), .ZN(G24));
  NAND2_X1  g598(.A1(new_n779), .A2(new_n570), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n682), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n707), .B2(new_n709), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n761), .A2(new_n329), .A3(new_n452), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n724), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n749), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n670), .A2(new_n253), .A3(KEYINPUT107), .A4(new_n717), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n787), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G125), .ZN(G27));
  AND3_X1   g609(.A1(new_n722), .A2(KEYINPUT110), .A3(new_n759), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT110), .B1(new_n722), .B2(new_n759), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n647), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n629), .B2(new_n644), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n723), .A2(new_n800), .A3(new_n595), .ZN(new_n801));
  INV_X1    g615(.A(new_n425), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n333), .B1(new_n802), .B2(new_n677), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n399), .A2(new_n425), .A3(new_n334), .ZN(new_n804));
  AOI21_X1  g618(.A(G902), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n453), .B1(new_n805), .B2(new_n449), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n328), .B1(new_n806), .B2(new_n448), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n801), .B1(new_n807), .B2(KEYINPUT108), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n681), .A2(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n808), .A2(new_n810), .A3(KEYINPUT109), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT109), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n648), .A2(new_n594), .A3(new_n649), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n681), .B2(new_n809), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n807), .A2(KEYINPUT108), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n798), .B(new_n793), .C1(new_n811), .C2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n593), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT109), .B1(new_n808), .B2(new_n810), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n814), .A2(new_n812), .A3(new_n815), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT42), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n793), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n817), .A2(KEYINPUT42), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G131), .ZN(G33));
  INV_X1    g639(.A(new_n718), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n593), .B(new_n826), .C1(new_n811), .C2(new_n816), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G134), .ZN(G36));
  INV_X1    g642(.A(new_n670), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n253), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT43), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(KEYINPUT44), .A3(new_n683), .A4(new_n710), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n832), .A2(new_n801), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n426), .B1(new_n678), .B2(new_n679), .ZN(new_n834));
  OAI21_X1  g648(.A(G469), .B1(new_n834), .B2(KEYINPUT45), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT45), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n836), .B(new_n426), .C1(new_n678), .C2(new_n679), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n454), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT46), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n840), .A2(new_n841), .B1(new_n449), .B2(new_n805), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n839), .A2(KEYINPUT46), .A3(new_n454), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n328), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n831), .A2(new_n683), .A3(new_n710), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT44), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n833), .A2(new_n736), .A3(new_n844), .A4(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(G137), .ZN(G39));
  NOR4_X1   g663(.A1(new_n722), .A2(new_n813), .A3(new_n759), .A4(new_n749), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n844), .A2(KEYINPUT47), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n844), .A2(KEYINPUT47), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(G140), .ZN(G42));
  AND4_X1   g668(.A1(new_n759), .A2(new_n831), .A3(new_n320), .A4(new_n780), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n742), .A2(new_n594), .A3(new_n788), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT50), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n844), .A2(KEYINPUT47), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n844), .A2(KEYINPUT47), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n761), .A2(new_n452), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n859), .B(new_n860), .C1(new_n329), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n855), .A2(new_n801), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n858), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n733), .A2(new_n759), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n252), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n868), .A2(new_n245), .B1(G475), .B2(new_n223), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n801), .A2(new_n762), .A3(new_n320), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n867), .A2(new_n869), .A3(new_n829), .A4(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n831), .A3(new_n787), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT112), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT51), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n873), .B2(new_n874), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n865), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n855), .A2(new_n789), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n867), .A2(new_n672), .A3(new_n870), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n798), .A2(new_n831), .A3(new_n870), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n881), .A2(KEYINPUT48), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(KEYINPUT48), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n877), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n873), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT51), .B1(new_n865), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n253), .A2(new_n318), .A3(new_n324), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n807), .A2(new_n801), .A3(new_n889), .A4(new_n717), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n769), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n821), .B2(new_n826), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n787), .B(new_n793), .C1(new_n811), .C2(new_n816), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT111), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n891), .ZN(new_n895));
  AND4_X1   g709(.A1(KEYINPUT111), .A2(new_n827), .A3(new_n893), .A4(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AND4_X1   g711(.A1(new_n655), .A2(new_n762), .A3(new_n791), .A4(new_n792), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n571), .A2(new_n574), .B1(G472), .B2(new_n591), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n899), .A2(new_n681), .A3(new_n724), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n898), .A2(new_n787), .B1(new_n900), .B2(new_n719), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT52), .ZN(new_n902));
  INV_X1    g716(.A(new_n699), .ZN(new_n903));
  INV_X1    g717(.A(new_n701), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n697), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n515), .B1(new_n905), .B2(new_n702), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n757), .B2(new_n758), .ZN(new_n907));
  AND4_X1   g721(.A1(new_n329), .A2(new_n455), .A3(new_n907), .A4(new_n717), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n724), .A2(new_n744), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n575), .A2(new_n732), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n901), .A2(new_n902), .A3(new_n751), .A4(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n726), .A2(new_n751), .A3(new_n794), .A4(new_n911), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT52), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n455), .A2(new_n759), .A3(new_n329), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n869), .B1(new_n324), .B2(new_n318), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n323), .B1(new_n916), .B2(new_n671), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n915), .A2(new_n917), .A3(new_n711), .A4(new_n650), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n712), .A2(new_n651), .A3(new_n918), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n769), .A2(new_n770), .B1(new_n781), .B2(new_n782), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n763), .B1(new_n673), .B2(new_n691), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n824), .A2(new_n912), .A3(new_n914), .A4(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n901), .A2(new_n902), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(KEYINPUT53), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n897), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n827), .A2(new_n893), .A3(new_n895), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT111), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n892), .A2(KEYINPUT111), .A3(new_n893), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n817), .A2(KEYINPUT42), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n821), .A2(new_n823), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n922), .A2(new_n912), .A3(new_n914), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT53), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT54), .B1(new_n926), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT53), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n897), .B2(new_n923), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n924), .A2(new_n939), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n931), .A2(new_n936), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n888), .A2(new_n938), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT113), .ZN(new_n946));
  OAI21_X1  g760(.A(G953), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n319), .A2(G953), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n945), .B2(KEYINPUT113), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n861), .A2(KEYINPUT49), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n861), .A2(KEYINPUT49), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n951), .A2(new_n830), .A3(new_n594), .A4(new_n329), .ZN(new_n952));
  OR4_X1    g766(.A1(new_n742), .A2(new_n866), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n947), .A2(new_n949), .A3(new_n953), .ZN(G75));
  AOI21_X1  g768(.A(new_n187), .B1(new_n940), .B2(new_n943), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n647), .ZN(new_n956));
  INV_X1    g770(.A(new_n618), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(KEYINPUT114), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(KEYINPUT114), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT55), .Z(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(new_n628), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT56), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n956), .A2(KEYINPUT115), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT115), .B1(new_n956), .B2(new_n964), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n200), .A2(G952), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT56), .B1(new_n955), .B2(G210), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n962), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n967), .A2(new_n971), .ZN(G51));
  XNOR2_X1  g786(.A(new_n453), .B(KEYINPUT57), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n931), .A2(new_n936), .A3(new_n942), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n974), .A2(new_n937), .A3(KEYINPUT54), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n941), .B1(new_n940), .B2(new_n943), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT116), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n803), .A2(new_n804), .ZN(new_n980));
  OAI211_X1 g794(.A(KEYINPUT116), .B(new_n973), .C1(new_n975), .C2(new_n976), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n955), .A2(new_n838), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n968), .B1(new_n982), .B2(new_n983), .ZN(G54));
  NAND3_X1  g798(.A1(new_n955), .A2(KEYINPUT58), .A3(G475), .ZN(new_n985));
  INV_X1    g799(.A(new_n251), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n987), .A2(new_n988), .A3(new_n968), .ZN(G60));
  NAND2_X1  g803(.A1(G478), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT59), .Z(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(new_n938), .B2(new_n944), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n661), .A2(new_n663), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n969), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n991), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n993), .B(new_n995), .C1(new_n975), .C2(new_n976), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(KEYINPUT117), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(KEYINPUT117), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(G63));
  NAND2_X1  g813(.A1(G217), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT60), .Z(new_n1001));
  OAI21_X1  g815(.A(new_n1001), .B1(new_n974), .B2(new_n937), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n968), .B1(new_n1002), .B2(new_n513), .ZN(new_n1003));
  AOI21_X1  g817(.A(KEYINPUT61), .B1(new_n1003), .B2(KEYINPUT119), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n703), .A2(new_n704), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT118), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1003), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  OAI221_X1 g822(.A(new_n1003), .B1(KEYINPUT119), .B2(KEYINPUT61), .C1(new_n1002), .C2(new_n1006), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(G66));
  OAI21_X1  g824(.A(G953), .B1(new_n624), .B2(new_n322), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1011), .B1(new_n922), .B2(G953), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n958), .B(new_n959), .C1(G898), .C2(new_n200), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT120), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1012), .B(new_n1014), .ZN(G69));
  NAND2_X1  g829(.A1(new_n529), .A2(new_n545), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n237), .B(KEYINPUT121), .Z(new_n1017));
  XNOR2_X1  g831(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT122), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n901), .A2(new_n751), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n747), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT62), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n916), .A2(new_n671), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n593), .A2(new_n737), .A3(new_n801), .A4(new_n1024), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n848), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n853), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1019), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1021), .B(KEYINPUT62), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1029), .A2(KEYINPUT122), .A3(new_n853), .A4(new_n1026), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1018), .B1(new_n1031), .B2(new_n200), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n200), .B1(G227), .B2(G900), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1018), .B1(new_n715), .B2(new_n200), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1020), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n844), .A2(new_n736), .A3(new_n909), .A4(new_n798), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n853), .A2(new_n848), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n824), .A2(new_n827), .ZN(new_n1038));
  OR2_X1    g852(.A1(new_n1038), .A2(KEYINPUT123), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(KEYINPUT123), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1034), .B1(new_n1041), .B2(new_n200), .ZN(new_n1042));
  OR3_X1    g856(.A1(new_n1032), .A2(new_n1033), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1033), .B1(new_n1032), .B2(new_n1042), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1043), .A2(new_n1044), .ZN(G72));
  XNOR2_X1  g859(.A(new_n576), .B(KEYINPUT125), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(new_n553), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1028), .A2(new_n922), .A3(new_n1030), .ZN(new_n1048));
  NAND2_X1  g862(.A1(G472), .A2(G902), .ZN(new_n1049));
  XOR2_X1   g863(.A(new_n1049), .B(KEYINPUT63), .Z(new_n1050));
  NAND2_X1  g864(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1051), .A2(KEYINPUT124), .ZN(new_n1052));
  INV_X1    g866(.A(KEYINPUT124), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1048), .A2(new_n1053), .A3(new_n1050), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1047), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g869(.A1(new_n1046), .A2(new_n553), .ZN(new_n1056));
  AND2_X1   g870(.A1(new_n1041), .A2(new_n922), .ZN(new_n1057));
  INV_X1    g871(.A(new_n1050), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n1058), .B1(new_n577), .B2(new_n554), .ZN(new_n1060));
  XOR2_X1   g874(.A(new_n1060), .B(KEYINPUT126), .Z(new_n1061));
  OAI21_X1  g875(.A(new_n1061), .B1(new_n926), .B2(new_n937), .ZN(new_n1062));
  NAND3_X1  g876(.A1(new_n1059), .A2(new_n969), .A3(new_n1062), .ZN(new_n1063));
  NOR2_X1   g877(.A1(new_n1055), .A2(new_n1063), .ZN(G57));
endmodule


