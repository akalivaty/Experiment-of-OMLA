//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1262, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(new_n202), .A2(new_n203), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n203), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n214), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n213), .B(new_n217), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  NAND2_X1  g0047(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT8), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G58), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n251), .A2(new_n253), .B1(G150), .B2(new_n254), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n255), .A2(KEYINPUT68), .B1(new_n204), .B2(G20), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(KEYINPUT68), .B2(new_n255), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n210), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(new_n211), .A3(G1), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n259), .ZN(new_n263));
  INV_X1    g0063(.A(G50), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(G20), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n263), .A2(new_n266), .B1(new_n264), .B2(new_n262), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT9), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  OAI211_X1 g0070(.A(G1), .B(G13), .C1(new_n252), .C2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(G274), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G226), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G222), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G223), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n283), .B1(new_n220), .B2(new_n281), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(G200), .B2(new_n289), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n269), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT10), .ZN(new_n294));
  INV_X1    g0094(.A(new_n289), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT69), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n268), .B1(new_n295), .B2(G169), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT17), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n252), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n281), .B2(KEYINPUT73), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n285), .A2(G1698), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT76), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G87), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT73), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT73), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(new_n309), .A3(G33), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(G226), .A3(G1698), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT76), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n317), .A3(new_n305), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n307), .A2(new_n308), .A3(new_n316), .A4(new_n318), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n319), .A2(KEYINPUT77), .A3(new_n287), .ZN(new_n320));
  AOI21_X1  g0120(.A(KEYINPUT77), .B1(new_n319), .B2(new_n287), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n276), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(KEYINPUT78), .A3(G232), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT78), .ZN(new_n325));
  INV_X1    g0125(.A(G232), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n276), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n327), .A3(new_n274), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(G190), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n319), .A2(new_n287), .ZN(new_n331));
  INV_X1    g0131(.A(new_n328), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n322), .A2(new_n329), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n258), .A2(new_n210), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G58), .A2(G68), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n207), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(KEYINPUT74), .A3(G20), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n254), .A2(G159), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n211), .B1(new_n207), .B2(new_n336), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(KEYINPUT74), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT7), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n281), .A2(new_n344), .A3(G20), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n310), .A2(new_n311), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT7), .B1(new_n346), .B2(new_n211), .ZN(new_n347));
  OAI21_X1  g0147(.A(G68), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT16), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n335), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT7), .B1(new_n315), .B2(G20), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n312), .A2(new_n344), .A3(new_n211), .A4(new_n314), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(G68), .A3(new_n353), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n340), .A2(new_n342), .A3(new_n350), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT75), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n356), .B1(new_n354), .B2(new_n355), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n351), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n263), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n265), .A2(G20), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n251), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n262), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n360), .A2(new_n362), .B1(new_n363), .B2(new_n251), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n359), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n302), .B1(new_n334), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT77), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n331), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n319), .A2(KEYINPUT77), .A3(new_n287), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(new_n370), .A3(new_n329), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n333), .A2(new_n330), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n344), .B1(new_n304), .B2(new_n211), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n353), .A2(G68), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n342), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n377), .A2(KEYINPUT16), .A3(new_n339), .A4(new_n338), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT75), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n364), .B1(new_n381), .B2(new_n351), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n373), .A2(KEYINPUT17), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n328), .A2(G179), .ZN(new_n384));
  INV_X1    g0184(.A(G169), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n322), .A2(new_n384), .B1(new_n385), .B2(new_n333), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT18), .B1(new_n386), .B2(new_n366), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n369), .A2(new_n370), .A3(new_n384), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n333), .A2(new_n385), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n390), .A2(new_n382), .A3(new_n391), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n367), .B(new_n383), .C1(new_n387), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n253), .A2(G77), .ZN(new_n394));
  INV_X1    g0194(.A(new_n254), .ZN(new_n395));
  OAI221_X1 g0195(.A(new_n394), .B1(new_n211), .B2(G68), .C1(new_n264), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n259), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT11), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n262), .A2(new_n203), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT12), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT71), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n263), .A2(G68), .A3(new_n361), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n405), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT71), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n401), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT72), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n409), .B(new_n410), .ZN(new_n411));
  XOR2_X1   g0211(.A(new_n274), .B(KEYINPUT70), .Z(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G97), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n326), .A2(G1698), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(G226), .B2(G1698), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n413), .B1(new_n415), .B2(new_n346), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(new_n287), .B1(new_n323), .B2(G238), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT13), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT13), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n412), .A2(new_n420), .A3(new_n417), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT14), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(G169), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n296), .B2(new_n422), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n423), .B1(new_n422), .B2(G169), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n411), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n409), .A2(KEYINPUT72), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n409), .A2(KEYINPUT72), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n419), .A2(G190), .A3(new_n421), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n422), .A2(G200), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  XOR2_X1   g0234(.A(KEYINPUT15), .B(G87), .Z(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n253), .ZN(new_n436));
  INV_X1    g0236(.A(new_n251), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n436), .B1(new_n211), .B2(new_n220), .C1(new_n395), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n259), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n263), .A2(G77), .A3(new_n361), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n440), .C1(G77), .C2(new_n363), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n274), .B1(new_n276), .B2(new_n221), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n281), .A2(G232), .A3(new_n282), .ZN(new_n443));
  INV_X1    g0243(.A(G107), .ZN(new_n444));
  OAI221_X1 g0244(.A(new_n443), .B1(new_n444), .B2(new_n281), .C1(new_n284), .C2(new_n219), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n442), .B1(new_n445), .B2(new_n287), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n441), .B1(G169), .B2(new_n446), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n446), .A2(new_n296), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n441), .B1(G190), .B2(new_n446), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n330), .B2(new_n446), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n301), .A2(new_n393), .A3(new_n434), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n444), .A2(KEYINPUT23), .A3(G20), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT23), .B1(new_n444), .B2(G20), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G116), .ZN(new_n458));
  OAI22_X1  g0258(.A1(new_n456), .A2(new_n457), .B1(G20), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n281), .A2(new_n211), .A3(G87), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n315), .A2(KEYINPUT22), .A3(new_n211), .A4(G87), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT24), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT24), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n462), .A2(new_n466), .A3(new_n463), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n335), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n262), .A2(new_n444), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT25), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n469), .B(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n263), .B1(G1), .B2(new_n252), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n444), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n270), .A2(KEYINPUT5), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n265), .B(G45), .C1(new_n270), .C2(KEYINPUT5), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n287), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G264), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(G1698), .B1(new_n312), .B2(new_n314), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT92), .B(G294), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n483), .A2(G250), .B1(G33), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n315), .A2(G257), .A3(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n482), .B1(new_n488), .B2(new_n287), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT83), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n478), .B1(new_n490), .B2(new_n477), .ZN(new_n491));
  INV_X1    g0291(.A(G274), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n287), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT84), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n476), .A2(KEYINPUT83), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n491), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  OR2_X1    g0296(.A1(new_n270), .A2(KEYINPUT5), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n490), .A2(new_n270), .A3(KEYINPUT5), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n272), .A2(G1), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n495), .A2(new_n497), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n271), .A2(G274), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT84), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n489), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(KEYINPUT93), .A3(G169), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n271), .B1(new_n486), .B2(new_n487), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n496), .A2(new_n502), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n506), .A2(new_n507), .A3(new_n482), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G179), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT93), .B1(new_n504), .B2(G169), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n475), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(G200), .B1(new_n489), .B2(new_n503), .ZN(new_n513));
  NOR4_X1   g0313(.A1(new_n506), .A2(new_n507), .A3(new_n482), .A4(G190), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n474), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT21), .ZN(new_n517));
  INV_X1    g0317(.A(new_n472), .ZN(new_n518));
  INV_X1    g0318(.A(G116), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n262), .A2(G116), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g0322(.A1(KEYINPUT79), .A2(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(KEYINPUT79), .A2(G97), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n252), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G283), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT81), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT81), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(G33), .A3(G283), .ZN(new_n530));
  AOI21_X1  g0330(.A(G20), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n259), .B1(new_n211), .B2(G116), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT20), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n535), .B(KEYINPUT90), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n532), .A2(new_n534), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT20), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(KEYINPUT91), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT91), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n533), .B1(new_n531), .B2(new_n526), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(KEYINPUT20), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n522), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n304), .A2(new_n282), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(G264), .B1(G303), .B2(new_n346), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n315), .A2(G257), .A3(new_n282), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n271), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n480), .A2(G270), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n503), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(G169), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n517), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT90), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n535), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n539), .A2(new_n542), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n554), .A2(new_n555), .B1(new_n521), .B2(new_n520), .ZN(new_n556));
  INV_X1    g0356(.A(G303), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n315), .A2(G1698), .ZN(new_n558));
  INV_X1    g0358(.A(G264), .ZN(new_n559));
  OAI221_X1 g0359(.A(new_n547), .B1(new_n557), .B2(new_n281), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n287), .ZN(new_n561));
  INV_X1    g0361(.A(new_n550), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n385), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n556), .A2(new_n563), .A3(KEYINPUT21), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(G190), .ZN(new_n565));
  OAI21_X1  g0365(.A(G200), .B1(new_n548), .B2(new_n550), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n544), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n548), .A2(new_n550), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n556), .A2(G179), .A3(new_n568), .ZN(new_n569));
  AND4_X1   g0369(.A1(new_n552), .A2(new_n564), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n528), .A2(new_n530), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n282), .A2(KEYINPUT4), .A3(G244), .ZN(new_n572));
  OR2_X1    g0372(.A1(new_n346), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n282), .A2(G244), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n312), .B2(new_n314), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n571), .B(new_n573), .C1(new_n575), .C2(KEYINPUT4), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n310), .A2(new_n311), .A3(G250), .A4(G1698), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT82), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n577), .B(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n287), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(G257), .B(new_n271), .C1(new_n477), .C2(new_n478), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n496), .B2(new_n502), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(KEYINPUT85), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT85), .ZN(new_n585));
  AOI211_X1 g0385(.A(new_n585), .B(new_n582), .C1(new_n496), .C2(new_n502), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n296), .B(new_n580), .C1(new_n584), .C2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n525), .A2(KEYINPUT6), .A3(new_n444), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT6), .ZN(new_n589));
  XNOR2_X1  g0389(.A(G97), .B(G107), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n588), .A2(KEYINPUT80), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n589), .B(G107), .C1(new_n523), .C2(new_n524), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT80), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n211), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(G107), .B1(new_n345), .B2(new_n347), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n254), .A2(G77), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n259), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n363), .A2(G97), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n518), .B2(G97), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n587), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT86), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n580), .B2(new_n583), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n580), .A2(new_n604), .A3(new_n583), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n385), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n580), .B1(new_n584), .B2(new_n586), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n602), .B1(new_n609), .B2(G200), .ZN(new_n610));
  INV_X1    g0410(.A(new_n607), .ZN(new_n611));
  OAI21_X1  g0411(.A(G190), .B1(new_n611), .B2(new_n605), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n603), .A2(new_n608), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n525), .A2(new_n253), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT19), .ZN(new_n615));
  INV_X1    g0415(.A(G87), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n523), .A2(new_n616), .A3(new_n444), .A4(new_n524), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n211), .B1(new_n413), .B2(new_n615), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n614), .A2(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n315), .A2(new_n211), .A3(G68), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n259), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n363), .A2(new_n435), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(KEYINPUT87), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT87), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n335), .B1(new_n619), .B2(new_n620), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n627), .B2(new_n623), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n518), .A2(new_n435), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n499), .A2(G250), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n499), .A2(new_n492), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n271), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n315), .A2(G238), .A3(new_n282), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n636), .B(new_n458), .C1(new_n558), .C2(new_n221), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n635), .B1(new_n637), .B2(new_n287), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n296), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(G169), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n631), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n638), .A2(new_n290), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(G200), .B2(new_n638), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT88), .B1(new_n472), .B2(new_n616), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT88), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n518), .A2(new_n646), .A3(G87), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n625), .A2(new_n628), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT89), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n642), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n642), .B2(new_n649), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n570), .B(new_n613), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n455), .A2(new_n516), .A3(new_n653), .ZN(G372));
  INV_X1    g0454(.A(new_n300), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n391), .B1(new_n390), .B2(new_n382), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n366), .A2(KEYINPUT18), .A3(new_n388), .A4(new_n389), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g0458(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n433), .A2(new_n449), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n664), .A2(new_n427), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n367), .A2(new_n383), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n655), .B1(new_n667), .B2(new_n294), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n552), .A2(new_n564), .A3(new_n569), .ZN(new_n669));
  INV_X1    g0469(.A(new_n511), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n505), .A2(new_n670), .A3(new_n509), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n669), .B1(new_n671), .B2(new_n475), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n640), .B1(new_n296), .B2(new_n638), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n673), .A2(new_n631), .B1(new_n644), .B2(new_n648), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n603), .A2(new_n608), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n610), .A2(new_n612), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .A4(new_n515), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n642), .B1(new_n672), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n603), .A2(KEYINPUT94), .A3(new_n608), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT94), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n611), .A2(G169), .A3(new_n605), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n587), .A2(new_n602), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n679), .A2(new_n674), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT26), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n675), .ZN(new_n687));
  OAI211_X1 g0487(.A(KEYINPUT26), .B(new_n687), .C1(new_n651), .C2(new_n652), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n678), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n668), .B1(new_n455), .B2(new_n689), .ZN(G369));
  AND2_X1   g0490(.A1(new_n512), .A2(new_n515), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n265), .A2(new_n211), .A3(G13), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(G213), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n691), .B1(new_n474), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n671), .A2(new_n475), .A3(new_n697), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n556), .A2(new_n697), .ZN(new_n703));
  MUX2_X1   g0503(.A(new_n669), .B(new_n570), .S(new_n703), .Z(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n697), .B(KEYINPUT97), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n512), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n669), .A2(new_n698), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n691), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT98), .Z(G399));
  INV_X1    g0514(.A(new_n215), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G41), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n265), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n617), .A2(G116), .ZN(new_n719));
  INV_X1    g0519(.A(new_n716), .ZN(new_n720));
  OAI22_X1  g0520(.A1(new_n718), .A2(new_n719), .B1(new_n208), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  INV_X1    g0522(.A(G330), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n568), .A2(G179), .A3(new_n489), .A4(new_n638), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n611), .A2(new_n605), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT30), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n561), .A2(new_n562), .A3(G179), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n489), .A2(new_n638), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n606), .A2(new_n607), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n638), .A2(G179), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n561), .A2(new_n562), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n609), .A2(new_n734), .A3(new_n504), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT31), .B1(new_n737), .B2(new_n697), .ZN(new_n738));
  INV_X1    g0538(.A(new_n736), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n726), .B2(new_n732), .ZN(new_n740));
  XNOR2_X1  g0540(.A(KEYINPUT99), .B(KEYINPUT31), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n740), .A2(new_n708), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n612), .ZN(new_n744));
  INV_X1    g0544(.A(new_n602), .ZN(new_n745));
  INV_X1    g0545(.A(new_n580), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n585), .B1(new_n507), .B2(new_n582), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n583), .A2(KEYINPUT85), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n745), .B1(new_n749), .B2(new_n330), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n744), .A2(new_n750), .B1(new_n681), .B2(new_n682), .ZN(new_n751));
  INV_X1    g0551(.A(new_n652), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n674), .A2(new_n650), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n754), .A2(new_n691), .A3(new_n570), .A4(new_n708), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n723), .B1(new_n743), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n685), .B(new_n687), .C1(new_n651), .C2(new_n652), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n684), .A2(KEYINPUT26), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g0560(.A(KEYINPUT29), .B(new_n698), .C1(new_n760), .C2(new_n678), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n688), .A2(new_n686), .ZN(new_n762));
  INV_X1    g0562(.A(new_n642), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n642), .A2(new_n515), .A3(new_n649), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n751), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n564), .A2(new_n569), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n512), .A2(new_n552), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n763), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n709), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n761), .B1(new_n769), .B2(KEYINPUT29), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n757), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n722), .B1(new_n772), .B2(G1), .ZN(G364));
  NOR3_X1   g0573(.A1(new_n261), .A2(new_n272), .A3(G20), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT100), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n718), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n704), .B2(G330), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G330), .B2(new_n704), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n715), .A2(new_n346), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G355), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G116), .B2(new_n215), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n315), .A2(new_n715), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(new_n272), .B2(new_n209), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n243), .A2(G45), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G13), .A2(G33), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n210), .B1(G20), .B2(new_n385), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT101), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n776), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT102), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n211), .A2(new_n296), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G190), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n281), .B1(new_n798), .B2(new_n220), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n796), .A2(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n290), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n799), .B1(G50), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n211), .A2(G179), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n803), .A2(G190), .A3(G200), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n616), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n803), .A2(new_n290), .A3(G200), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n805), .B1(G107), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n796), .A2(G190), .A3(new_n330), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT103), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n802), .B(new_n808), .C1(new_n202), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n803), .A2(new_n797), .ZN(new_n812));
  INV_X1    g0612(.A(G159), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(KEYINPUT104), .B(KEYINPUT32), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n290), .A2(G179), .A3(G200), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n211), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n800), .A2(G190), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G97), .A2(new_n819), .B1(new_n820), .B2(G68), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G317), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT33), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n823), .A2(KEYINPUT33), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n820), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n801), .A2(G326), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(new_n557), .C2(new_n804), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n819), .A2(new_n485), .B1(new_n807), .B2(G283), .ZN(new_n829));
  INV_X1    g0629(.A(new_n809), .ZN(new_n830));
  INV_X1    g0630(.A(new_n812), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n830), .A2(G322), .B1(new_n831), .B2(G329), .ZN(new_n832));
  INV_X1    g0632(.A(new_n798), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n281), .B1(new_n833), .B2(G311), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n829), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n811), .A2(new_n822), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n795), .B1(new_n790), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n789), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n837), .B1(new_n794), .B2(new_n793), .C1(new_n704), .C2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n778), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  NAND2_X1  g0641(.A1(new_n441), .A2(new_n697), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n452), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n450), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n449), .A2(new_n698), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n769), .B(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(new_n757), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT106), .Z(new_n850));
  AOI21_X1  g0650(.A(new_n776), .B1(new_n848), .B2(new_n757), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n790), .A2(new_n787), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n776), .B1(G77), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT105), .ZN(new_n856));
  INV_X1    g0656(.A(new_n801), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n857), .A2(new_n557), .B1(new_n806), .B2(new_n616), .ZN(new_n858));
  INV_X1    g0658(.A(new_n804), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(G107), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(G294), .ZN(new_n861));
  INV_X1    g0661(.A(G311), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n809), .A2(new_n861), .B1(new_n812), .B2(new_n862), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n281), .B(new_n863), .C1(G116), .C2(new_n833), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G97), .A2(new_n819), .B1(new_n820), .B2(G283), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n860), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n807), .A2(G68), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n867), .B1(new_n264), .B2(new_n804), .C1(new_n202), .C2(new_n818), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n304), .B(new_n868), .C1(G132), .C2(new_n831), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT34), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n801), .A2(G137), .B1(new_n833), .B2(G159), .ZN(new_n871));
  INV_X1    g0671(.A(G150), .ZN(new_n872));
  INV_X1    g0672(.A(new_n820), .ZN(new_n873));
  INV_X1    g0673(.A(G143), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n871), .B1(new_n872), .B2(new_n873), .C1(new_n810), .C2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n869), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n875), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(KEYINPUT34), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n866), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n856), .B1(new_n879), .B2(new_n790), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n847), .B2(new_n788), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n852), .A2(new_n881), .ZN(G384));
  AOI21_X1  g0682(.A(new_n265), .B1(G13), .B2(new_n211), .ZN(new_n883));
  INV_X1    g0683(.A(new_n695), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n663), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT107), .B1(new_n430), .B2(new_n698), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT107), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n411), .A2(new_n887), .A3(new_n697), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n427), .A2(new_n886), .A3(new_n433), .A4(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n427), .A2(new_n433), .B1(new_n886), .B2(new_n888), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n709), .B(new_n846), .C1(new_n762), .C2(new_n768), .ZN(new_n894));
  INV_X1    g0694(.A(new_n845), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n354), .A2(new_n343), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n335), .B1(new_n898), .B2(new_n350), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n381), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n365), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n386), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n695), .B1(new_n900), .B2(new_n365), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n373), .A2(new_n382), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT37), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n366), .A2(new_n388), .A3(new_n389), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n366), .A2(new_n884), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n907), .B1(KEYINPUT37), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n373), .A2(KEYINPUT17), .A3(new_n382), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT17), .B1(new_n373), .B2(new_n382), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI211_X1 g0714(.A(KEYINPUT108), .B(new_n904), .C1(new_n914), .C2(new_n658), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT108), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n393), .B2(new_n903), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n911), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(KEYINPUT38), .B(new_n911), .C1(new_n915), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n885), .B1(new_n897), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  INV_X1    g0724(.A(new_n921), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT95), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n905), .A2(new_n926), .A3(new_n909), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT37), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n910), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n695), .B1(new_n359), .B2(new_n365), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n382), .B2(new_n373), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n931), .A2(KEYINPUT95), .A3(KEYINPUT37), .A4(new_n908), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n661), .A2(new_n914), .A3(new_n662), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n930), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n924), .B1(new_n925), .B2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n427), .A2(new_n697), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n920), .A2(KEYINPUT39), .A3(new_n921), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n923), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n454), .B(new_n761), .C1(KEYINPUT29), .C2(new_n769), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n668), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n886), .A2(new_n888), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n434), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n846), .B1(new_n947), .B2(new_n889), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n653), .A2(new_n516), .A3(new_n709), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n741), .B1(new_n740), .B2(new_n698), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n948), .B(new_n949), .C1(new_n950), .C2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n922), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n948), .B1(new_n950), .B2(new_n953), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n933), .A2(new_n935), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n919), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n957), .B1(new_n959), .B2(new_n921), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n956), .B1(new_n949), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n950), .A2(new_n953), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n962), .B1(new_n455), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n755), .A2(new_n952), .A3(new_n951), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n961), .A2(new_n454), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(G330), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n883), .B1(new_n945), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n945), .B2(new_n967), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n591), .A2(new_n594), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT35), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT35), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n972), .A2(G116), .A3(new_n212), .A4(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT36), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n209), .A2(G77), .A3(new_n336), .ZN(new_n976));
  INV_X1    g0776(.A(new_n201), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n976), .B1(new_n203), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(G1), .A3(new_n261), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n969), .A2(new_n975), .A3(new_n979), .ZN(G367));
  OAI21_X1  g0780(.A(new_n613), .B1(new_n745), .B2(new_n708), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n687), .A2(new_n709), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n691), .A2(new_n711), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT42), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n675), .B1(new_n981), .B2(new_n512), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT109), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n709), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n989), .B2(new_n988), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n648), .A2(new_n698), .ZN(new_n992));
  MUX2_X1   g0792(.A(new_n674), .B(new_n763), .S(new_n992), .Z(new_n993));
  AOI22_X1  g0793(.A1(new_n987), .A2(new_n991), .B1(KEYINPUT43), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n706), .A2(new_n983), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n775), .A2(new_n265), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n712), .A2(new_n983), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT45), .Z(new_n1001));
  NOR2_X1   g0801(.A1(new_n712), .A2(new_n983), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT44), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(new_n707), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n985), .B1(new_n701), .B2(new_n711), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(new_n705), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n771), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n716), .B(KEYINPUT41), .Z(new_n1010));
  OAI21_X1  g0810(.A(new_n999), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n998), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n792), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n435), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1013), .B1(new_n215), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n783), .A2(new_n239), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n776), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(G283), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n304), .B1(new_n1018), .B2(new_n798), .C1(new_n823), .C2(new_n812), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n810), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(G303), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n859), .A2(G116), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT46), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G107), .A2(new_n819), .B1(new_n820), .B2(new_n485), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n801), .A2(G311), .B1(new_n807), .B2(new_n525), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT110), .Z(new_n1027));
  NOR2_X1   g0827(.A1(new_n818), .A2(new_n203), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G150), .B2(new_n830), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT111), .ZN(new_n1030));
  INV_X1    g0830(.A(G137), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n804), .A2(new_n202), .B1(new_n812), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1032), .A2(KEYINPUT112), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n873), .A2(new_n813), .B1(new_n857), .B2(new_n874), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1032), .A2(KEYINPUT112), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n807), .A2(G77), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1036), .B(new_n281), .C1(new_n201), .C2(new_n798), .ZN(new_n1037));
  OR4_X1    g0837(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1027), .B1(new_n1030), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT47), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1017), .B1(new_n1040), .B2(new_n790), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n838), .B2(new_n993), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1012), .A2(new_n1042), .ZN(G387));
  OAI22_X1  g0843(.A1(new_n809), .A2(new_n264), .B1(new_n798), .B2(new_n203), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(KEYINPUT113), .B(G150), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1044), .B1(new_n831), .B2(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n820), .A2(new_n251), .B1(new_n859), .B2(G77), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n819), .A2(new_n435), .B1(new_n807), .B2(G97), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n304), .B1(new_n801), .B2(G159), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n315), .B1(G326), .B2(new_n831), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n820), .A2(G311), .B1(new_n833), .B2(G303), .ZN(new_n1053));
  INV_X1    g0853(.A(G322), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n857), .C1(new_n810), .C2(new_n823), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n819), .A2(G283), .B1(new_n859), .B2(new_n485), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT49), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1052), .B1(new_n519), .B2(new_n806), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1051), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n790), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n776), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n236), .A2(new_n272), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1067), .A2(new_n782), .B1(new_n719), .B2(new_n779), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n251), .A2(new_n264), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT50), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n272), .B1(new_n203), .B2(new_n220), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n1070), .A2(new_n719), .A3(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1068), .A2(new_n1072), .B1(G107), .B2(new_n215), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1066), .B1(new_n1073), .B2(new_n1013), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1065), .B(new_n1074), .C1(new_n701), .C2(new_n838), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1007), .A2(new_n771), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n716), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1008), .A2(new_n772), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1075), .B1(new_n1007), .B2(new_n999), .C1(new_n1078), .C2(new_n1079), .ZN(G393));
  AOI21_X1  g0880(.A(new_n792), .B1(new_n715), .B2(new_n525), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n783), .A2(new_n246), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1066), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n790), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n873), .A2(new_n201), .B1(new_n616), .B2(new_n806), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n315), .B1(new_n874), .B2(new_n812), .C1(new_n437), .C2(new_n798), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n804), .A2(new_n203), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n818), .A2(new_n220), .ZN(new_n1089));
  NOR4_X1   g0889(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n857), .A2(new_n872), .B1(new_n813), .B2(new_n809), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n857), .A2(new_n823), .B1(new_n862), .B2(new_n809), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT52), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n873), .A2(new_n557), .B1(new_n806), .B2(new_n444), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n346), .B1(new_n812), .B2(new_n1054), .C1(new_n861), .C2(new_n798), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n818), .A2(new_n519), .B1(new_n804), .B2(new_n1018), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1090), .A2(new_n1092), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1084), .B1(new_n1085), .B2(new_n1099), .C1(new_n983), .C2(new_n838), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1004), .B(new_n706), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(new_n999), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1077), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT114), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n720), .B1(new_n1005), .B2(new_n1076), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G390));
  OAI21_X1  g0907(.A(new_n847), .B1(new_n890), .B2(new_n891), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n963), .A2(new_n1108), .A3(new_n723), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n937), .A2(new_n940), .B1(new_n896), .B2(new_n938), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n698), .B(new_n844), .C1(new_n760), .C2(new_n678), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n845), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n893), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n929), .A2(new_n932), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n930), .B2(new_n934), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n921), .B1(new_n1115), .B2(KEYINPUT38), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1113), .A2(new_n938), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1109), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n895), .B1(new_n769), .B2(new_n847), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n938), .B1(new_n1119), .B2(new_n892), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n920), .A2(KEYINPUT39), .A3(new_n921), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT39), .B1(new_n959), .B2(new_n921), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1113), .A2(new_n938), .A3(new_n1116), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n756), .A2(new_n847), .A3(new_n893), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n454), .A2(new_n965), .A3(G330), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n943), .A2(new_n668), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n893), .B1(new_n756), .B2(new_n847), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n1129), .A2(new_n1109), .B1(new_n895), .B2(new_n894), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1111), .A2(new_n845), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n963), .A2(new_n723), .A3(new_n846), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1125), .B(new_n1131), .C1(new_n1132), .C2(new_n893), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1128), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1118), .A2(new_n1126), .A3(new_n1134), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1135), .A2(new_n716), .ZN(new_n1136));
  AOI211_X1 g0936(.A(KEYINPUT115), .B(new_n1134), .C1(new_n1118), .C2(new_n1126), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT115), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1118), .A2(new_n1126), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1134), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1136), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n999), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1118), .A2(new_n1126), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n787), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n776), .B1(new_n251), .B2(new_n854), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n859), .A2(new_n1046), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT53), .ZN(new_n1148));
  INV_X1    g0948(.A(G125), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n281), .B1(new_n812), .B2(new_n1149), .C1(new_n798), .C2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n873), .A2(new_n1031), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n818), .A2(new_n813), .B1(new_n806), .B2(new_n201), .ZN(new_n1153));
  OR4_X1    g0953(.A1(new_n1148), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G128), .A2(new_n801), .B1(new_n830), .B2(G132), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT116), .Z(new_n1156));
  NAND2_X1  g0956(.A1(new_n833), .A2(new_n525), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n873), .B2(new_n444), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT117), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1089), .B1(G283), .B2(new_n801), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n830), .A2(G116), .B1(new_n831), .B2(G294), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n867), .A4(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(KEYINPUT118), .B(new_n346), .C1(new_n804), .C2(new_n616), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT118), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n805), .B2(new_n281), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n1154), .A2(new_n1156), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1146), .B1(new_n1168), .B2(new_n790), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1145), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1142), .A2(new_n1144), .A3(new_n1170), .ZN(G378));
  AOI21_X1  g0971(.A(new_n301), .B1(new_n268), .B2(new_n884), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n268), .A2(new_n884), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n294), .B2(new_n300), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OR3_X1    g0976(.A1(new_n1172), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1176), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n961), .B2(G330), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n963), .A2(new_n1108), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n949), .B1(new_n1116), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n954), .B1(new_n920), .B2(new_n921), .ZN(new_n1183));
  OAI211_X1 g0983(.A(G330), .B(new_n1179), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n942), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(G330), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1179), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1189), .A2(new_n941), .A3(new_n923), .A4(new_n1184), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n999), .B1(new_n1186), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1066), .B1(new_n201), .B2(new_n853), .ZN(new_n1192));
  INV_X1    g0992(.A(G132), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n873), .A2(new_n1193), .B1(new_n857), .B2(new_n1149), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n830), .A2(G128), .B1(new_n833), .B2(G137), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n804), .B2(new_n1150), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(G150), .C2(new_n819), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n807), .A2(G159), .ZN(new_n1201));
  AOI211_X1 g1001(.A(G33), .B(G41), .C1(new_n831), .C2(G124), .ZN(new_n1202));
  AND4_X1   g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n830), .A2(G107), .B1(new_n831), .B2(G283), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1014), .B2(new_n798), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1028), .B(new_n1205), .C1(G77), .C2(new_n859), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n857), .A2(new_n519), .B1(new_n806), .B2(new_n202), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G97), .B2(new_n820), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n315), .A2(G41), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G50), .B(new_n1209), .C1(new_n252), .C2(new_n270), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(new_n1203), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1192), .B1(new_n1085), .B2(new_n1215), .C1(new_n1179), .C2(new_n788), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT120), .Z(new_n1217));
  NOR2_X1   g1017(.A1(new_n1191), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1128), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1186), .A2(new_n1190), .B1(new_n1135), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n716), .B1(new_n1220), .B2(KEYINPUT57), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1186), .A2(new_n1190), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1135), .A2(new_n1219), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1222), .A2(KEYINPUT57), .A3(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1218), .B1(new_n1221), .B2(new_n1224), .ZN(G375));
  NAND2_X1  g1025(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1143), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n873), .A2(new_n519), .B1(new_n857), .B2(new_n861), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G97), .B2(new_n859), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n819), .A2(new_n435), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n809), .A2(new_n1018), .B1(new_n798), .B2(new_n444), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n281), .B(new_n1231), .C1(G303), .C2(new_n831), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1229), .A2(new_n1036), .A3(new_n1230), .A4(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n819), .A2(G50), .B1(new_n859), .B2(G159), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1193), .B2(new_n857), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1020), .A2(G137), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G150), .A2(new_n833), .B1(new_n831), .B2(G128), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1150), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n820), .A2(new_n1238), .B1(new_n807), .B2(G58), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n315), .A3(new_n1237), .A4(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1233), .B1(new_n1235), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n790), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1066), .B1(new_n203), .B2(new_n853), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(new_n893), .C2(new_n788), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1227), .A2(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT121), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1010), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1130), .A2(new_n1133), .A3(new_n1128), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1140), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1246), .A2(new_n1249), .ZN(G381));
  OR4_X1    g1050(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1251));
  OR2_X1    g1051(.A1(G378), .A2(KEYINPUT122), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT57), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n720), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1220), .A2(KEYINPUT57), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G378), .A2(KEYINPUT122), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1252), .A2(new_n1218), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OR4_X1    g1059(.A1(G387), .A2(new_n1251), .A3(G381), .A4(new_n1259), .ZN(G407));
  NAND2_X1  g1060(.A1(new_n696), .A2(G213), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT123), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G407), .B(G213), .C1(new_n1259), .C2(new_n1263), .ZN(G409));
  OR2_X1    g1064(.A1(G387), .A2(new_n1106), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G387), .A2(new_n1106), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(G393), .B(new_n840), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1265), .A2(new_n1266), .A3(new_n1268), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT124), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1142), .A2(new_n1144), .A3(new_n1170), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(G375), .B2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1257), .A2(KEYINPUT124), .A3(G378), .A4(new_n1218), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1218), .B1(new_n1010), .B2(new_n1253), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1252), .A2(new_n1258), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1262), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT60), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1248), .B1(new_n1134), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT125), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT125), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1285), .B(new_n1248), .C1(new_n1134), .C2(new_n1282), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1248), .A2(new_n1282), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1287), .A2(new_n720), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1284), .A2(new_n1286), .A3(new_n1288), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1246), .A2(G384), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G384), .B1(new_n1246), .B2(new_n1289), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1273), .B1(new_n1281), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1261), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT126), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1262), .A2(G2897), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1246), .A2(new_n1289), .ZN(new_n1300));
  INV_X1    g1100(.A(G384), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1246), .A2(G384), .A3(new_n1289), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n696), .A2(G213), .A3(G2897), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1302), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1297), .B1(new_n1299), .B2(new_n1305), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1299), .A2(new_n1305), .A3(new_n1297), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1296), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1295), .A2(new_n1261), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1292), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1294), .A2(new_n1308), .A3(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1307), .A2(new_n1306), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1271), .B1(new_n1281), .B2(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1310), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1281), .A2(KEYINPUT62), .A3(new_n1309), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1314), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1312), .B1(new_n1318), .B2(new_n1320), .ZN(G405));
  NAND3_X1  g1121(.A1(new_n1252), .A2(G375), .A3(new_n1258), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1278), .A2(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1323), .A2(new_n1309), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1309), .ZN(new_n1325));
  OR3_X1    g1125(.A1(new_n1324), .A2(new_n1325), .A3(new_n1319), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1319), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(G402));
endmodule


