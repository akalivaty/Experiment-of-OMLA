//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n205), .A2(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  OR3_X1    g009(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n210), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(new_n207), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(KEYINPUT17), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT86), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  AOI21_X1  g018(.A(G1gat), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT84), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(KEYINPUT85), .A2(G8gat), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n218), .B(new_n221), .C1(new_n219), .C2(G1gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(KEYINPUT85), .A2(G8gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n214), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n217), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n228), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n229), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT87), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(KEYINPUT18), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n235), .B(KEYINPUT88), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(KEYINPUT13), .ZN(new_n241));
  INV_X1    g040(.A(new_n234), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n233), .A2(new_n229), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n238), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n232), .A2(new_n234), .A3(new_n235), .A4(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n239), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT11), .B(G169gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G197gat), .ZN(new_n249));
  XOR2_X1   g048(.A(G113gat), .B(G141gat), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n251), .B(KEYINPUT83), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT12), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n253), .A2(new_n239), .A3(new_n244), .A4(new_n246), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259));
  XNOR2_X1  g058(.A(G127gat), .B(G134gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT70), .B(G113gat), .ZN(new_n261));
  INV_X1    g060(.A(G120gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n262), .A2(G113gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n259), .B(new_n260), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G113gat), .B(G120gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(KEYINPUT1), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n267), .A2(new_n260), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT26), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n272), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n276), .B1(KEYINPUT26), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n274), .A2(new_n275), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT27), .B(G183gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT28), .B1(new_n283), .B2(G190gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT27), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G183gat), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT28), .B1(new_n286), .B2(KEYINPUT67), .ZN(new_n287));
  INV_X1    g086(.A(G190gat), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n287), .B(new_n288), .C1(KEYINPUT67), .C2(new_n282), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n284), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n284), .A2(new_n289), .A3(KEYINPUT68), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n281), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n297), .A2(G169gat), .A3(G176gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n299));
  INV_X1    g098(.A(new_n271), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G169gat), .ZN(new_n302));
  INV_X1    g101(.A(G176gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT23), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT64), .B1(new_n304), .B2(new_n271), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n297), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(G183gat), .A3(G190gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n311));
  AND2_X1   g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT25), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n310), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT65), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n306), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n299), .B1(new_n298), .B2(new_n300), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n304), .A2(KEYINPUT64), .A3(new_n271), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G183gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n288), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(KEYINPUT24), .A3(new_n279), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n323), .A2(KEYINPUT25), .A3(new_n307), .A4(new_n309), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT65), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n317), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n313), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n298), .A2(new_n300), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT25), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n296), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  AOI211_X1 g130(.A(KEYINPUT66), .B(new_n329), .C1(new_n317), .C2(new_n325), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n270), .B(new_n295), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT71), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n316), .B1(new_n306), .B2(new_n315), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n320), .A2(new_n324), .A3(KEYINPUT65), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n330), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT66), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n329), .B1(new_n317), .B2(new_n325), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n296), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT71), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n341), .A2(new_n342), .A3(new_n270), .A4(new_n295), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n295), .B1(new_n331), .B2(new_n332), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n269), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n334), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT32), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT33), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G15gat), .B(G43gat), .ZN(new_n353));
  INV_X1    g152(.A(G71gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  XOR2_X1   g154(.A(KEYINPUT72), .B(G99gat), .Z(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  NAND3_X1  g156(.A1(new_n350), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n334), .A2(new_n343), .A3(new_n345), .A4(new_n347), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT73), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT34), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT34), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(KEYINPUT73), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT32), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n346), .B2(new_n348), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT33), .B1(new_n346), .B2(new_n348), .ZN(new_n367));
  INV_X1    g166(.A(new_n357), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n358), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n358), .A2(new_n364), .A3(KEYINPUT74), .A4(new_n369), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(G141gat), .B(G148gat), .Z(new_n375));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT2), .ZN(new_n378));
  XNOR2_X1  g177(.A(G141gat), .B(G148gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT77), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(G155gat), .B(G162gat), .Z(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G155gat), .ZN(new_n384));
  INV_X1    g183(.A(G162gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n378), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(new_n384), .B2(new_n385), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n375), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT4), .B1(new_n389), .B2(new_n269), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n381), .A2(new_n382), .B1(new_n387), .B2(new_n375), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n270), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n389), .B2(new_n269), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n389), .A2(KEYINPUT3), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n269), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n394), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n270), .A2(new_n392), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n389), .A2(new_n269), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n396), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n405), .A3(KEYINPUT5), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n396), .A2(KEYINPUT5), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n394), .A2(new_n401), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT0), .B(G57gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(G85gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n411), .B(new_n412), .Z(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n406), .A2(new_n408), .A3(new_n413), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n409), .A2(KEYINPUT6), .A3(new_n414), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G226gat), .A2(G233gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n422), .B(new_n295), .C1(new_n331), .C2(new_n332), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(KEYINPUT29), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(new_n294), .B2(new_n339), .ZN(new_n425));
  XNOR2_X1  g224(.A(G197gat), .B(G204gat), .ZN(new_n426));
  AND2_X1   g225(.A1(G211gat), .A2(G218gat), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(KEYINPUT22), .B2(new_n427), .ZN(new_n428));
  XOR2_X1   g227(.A(G211gat), .B(G218gat), .Z(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G8gat), .B(G36gat), .Z(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(G64gat), .ZN(new_n433));
  INV_X1    g232(.A(G92gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n294), .A2(new_n339), .A3(new_n421), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n436), .B1(new_n344), .B2(new_n424), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n431), .B(new_n435), .C1(new_n437), .C2(new_n430), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT30), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n431), .B1(new_n437), .B2(new_n430), .ZN(new_n440));
  INV_X1    g239(.A(new_n435), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(KEYINPUT30), .A3(new_n441), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT76), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n440), .A2(KEYINPUT76), .A3(KEYINPUT30), .A4(new_n441), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n420), .A2(new_n443), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n358), .A2(new_n369), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n361), .A2(new_n363), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT29), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n430), .B1(new_n400), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT3), .B1(new_n430), .B2(new_n453), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n392), .ZN(new_n456));
  NAND2_X1  g255(.A1(G228gat), .A2(G233gat), .ZN(new_n457));
  OR3_X1    g256(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(KEYINPUT79), .Z(new_n459));
  NAND3_X1  g258(.A1(new_n428), .A2(KEYINPUT80), .A3(new_n429), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n453), .B(new_n460), .C1(new_n430), .C2(KEYINPUT80), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n392), .B1(new_n461), .B2(new_n399), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n459), .B1(new_n462), .B2(new_n454), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G22gat), .ZN(new_n465));
  INV_X1    g264(.A(G22gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n458), .A2(new_n466), .A3(new_n463), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT81), .ZN(new_n469));
  XNOR2_X1  g268(.A(G78gat), .B(G106gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT78), .ZN(new_n471));
  XOR2_X1   g270(.A(KEYINPUT31), .B(G50gat), .Z(new_n472));
  XOR2_X1   g271(.A(new_n471), .B(new_n472), .Z(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT81), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n465), .A2(new_n475), .A3(new_n467), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n469), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n468), .A2(KEYINPUT81), .A3(new_n473), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n374), .A2(new_n449), .A3(new_n452), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT75), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n484));
  AOI221_X4 g283(.A(new_n365), .B1(KEYINPUT33), .B2(new_n357), .C1(new_n346), .C2(new_n348), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n451), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n483), .B1(new_n450), .B2(new_n451), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n449), .A4(new_n374), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n482), .B1(new_n491), .B2(new_n479), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n374), .A2(new_n452), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT36), .ZN(new_n494));
  INV_X1    g293(.A(new_n488), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n374), .A2(new_n495), .A3(new_n496), .A4(new_n486), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n446), .A2(new_n443), .A3(new_n447), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT39), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n395), .B1(new_n394), .B2(new_n401), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n403), .A2(new_n404), .ZN(new_n501));
  AOI211_X1 g300(.A(new_n499), .B(new_n500), .C1(new_n395), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n499), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n413), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT40), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n500), .B1(new_n395), .B2(new_n501), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT39), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n413), .A4(new_n503), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n498), .A2(new_n415), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n498), .A2(KEYINPUT82), .A3(new_n415), .A4(new_n510), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n430), .B1(new_n423), .B2(new_n425), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n430), .B2(new_n437), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT38), .B1(new_n517), .B2(KEYINPUT37), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT37), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n441), .B1(new_n440), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n420), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n519), .B2(new_n440), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n522), .A2(KEYINPUT38), .B1(new_n440), .B2(new_n441), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n479), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n515), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n448), .A2(new_n479), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n494), .A2(new_n497), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n258), .B1(new_n492), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT9), .ZN(new_n529));
  INV_X1    g328(.A(G78gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n354), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT89), .ZN(new_n532));
  XOR2_X1   g331(.A(G57gat), .B(G64gat), .Z(new_n533));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n534), .B(new_n529), .C1(new_n354), .C2(new_n530), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G71gat), .B(G78gat), .Z(new_n537));
  OR2_X1    g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT21), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n543), .B(G211gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n542), .B(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(G127gat), .B(G155gat), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n228), .B1(new_n541), .B2(new_n540), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(new_n321), .ZN(new_n550));
  AND2_X1   g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n551), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n556), .B1(new_n553), .B2(new_n554), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n548), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n554), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n555), .B1(new_n560), .B2(new_n552), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n562), .A3(new_n547), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  INV_X1    g364(.A(G85gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(KEYINPUT8), .A2(new_n565), .B1(new_n566), .B2(new_n434), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT7), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n568), .B1(new_n566), .B2(new_n434), .ZN(new_n569));
  NAND3_X1  g368(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n571), .B(new_n572), .Z(new_n573));
  NAND3_X1  g372(.A1(new_n217), .A2(new_n231), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n571), .B(new_n572), .ZN(new_n575));
  AND2_X1   g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n229), .A2(new_n575), .B1(KEYINPUT41), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n576), .A2(KEYINPUT41), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT92), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G190gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G218gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n580), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n540), .A2(new_n573), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT10), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n575), .A2(new_n539), .A3(new_n538), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n575), .A2(KEYINPUT10), .A3(new_n538), .A4(new_n539), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n591), .A2(KEYINPUT93), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT93), .B1(new_n591), .B2(new_n592), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n587), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n588), .A2(new_n590), .ZN(new_n596));
  INV_X1    g395(.A(new_n587), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(new_n303), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n600), .B(G204gat), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n591), .A2(new_n592), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n587), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n598), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n601), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n564), .A2(new_n586), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n528), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n420), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g415(.A(KEYINPUT16), .B(G8gat), .Z(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n498), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT94), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n619), .A2(KEYINPUT42), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(KEYINPUT42), .ZN(new_n621));
  INV_X1    g420(.A(new_n498), .ZN(new_n622));
  OAI21_X1  g421(.A(G8gat), .B1(new_n612), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n623), .A2(KEYINPUT95), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(KEYINPUT95), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n620), .B(new_n621), .C1(new_n624), .C2(new_n625), .ZN(G1325gat));
  INV_X1    g425(.A(G15gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n494), .A2(new_n497), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n612), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n489), .A2(new_n374), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n630), .B1(new_n627), .B2(new_n632), .ZN(G1326gat));
  NOR2_X1   g432(.A1(new_n612), .A2(new_n480), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT43), .B(G22gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(G1327gat));
  AOI21_X1  g435(.A(new_n586), .B1(new_n492), .B2(new_n527), .ZN(new_n637));
  INV_X1    g436(.A(new_n564), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n609), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(new_n258), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n641), .A2(G29gat), .A3(new_n420), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT45), .Z(new_n643));
  NAND2_X1  g442(.A1(new_n492), .A2(new_n527), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(KEYINPUT44), .A3(new_n585), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT96), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n257), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n255), .A2(KEYINPUT96), .A3(new_n256), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n639), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n448), .A2(new_n479), .A3(KEYINPUT97), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n515), .B2(new_n524), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n526), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n653), .A2(new_n494), .A3(new_n497), .A4(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n586), .B1(new_n492), .B2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n645), .B(new_n651), .C1(KEYINPUT44), .C2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(G29gat), .B1(new_n658), .B2(new_n420), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n659), .ZN(G1328gat));
  OR3_X1    g459(.A1(new_n658), .A2(KEYINPUT98), .A3(new_n622), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT98), .B1(new_n658), .B2(new_n622), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(G36gat), .A3(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n641), .A2(G36gat), .A3(new_n622), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT46), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(G1329gat));
  NAND2_X1  g465(.A1(new_n628), .A2(G43gat), .ZN(new_n667));
  INV_X1    g466(.A(new_n631), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n641), .A2(new_n668), .ZN(new_n669));
  OAI22_X1  g468(.A1(new_n658), .A2(new_n667), .B1(new_n669), .B2(G43gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g470(.A(G50gat), .B1(new_n658), .B2(new_n480), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT48), .B1(new_n672), .B2(KEYINPUT99), .ZN(new_n673));
  OR3_X1    g472(.A1(new_n641), .A2(G50gat), .A3(new_n480), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n672), .B(new_n674), .C1(KEYINPUT99), .C2(KEYINPUT48), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(G1331gat));
  NAND4_X1  g477(.A1(new_n650), .A2(new_n564), .A3(new_n586), .A4(new_n608), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT100), .Z(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n492), .B2(new_n656), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n614), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g482(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n681), .A2(new_n498), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT101), .ZN(new_n686));
  NOR2_X1   g485(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n686), .B(new_n688), .ZN(G1333gat));
  AOI21_X1  g488(.A(new_n354), .B1(new_n681), .B2(new_n628), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n681), .A2(new_n631), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n354), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT102), .B(KEYINPUT50), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1334gat));
  NAND2_X1  g493(.A1(new_n681), .A2(new_n479), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G78gat), .ZN(G1335gat));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n492), .A2(new_n656), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n585), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n564), .A2(new_n649), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT51), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT51), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n657), .A2(new_n703), .A3(new_n700), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n702), .A2(new_n614), .A3(new_n608), .A4(new_n704), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n705), .A2(new_n566), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n708), .A2(new_n608), .A3(new_n645), .A4(new_n700), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n566), .A3(new_n420), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n697), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n657), .A2(KEYINPUT44), .ZN(new_n712));
  AOI211_X1 g511(.A(new_n707), .B(new_n586), .C1(new_n492), .C2(new_n527), .ZN(new_n713));
  NOR4_X1   g512(.A1(new_n712), .A2(new_n713), .A3(new_n609), .A4(new_n701), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(G85gat), .A3(new_n614), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n705), .A2(new_n566), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(KEYINPUT103), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n711), .A2(new_n717), .ZN(G1336gat));
  AOI21_X1  g517(.A(new_n434), .B1(new_n714), .B2(new_n498), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n702), .A2(new_n434), .A3(new_n608), .A4(new_n704), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n622), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT52), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G92gat), .B1(new_n709), .B2(new_n622), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n723), .B(new_n724), .C1(new_n622), .C2(new_n720), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n725), .ZN(G1337gat));
  OAI21_X1  g525(.A(G99gat), .B1(new_n709), .B2(new_n629), .ZN(new_n727));
  AND4_X1   g526(.A1(new_n703), .A2(new_n698), .A3(new_n585), .A4(new_n700), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n703), .B1(new_n657), .B2(new_n700), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(G99gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n731), .A3(new_n608), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n727), .B1(new_n732), .B2(new_n668), .ZN(G1338gat));
  OAI21_X1  g532(.A(G106gat), .B1(new_n709), .B2(new_n480), .ZN(new_n734));
  INV_X1    g533(.A(G106gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n730), .A2(new_n735), .A3(new_n479), .A4(new_n608), .ZN(new_n736));
  XNOR2_X1  g535(.A(KEYINPUT104), .B(KEYINPUT53), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n734), .B2(new_n736), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(G1339gat));
  AND4_X1   g539(.A1(new_n564), .A2(new_n650), .A3(new_n586), .A4(new_n609), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n742));
  AOI211_X1 g541(.A(KEYINPUT54), .B(new_n597), .C1(new_n591), .C2(new_n592), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(new_n602), .ZN(new_n744));
  OAI211_X1 g543(.A(KEYINPUT105), .B(new_n601), .C1(new_n605), .C2(KEYINPUT54), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n591), .A2(new_n597), .A3(new_n592), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n595), .A2(KEYINPUT54), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n746), .A2(KEYINPUT55), .A3(new_n748), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n751), .A2(new_n603), .A3(new_n752), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n242), .A2(new_n243), .A3(new_n241), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n235), .B1(new_n232), .B2(new_n234), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n251), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n256), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n753), .A2(new_n585), .A3(new_n757), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n649), .A2(new_n753), .B1(new_n608), .B2(new_n757), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(new_n585), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n741), .B1(new_n760), .B2(new_n638), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n479), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n762), .A2(new_n614), .A3(new_n622), .A4(new_n631), .ZN(new_n763));
  OAI21_X1  g562(.A(G113gat), .B1(new_n763), .B2(new_n258), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n746), .A2(KEYINPUT55), .A3(new_n748), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT55), .B1(new_n746), .B2(new_n748), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n255), .A2(KEYINPUT96), .A3(new_n256), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT96), .B1(new_n255), .B2(new_n256), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n767), .B(new_n603), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n757), .A2(new_n608), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n585), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n758), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n638), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n650), .A2(new_n564), .A3(new_n586), .A4(new_n609), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n614), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n374), .A2(new_n452), .A3(new_n480), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n777), .A2(new_n498), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n650), .A2(new_n261), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n764), .B1(new_n780), .B2(new_n781), .ZN(G1340gat));
  NAND3_X1  g581(.A1(new_n779), .A2(new_n262), .A3(new_n608), .ZN(new_n783));
  OAI21_X1  g582(.A(G120gat), .B1(new_n763), .B2(new_n609), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT106), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(KEYINPUT107), .B(new_n783), .C1(new_n786), .C2(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1341gat));
  AOI21_X1  g591(.A(G127gat), .B1(new_n779), .B2(new_n564), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n763), .A2(new_n638), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(G127gat), .B2(new_n794), .ZN(G1342gat));
  NOR3_X1   g594(.A1(new_n780), .A2(G134gat), .A3(new_n586), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT56), .ZN(new_n797));
  OAI21_X1  g596(.A(G134gat), .B1(new_n763), .B2(new_n586), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1343gat));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n761), .B2(new_n480), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n257), .A2(new_n751), .A3(new_n603), .A4(new_n752), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n771), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n586), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n758), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n638), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n775), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(KEYINPUT108), .A3(KEYINPUT57), .A4(new_n479), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n564), .B1(new_n804), .B2(new_n758), .ZN(new_n809));
  OAI211_X1 g608(.A(KEYINPUT57), .B(new_n479), .C1(new_n809), .C2(new_n741), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT108), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n801), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n628), .A2(new_n420), .A3(new_n498), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n257), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT58), .B1(new_n817), .B2(G141gat), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n629), .B1(new_n777), .B2(KEYINPUT109), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n420), .B1(new_n774), .B2(new_n775), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT109), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n622), .B(new_n479), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(G141gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n824), .A3(new_n257), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(KEYINPUT110), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(KEYINPUT110), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n818), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(G141gat), .B1(new_n815), .B2(new_n650), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n825), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT58), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n831), .ZN(G1344gat));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n833), .A3(new_n608), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n611), .A2(new_n258), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n806), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n800), .A3(new_n479), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n761), .A2(new_n480), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n608), .B(new_n837), .C1(new_n838), .C2(new_n800), .ZN(new_n839));
  INV_X1    g638(.A(new_n814), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT59), .B(G148gat), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n833), .B1(new_n823), .B2(new_n608), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n834), .B(new_n841), .C1(G148gat), .C2(new_n842), .ZN(G1345gat));
  NOR3_X1   g642(.A1(new_n815), .A2(new_n384), .A3(new_n638), .ZN(new_n844));
  AOI21_X1  g643(.A(G155gat), .B1(new_n823), .B2(new_n564), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(G1346gat));
  INV_X1    g645(.A(new_n822), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n628), .B1(new_n820), .B2(new_n821), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n847), .A2(new_n385), .A3(new_n585), .A4(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT111), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n823), .A2(KEYINPUT111), .A3(new_n385), .A4(new_n585), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n813), .A2(new_n585), .A3(new_n814), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT112), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n813), .A2(new_n856), .A3(new_n585), .A4(new_n814), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(G162gat), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n853), .A2(new_n858), .A3(KEYINPUT113), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1347gat));
  NOR2_X1   g662(.A1(new_n778), .A2(new_n622), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n614), .B1(new_n864), .B2(KEYINPUT114), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n865), .B(new_n776), .C1(KEYINPUT114), .C2(new_n864), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(KEYINPUT115), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(KEYINPUT115), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n302), .A3(new_n649), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n622), .A2(new_n614), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n762), .A2(new_n631), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G169gat), .B1(new_n873), .B2(new_n258), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(KEYINPUT116), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(KEYINPUT116), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(G1348gat));
  NOR3_X1   g676(.A1(new_n873), .A2(new_n303), .A3(new_n609), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n870), .A2(new_n608), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n303), .ZN(G1349gat));
  OR3_X1    g679(.A1(new_n866), .A2(new_n283), .A3(new_n638), .ZN(new_n881));
  OAI21_X1  g680(.A(G183gat), .B1(new_n873), .B2(new_n638), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g682(.A(KEYINPUT117), .B(KEYINPUT60), .Z(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT118), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n887), .B1(new_n883), .B2(KEYINPUT60), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n886), .B1(new_n888), .B2(new_n885), .ZN(G1350gat));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n586), .A2(G190gat), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n869), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n762), .A2(new_n631), .A3(new_n585), .A4(new_n872), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n894), .A2(new_n895), .A3(G190gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n894), .B2(G190gat), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n890), .B1(new_n893), .B2(new_n898), .ZN(new_n899));
  OAI221_X1 g698(.A(KEYINPUT119), .B1(new_n896), .B2(new_n897), .C1(new_n869), .C2(new_n892), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1351gat));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902));
  AOI211_X1 g701(.A(KEYINPUT57), .B(new_n480), .C1(new_n835), .C2(new_n806), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n800), .B1(new_n776), .B2(new_n479), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g704(.A(KEYINPUT120), .B(new_n837), .C1(new_n838), .C2(new_n800), .ZN(new_n906));
  INV_X1    g705(.A(new_n872), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT121), .B1(new_n628), .B2(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n628), .A2(new_n614), .A3(new_n622), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n905), .A2(new_n906), .A3(new_n908), .A4(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G197gat), .B1(new_n912), .B2(new_n258), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n838), .A2(new_n909), .ZN(new_n915));
  OR3_X1    g714(.A1(new_n915), .A2(G197gat), .A3(new_n650), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n914), .B1(new_n913), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(G1352gat));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n920));
  OR3_X1    g719(.A1(new_n912), .A2(new_n920), .A3(new_n609), .ZN(new_n921));
  XOR2_X1   g720(.A(KEYINPUT123), .B(G204gat), .Z(new_n922));
  OAI21_X1  g721(.A(new_n920), .B1(new_n912), .B2(new_n609), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n915), .B1(new_n925), .B2(KEYINPUT62), .ZN(new_n926));
  INV_X1    g725(.A(new_n922), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n608), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n925), .A2(KEYINPUT62), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n924), .A2(new_n930), .ZN(G1353gat));
  NAND2_X1  g730(.A1(new_n911), .A2(new_n908), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n564), .B(new_n837), .C1(new_n838), .C2(new_n800), .ZN(new_n933));
  OAI21_X1  g732(.A(G211gat), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(KEYINPUT126), .A3(new_n937), .ZN(new_n938));
  OR3_X1    g737(.A1(new_n915), .A2(G211gat), .A3(new_n638), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n940), .A3(new_n935), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n912), .B2(new_n586), .ZN(new_n943));
  OR3_X1    g742(.A1(new_n915), .A2(G218gat), .A3(new_n586), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n943), .A2(KEYINPUT127), .A3(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1355gat));
endmodule


