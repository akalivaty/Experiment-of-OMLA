

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577;

  XNOR2_X1 U320 ( .A(n377), .B(n376), .ZN(n549) );
  XNOR2_X1 U321 ( .A(n308), .B(n307), .ZN(n526) );
  XNOR2_X1 U322 ( .A(n430), .B(n375), .ZN(n376) );
  XOR2_X1 U323 ( .A(n458), .B(KEYINPUT28), .Z(n524) );
  XNOR2_X1 U324 ( .A(n440), .B(G183GAT), .ZN(n441) );
  XNOR2_X1 U325 ( .A(n442), .B(n441), .ZN(G1350GAT) );
  XOR2_X1 U326 ( .A(KEYINPUT79), .B(KEYINPUT82), .Z(n289) );
  XNOR2_X1 U327 ( .A(KEYINPUT20), .B(G120GAT), .ZN(n288) );
  XNOR2_X1 U328 ( .A(n289), .B(n288), .ZN(n308) );
  XOR2_X1 U329 ( .A(G99GAT), .B(G134GAT), .Z(n291) );
  XNOR2_X1 U330 ( .A(G43GAT), .B(G190GAT), .ZN(n290) );
  XNOR2_X1 U331 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U332 ( .A(KEYINPUT78), .B(G71GAT), .Z(n293) );
  XNOR2_X1 U333 ( .A(G15GAT), .B(KEYINPUT81), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U335 ( .A(n295), .B(n294), .Z(n306) );
  XNOR2_X1 U336 ( .A(KEYINPUT80), .B(KEYINPUT18), .ZN(n296) );
  XNOR2_X1 U337 ( .A(n296), .B(KEYINPUT19), .ZN(n297) );
  XOR2_X1 U338 ( .A(n297), .B(KEYINPUT17), .Z(n299) );
  XNOR2_X1 U339 ( .A(G169GAT), .B(G183GAT), .ZN(n298) );
  XNOR2_X1 U340 ( .A(n299), .B(n298), .ZN(n431) );
  XOR2_X1 U341 ( .A(G127GAT), .B(KEYINPUT77), .Z(n301) );
  XNOR2_X1 U342 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n300) );
  XNOR2_X1 U343 ( .A(n301), .B(n300), .ZN(n331) );
  XOR2_X1 U344 ( .A(n331), .B(G176GAT), .Z(n303) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U347 ( .A(n431), .B(n304), .ZN(n305) );
  XNOR2_X1 U348 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U349 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n310) );
  XNOR2_X1 U350 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n309) );
  XNOR2_X1 U351 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U352 ( .A(G141GAT), .B(n311), .ZN(n340) );
  XOR2_X1 U353 ( .A(G148GAT), .B(KEYINPUT85), .Z(n313) );
  XNOR2_X1 U354 ( .A(KEYINPUT23), .B(KEYINPUT83), .ZN(n312) );
  XNOR2_X1 U355 ( .A(n313), .B(n312), .ZN(n324) );
  XOR2_X1 U356 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n315) );
  XOR2_X1 U357 ( .A(G50GAT), .B(G162GAT), .Z(n364) );
  XOR2_X1 U358 ( .A(G204GAT), .B(G78GAT), .Z(n396) );
  XNOR2_X1 U359 ( .A(n364), .B(n396), .ZN(n314) );
  XNOR2_X1 U360 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U361 ( .A(n316), .B(G106GAT), .Z(n322) );
  XNOR2_X1 U362 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n317) );
  XNOR2_X1 U363 ( .A(n317), .B(G211GAT), .ZN(n422) );
  XOR2_X1 U364 ( .A(n422), .B(G22GAT), .Z(n319) );
  NAND2_X1 U365 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U367 ( .A(n320), .B(G218GAT), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U369 ( .A(n324), .B(n323), .Z(n325) );
  XNOR2_X1 U370 ( .A(n340), .B(n325), .ZN(n458) );
  XNOR2_X1 U371 ( .A(G120GAT), .B(G148GAT), .ZN(n326) );
  XNOR2_X1 U372 ( .A(n326), .B(G57GAT), .ZN(n399) );
  XOR2_X1 U373 ( .A(KEYINPUT86), .B(n399), .Z(n328) );
  XNOR2_X1 U374 ( .A(G162GAT), .B(KEYINPUT88), .ZN(n327) );
  XNOR2_X1 U375 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U376 ( .A(n329), .B(KEYINPUT5), .Z(n333) );
  XNOR2_X1 U377 ( .A(G29GAT), .B(G134GAT), .ZN(n330) );
  XNOR2_X1 U378 ( .A(n330), .B(G85GAT), .ZN(n373) );
  XNOR2_X1 U379 ( .A(n331), .B(n373), .ZN(n332) );
  XNOR2_X1 U380 ( .A(n333), .B(n332), .ZN(n345) );
  XOR2_X1 U381 ( .A(KEYINPUT87), .B(KEYINPUT1), .Z(n335) );
  XNOR2_X1 U382 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U384 ( .A(KEYINPUT89), .B(n336), .Z(n338) );
  NAND2_X1 U385 ( .A1(G225GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U386 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U387 ( .A(n339), .B(KEYINPUT4), .Z(n343) );
  INV_X1 U388 ( .A(n340), .ZN(n341) );
  XNOR2_X1 U389 ( .A(G1GAT), .B(n341), .ZN(n342) );
  XNOR2_X1 U390 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U391 ( .A(n345), .B(n344), .Z(n456) );
  XNOR2_X1 U392 ( .A(KEYINPUT91), .B(n456), .ZN(n513) );
  INV_X1 U393 ( .A(KEYINPUT54), .ZN(n435) );
  XOR2_X1 U394 ( .A(G36GAT), .B(G29GAT), .Z(n347) );
  NAND2_X1 U395 ( .A1(G229GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U396 ( .A(n347), .B(n346), .ZN(n360) );
  XOR2_X1 U397 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n349) );
  XNOR2_X1 U398 ( .A(G141GAT), .B(KEYINPUT29), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U400 ( .A(G197GAT), .B(G113GAT), .Z(n351) );
  XNOR2_X1 U401 ( .A(G169GAT), .B(G50GAT), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U403 ( .A(n353), .B(n352), .Z(n358) );
  XNOR2_X1 U404 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n354) );
  XNOR2_X1 U405 ( .A(n354), .B(KEYINPUT7), .ZN(n374) );
  XOR2_X1 U406 ( .A(G8GAT), .B(G1GAT), .Z(n356) );
  XNOR2_X1 U407 ( .A(G15GAT), .B(G22GAT), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n356), .B(n355), .ZN(n378) );
  XNOR2_X1 U409 ( .A(n374), .B(n378), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U411 ( .A(n360), .B(n359), .ZN(n561) );
  XOR2_X1 U412 ( .A(KEYINPUT72), .B(KEYINPUT9), .Z(n362) );
  XNOR2_X1 U413 ( .A(KEYINPUT10), .B(KEYINPUT11), .ZN(n361) );
  XOR2_X1 U414 ( .A(n362), .B(n361), .Z(n367) );
  XOR2_X1 U415 ( .A(KEYINPUT73), .B(KEYINPUT65), .Z(n363) );
  XNOR2_X1 U416 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U417 ( .A(G99GAT), .B(G106GAT), .Z(n395) );
  XNOR2_X1 U418 ( .A(n365), .B(n395), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n367), .B(n366), .ZN(n369) );
  NAND2_X1 U420 ( .A1(G232GAT), .A2(G233GAT), .ZN(n368) );
  XOR2_X1 U421 ( .A(n369), .B(n368), .Z(n377) );
  XOR2_X1 U422 ( .A(G92GAT), .B(KEYINPUT74), .Z(n371) );
  XNOR2_X1 U423 ( .A(G190GAT), .B(G218GAT), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U425 ( .A(G36GAT), .B(n372), .Z(n430) );
  XNOR2_X1 U426 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U427 ( .A(KEYINPUT75), .B(n549), .Z(n534) );
  XNOR2_X1 U428 ( .A(n534), .B(KEYINPUT36), .ZN(n573) );
  XOR2_X1 U429 ( .A(KEYINPUT15), .B(n378), .Z(n380) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U431 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U432 ( .A(G71GAT), .B(KEYINPUT13), .Z(n394) );
  XOR2_X1 U433 ( .A(n381), .B(n394), .Z(n383) );
  XNOR2_X1 U434 ( .A(G183GAT), .B(G127GAT), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n383), .B(n382), .ZN(n391) );
  XOR2_X1 U436 ( .A(G57GAT), .B(G78GAT), .Z(n385) );
  XNOR2_X1 U437 ( .A(G155GAT), .B(G211GAT), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U439 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n387) );
  XNOR2_X1 U440 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U442 ( .A(n389), .B(n388), .Z(n390) );
  XNOR2_X1 U443 ( .A(n391), .B(n390), .ZN(n571) );
  NAND2_X1 U444 ( .A1(n573), .A2(n571), .ZN(n393) );
  XNOR2_X1 U445 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n393), .B(n392), .ZN(n412) );
  XOR2_X1 U447 ( .A(G176GAT), .B(G64GAT), .Z(n423) );
  XOR2_X1 U448 ( .A(n423), .B(n394), .Z(n398) );
  XNOR2_X1 U449 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n398), .B(n397), .ZN(n403) );
  XOR2_X1 U451 ( .A(n399), .B(KEYINPUT68), .Z(n401) );
  NAND2_X1 U452 ( .A1(G230GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U453 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U454 ( .A(n403), .B(n402), .Z(n411) );
  XOR2_X1 U455 ( .A(KEYINPUT31), .B(KEYINPUT69), .Z(n405) );
  XNOR2_X1 U456 ( .A(G85GAT), .B(G92GAT), .ZN(n404) );
  XNOR2_X1 U457 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U458 ( .A(KEYINPUT67), .B(KEYINPUT33), .Z(n407) );
  XNOR2_X1 U459 ( .A(KEYINPUT32), .B(KEYINPUT70), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U461 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U462 ( .A(n411), .B(n410), .ZN(n566) );
  NAND2_X1 U463 ( .A1(n412), .A2(n566), .ZN(n413) );
  OR2_X1 U464 ( .A1(n561), .A2(n413), .ZN(n420) );
  XOR2_X1 U465 ( .A(n566), .B(KEYINPUT41), .Z(n499) );
  INV_X1 U466 ( .A(n499), .ZN(n553) );
  NAND2_X1 U467 ( .A1(n561), .A2(n553), .ZN(n414) );
  XNOR2_X1 U468 ( .A(KEYINPUT46), .B(n414), .ZN(n415) );
  INV_X1 U469 ( .A(n571), .ZN(n463) );
  NAND2_X1 U470 ( .A1(n415), .A2(n463), .ZN(n416) );
  NOR2_X1 U471 ( .A1(n549), .A2(n416), .ZN(n418) );
  XNOR2_X1 U472 ( .A(KEYINPUT112), .B(KEYINPUT47), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n419) );
  NAND2_X1 U474 ( .A1(n420), .A2(n419), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n421), .B(KEYINPUT48), .ZN(n521) );
  XOR2_X1 U476 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U477 ( .A1(G226GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U479 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n427) );
  XNOR2_X1 U480 ( .A(G8GAT), .B(G204GAT), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U482 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U483 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U484 ( .A(n433), .B(n432), .ZN(n452) );
  NAND2_X1 U485 ( .A1(n521), .A2(n452), .ZN(n434) );
  XNOR2_X1 U486 ( .A(n435), .B(n434), .ZN(n436) );
  NAND2_X1 U487 ( .A1(n513), .A2(n436), .ZN(n437) );
  XNOR2_X1 U488 ( .A(n437), .B(KEYINPUT64), .ZN(n560) );
  NOR2_X1 U489 ( .A1(n458), .A2(n560), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n438), .B(KEYINPUT55), .ZN(n439) );
  NOR2_X2 U491 ( .A1(n526), .A2(n439), .ZN(n554) );
  NAND2_X1 U492 ( .A1(n554), .A2(n571), .ZN(n442) );
  XOR2_X1 U493 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n440) );
  INV_X1 U494 ( .A(G190GAT), .ZN(n446) );
  XOR2_X1 U495 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n444) );
  NAND2_X1 U496 ( .A1(n554), .A2(n534), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(G1351GAT) );
  NAND2_X1 U499 ( .A1(n561), .A2(n566), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n447), .B(KEYINPUT71), .ZN(n482) );
  INV_X1 U501 ( .A(n452), .ZN(n515) );
  NOR2_X1 U502 ( .A1(n526), .A2(n515), .ZN(n448) );
  NOR2_X1 U503 ( .A1(n458), .A2(n448), .ZN(n449) );
  XOR2_X1 U504 ( .A(n449), .B(KEYINPUT25), .Z(n450) );
  XNOR2_X1 U505 ( .A(KEYINPUT94), .B(n450), .ZN(n454) );
  NAND2_X1 U506 ( .A1(n526), .A2(n458), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n451), .B(KEYINPUT26), .ZN(n559) );
  XOR2_X1 U508 ( .A(n452), .B(KEYINPUT27), .Z(n457) );
  NOR2_X1 U509 ( .A1(n559), .A2(n457), .ZN(n453) );
  NOR2_X1 U510 ( .A1(n454), .A2(n453), .ZN(n455) );
  NOR2_X1 U511 ( .A1(n456), .A2(n455), .ZN(n462) );
  INV_X1 U512 ( .A(n526), .ZN(n460) );
  NOR2_X1 U513 ( .A1(n457), .A2(n513), .ZN(n522) );
  NAND2_X1 U514 ( .A1(n522), .A2(n524), .ZN(n459) );
  NOR2_X1 U515 ( .A1(n460), .A2(n459), .ZN(n461) );
  NOR2_X1 U516 ( .A1(n462), .A2(n461), .ZN(n478) );
  NOR2_X1 U517 ( .A1(n534), .A2(n463), .ZN(n464) );
  XOR2_X1 U518 ( .A(KEYINPUT16), .B(n464), .Z(n465) );
  NOR2_X1 U519 ( .A1(n478), .A2(n465), .ZN(n500) );
  NAND2_X1 U520 ( .A1(n482), .A2(n500), .ZN(n466) );
  XOR2_X1 U521 ( .A(KEYINPUT95), .B(n466), .Z(n475) );
  NOR2_X1 U522 ( .A1(n513), .A2(n475), .ZN(n468) );
  XNOR2_X1 U523 ( .A(KEYINPUT34), .B(KEYINPUT96), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n468), .B(n467), .ZN(n469) );
  XOR2_X1 U525 ( .A(G1GAT), .B(n469), .Z(G1324GAT) );
  NOR2_X1 U526 ( .A1(n515), .A2(n475), .ZN(n470) );
  XOR2_X1 U527 ( .A(G8GAT), .B(n470), .Z(G1325GAT) );
  NOR2_X1 U528 ( .A1(n475), .A2(n526), .ZN(n474) );
  XOR2_X1 U529 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n472) );
  XNOR2_X1 U530 ( .A(G15GAT), .B(KEYINPUT98), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(G1326GAT) );
  NOR2_X1 U533 ( .A1(n524), .A2(n475), .ZN(n477) );
  XNOR2_X1 U534 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(G1327GAT) );
  XNOR2_X1 U536 ( .A(KEYINPUT37), .B(KEYINPUT100), .ZN(n481) );
  NOR2_X1 U537 ( .A1(n478), .A2(n571), .ZN(n479) );
  NAND2_X1 U538 ( .A1(n479), .A2(n573), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(n511) );
  NAND2_X1 U540 ( .A1(n511), .A2(n482), .ZN(n485) );
  XOR2_X1 U541 ( .A(KEYINPUT38), .B(KEYINPUT101), .Z(n483) );
  XNOR2_X1 U542 ( .A(KEYINPUT102), .B(n483), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(n493) );
  NOR2_X1 U544 ( .A1(n493), .A2(n513), .ZN(n488) );
  XOR2_X1 U545 ( .A(G29GAT), .B(KEYINPUT39), .Z(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT103), .B(n486), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  NOR2_X1 U548 ( .A1(n515), .A2(n493), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT104), .B(n489), .Z(n490) );
  XNOR2_X1 U550 ( .A(G36GAT), .B(n490), .ZN(G1329GAT) );
  NOR2_X1 U551 ( .A1(n526), .A2(n493), .ZN(n491) );
  XOR2_X1 U552 ( .A(KEYINPUT40), .B(n491), .Z(n492) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(n492), .ZN(G1330GAT) );
  NOR2_X1 U554 ( .A1(n524), .A2(n493), .ZN(n495) );
  XNOR2_X1 U555 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U557 ( .A(G50GAT), .B(n496), .ZN(G1331GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n498) );
  XNOR2_X1 U559 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n502) );
  NOR2_X1 U561 ( .A1(n499), .A2(n561), .ZN(n510) );
  NAND2_X1 U562 ( .A1(n510), .A2(n500), .ZN(n505) );
  NOR2_X1 U563 ( .A1(n513), .A2(n505), .ZN(n501) );
  XOR2_X1 U564 ( .A(n502), .B(n501), .Z(G1332GAT) );
  NOR2_X1 U565 ( .A1(n515), .A2(n505), .ZN(n503) );
  XOR2_X1 U566 ( .A(G64GAT), .B(n503), .Z(G1333GAT) );
  NOR2_X1 U567 ( .A1(n526), .A2(n505), .ZN(n504) );
  XOR2_X1 U568 ( .A(G71GAT), .B(n504), .Z(G1334GAT) );
  NOR2_X1 U569 ( .A1(n505), .A2(n524), .ZN(n509) );
  XOR2_X1 U570 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n507) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT110), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n510), .ZN(n512) );
  XOR2_X1 U575 ( .A(KEYINPUT111), .B(n512), .Z(n518) );
  NOR2_X1 U576 ( .A1(n513), .A2(n518), .ZN(n514) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n514), .Z(G1336GAT) );
  NOR2_X1 U578 ( .A1(n515), .A2(n518), .ZN(n516) );
  XOR2_X1 U579 ( .A(G92GAT), .B(n516), .Z(G1337GAT) );
  NOR2_X1 U580 ( .A1(n526), .A2(n518), .ZN(n517) );
  XOR2_X1 U581 ( .A(G99GAT), .B(n517), .Z(G1338GAT) );
  NOR2_X1 U582 ( .A1(n524), .A2(n518), .ZN(n519) );
  XOR2_X1 U583 ( .A(KEYINPUT44), .B(n519), .Z(n520) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  NAND2_X1 U585 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U586 ( .A(KEYINPUT114), .B(n523), .Z(n539) );
  NAND2_X1 U587 ( .A1(n524), .A2(n539), .ZN(n525) );
  NOR2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n535), .A2(n561), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .Z(n529) );
  NAND2_X1 U592 ( .A1(n535), .A2(n553), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(G1341GAT) );
  NAND2_X1 U594 ( .A1(n571), .A2(n535), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(KEYINPUT50), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n533) );
  XNOR2_X1 U598 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(KEYINPUT115), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  INV_X1 U603 ( .A(n539), .ZN(n540) );
  NOR2_X1 U604 ( .A1(n559), .A2(n540), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n550), .A2(n561), .ZN(n541) );
  XNOR2_X1 U606 ( .A(KEYINPUT118), .B(n541), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n544) );
  NAND2_X1 U609 ( .A1(n550), .A2(n553), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n546) );
  XOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT52), .Z(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U613 ( .A1(n571), .A2(n550), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(KEYINPUT120), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G155GAT), .B(n548), .ZN(G1346GAT) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U618 ( .A1(n561), .A2(n554), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n556) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n558) );
  XOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT56), .Z(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  XOR2_X1 U625 ( .A(G197GAT), .B(KEYINPUT60), .Z(n563) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n574) );
  NAND2_X1 U627 ( .A1(n574), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U629 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1352GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n569) );
  INV_X1 U632 ( .A(n566), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n574), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(n570), .ZN(G1353GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n574), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n576) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(n577), .ZN(G1355GAT) );
endmodule

