

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n369, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n390, n392, n393, n394, n395, n397, n398, n400, n401,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n537,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792;

  INV_X1 U375 ( .A(n574), .ZN(n358) );
  INV_X1 U376 ( .A(n569), .ZN(n361) );
  INV_X1 U377 ( .A(n664), .ZN(n354) );
  NOR2_X1 U378 ( .A1(n790), .A2(n791), .ZN(n617) );
  BUF_X1 U379 ( .A(n747), .Z(n364) );
  INV_X1 U380 ( .A(n537), .ZN(n366) );
  XNOR2_X1 U381 ( .A(n604), .B(KEYINPUT1), .ZN(n747) );
  XNOR2_X1 U382 ( .A(n363), .B(n782), .ZN(n511) );
  XNOR2_X1 U383 ( .A(n508), .B(KEYINPUT72), .ZN(n363) );
  XNOR2_X1 U384 ( .A(n437), .B(n663), .ZN(n418) );
  XNOR2_X1 U385 ( .A(G107), .B(G104), .ZN(n417) );
  XOR2_X1 U386 ( .A(KEYINPUT5), .B(KEYINPUT100), .Z(n494) );
  XNOR2_X1 U387 ( .A(n352), .B(KEYINPUT84), .ZN(n390) );
  NAND2_X1 U388 ( .A1(n356), .A2(n388), .ZN(n352) );
  XNOR2_X1 U389 ( .A(n357), .B(n574), .ZN(n380) );
  NAND2_X1 U390 ( .A1(n400), .A2(n403), .ZN(n357) );
  NAND2_X1 U391 ( .A1(n353), .A2(KEYINPUT44), .ZN(n556) );
  NAND2_X1 U392 ( .A1(n355), .A2(n354), .ZN(n353) );
  INV_X1 U393 ( .A(n665), .ZN(n355) );
  NAND2_X1 U394 ( .A1(n394), .A2(n393), .ZN(n356) );
  XNOR2_X2 U395 ( .A(n567), .B(KEYINPUT35), .ZN(n666) );
  XNOR2_X1 U396 ( .A(n359), .B(n358), .ZN(n367) );
  NAND2_X1 U397 ( .A1(n400), .A2(n403), .ZN(n359) );
  NAND2_X2 U398 ( .A1(n360), .A2(n401), .ZN(n400) );
  XNOR2_X2 U399 ( .A(n572), .B(n571), .ZN(n360) );
  AND2_X2 U400 ( .A1(n406), .A2(n377), .ZN(n395) );
  OR2_X2 U401 ( .A1(n666), .A2(n361), .ZN(n572) );
  OR2_X2 U402 ( .A1(n669), .A2(G902), .ZN(n504) );
  XNOR2_X2 U403 ( .A(n362), .B(n378), .ZN(n631) );
  NAND2_X2 U404 ( .A1(n611), .A2(n424), .ZN(n362) );
  XNOR2_X2 U405 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X2 U406 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X2 U407 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U408 ( .A(n543), .B(n366), .ZN(n560) );
  OR2_X2 U409 ( .A1(n685), .A2(G902), .ZN(n428) );
  XNOR2_X2 U410 ( .A(n621), .B(KEYINPUT19), .ZN(n607) );
  NAND2_X2 U411 ( .A1(n425), .A2(n430), .ZN(n456) );
  XNOR2_X1 U412 ( .A(n365), .B(n509), .ZN(n690) );
  XNOR2_X1 U413 ( .A(n781), .B(n446), .ZN(n365) );
  NOR2_X2 U414 ( .A1(n607), .A2(n462), .ZN(n463) );
  XNOR2_X2 U415 ( .A(n463), .B(KEYINPUT0), .ZN(n543) );
  NAND2_X1 U416 ( .A1(G953), .A2(G902), .ZN(n580) );
  INV_X1 U417 ( .A(G237), .ZN(n448) );
  XNOR2_X1 U418 ( .A(G131), .B(G101), .ZN(n496) );
  AND2_X1 U419 ( .A1(n465), .A2(G224), .ZN(n442) );
  XNOR2_X1 U420 ( .A(G116), .B(G119), .ZN(n413) );
  XNOR2_X1 U421 ( .A(G116), .B(G107), .ZN(n470) );
  INV_X2 U422 ( .A(G953), .ZN(n465) );
  BUF_X1 U423 ( .A(G104), .Z(n661) );
  XNOR2_X1 U424 ( .A(n384), .B(KEYINPUT105), .ZN(n712) );
  NAND2_X1 U425 ( .A1(n748), .A2(n604), .ZN(n588) );
  INV_X1 U426 ( .A(G110), .ZN(n663) );
  OR2_X1 U427 ( .A1(n642), .A2(n775), .ZN(n727) );
  XNOR2_X1 U428 ( .A(n548), .B(n547), .ZN(n715) );
  INV_X1 U429 ( .A(n576), .ZN(n737) );
  OR2_X1 U430 ( .A1(n712), .A2(n714), .ZN(n576) );
  XNOR2_X1 U431 ( .A(n559), .B(n558), .ZN(n735) );
  OR2_X1 U432 ( .A1(n563), .A2(n564), .ZN(n384) );
  XNOR2_X1 U433 ( .A(n541), .B(KEYINPUT69), .ZN(n748) );
  NOR2_X1 U434 ( .A1(n577), .A2(n736), .ZN(n579) );
  XNOR2_X1 U435 ( .A(n522), .B(n521), .ZN(n675) );
  XNOR2_X1 U436 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U437 ( .A(n490), .B(n427), .ZN(n653) );
  XNOR2_X1 U438 ( .A(n464), .B(G134), .ZN(n490) );
  XNOR2_X1 U439 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n574) );
  XNOR2_X1 U440 ( .A(KEYINPUT73), .B(KEYINPUT34), .ZN(n561) );
  XNOR2_X2 U441 ( .A(G146), .B(G125), .ZN(n478) );
  XNOR2_X2 U442 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n489) );
  BUF_X1 U443 ( .A(n781), .Z(n369) );
  XNOR2_X1 U444 ( .A(n491), .B(n440), .ZN(n781) );
  XNOR2_X1 U445 ( .A(n414), .B(n413), .ZN(n491) );
  XNOR2_X1 U446 ( .A(n438), .B(n415), .ZN(n414) );
  XNOR2_X1 U447 ( .A(n782), .B(KEYINPUT72), .ZN(n509) );
  NOR2_X1 U448 ( .A1(G953), .A2(G237), .ZN(n492) );
  AND2_X1 U449 ( .A1(n747), .A2(n748), .ZN(n557) );
  XNOR2_X1 U450 ( .A(n474), .B(KEYINPUT104), .ZN(n387) );
  XNOR2_X1 U451 ( .A(G113), .B(G122), .ZN(n474) );
  XOR2_X1 U452 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n475) );
  XNOR2_X1 U453 ( .A(G902), .B(KEYINPUT15), .ZN(n641) );
  INV_X1 U454 ( .A(KEYINPUT10), .ZN(n477) );
  INV_X1 U455 ( .A(KEYINPUT40), .ZN(n612) );
  XNOR2_X1 U456 ( .A(n598), .B(n597), .ZN(n609) );
  INV_X1 U457 ( .A(KEYINPUT68), .ZN(n571) );
  XNOR2_X1 U458 ( .A(n573), .B(n416), .ZN(n401) );
  INV_X1 U459 ( .A(KEYINPUT89), .ZN(n416) );
  NOR2_X1 U460 ( .A1(n409), .A2(n408), .ZN(n407) );
  INV_X1 U461 ( .A(KEYINPUT76), .ZN(n408) );
  NAND2_X1 U462 ( .A1(n450), .A2(n575), .ZN(n433) );
  NOR2_X1 U463 ( .A1(n789), .A2(n412), .ZN(n411) );
  INV_X1 U464 ( .A(n721), .ZN(n412) );
  XNOR2_X1 U465 ( .A(n489), .B(G137), .ZN(n427) );
  AND2_X1 U466 ( .A1(n392), .A2(n379), .ZN(n388) );
  XNOR2_X1 U467 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n441) );
  NAND2_X1 U468 ( .A1(G237), .A2(G234), .ZN(n460) );
  NAND2_X1 U469 ( .A1(n432), .A2(n641), .ZN(n431) );
  INV_X1 U470 ( .A(n450), .ZN(n432) );
  INV_X1 U471 ( .A(G902), .ZN(n523) );
  XNOR2_X1 U472 ( .A(KEYINPUT16), .B(G122), .ZN(n439) );
  XNOR2_X1 U473 ( .A(n422), .B(n421), .ZN(n518) );
  INV_X1 U474 ( .A(KEYINPUT8), .ZN(n421) );
  NAND2_X1 U475 ( .A1(n465), .A2(G234), .ZN(n422) );
  XNOR2_X1 U476 ( .A(G128), .B(G137), .ZN(n512) );
  XNOR2_X1 U477 ( .A(G119), .B(KEYINPUT23), .ZN(n514) );
  INV_X1 U478 ( .A(KEYINPUT9), .ZN(n466) );
  XOR2_X2 U479 ( .A(G122), .B(KEYINPUT7), .Z(n467) );
  XNOR2_X1 U480 ( .A(n386), .B(n385), .ZN(n479) );
  XNOR2_X1 U481 ( .A(n475), .B(n373), .ZN(n385) );
  XNOR2_X1 U482 ( .A(n476), .B(n387), .ZN(n386) );
  XOR2_X1 U483 ( .A(G131), .B(G140), .Z(n507) );
  INV_X1 U484 ( .A(KEYINPUT98), .ZN(n537) );
  NAND2_X1 U485 ( .A1(n648), .A2(G953), .ZN(n696) );
  INV_X1 U486 ( .A(KEYINPUT122), .ZN(n771) );
  OR2_X1 U487 ( .A1(n632), .A2(KEYINPUT76), .ZN(n371) );
  AND2_X1 U488 ( .A1(n632), .A2(n411), .ZN(n372) );
  AND2_X1 U489 ( .A1(G214), .A2(n492), .ZN(n373) );
  XOR2_X1 U490 ( .A(n610), .B(KEYINPUT82), .Z(n374) );
  AND2_X1 U491 ( .A1(n430), .A2(n433), .ZN(n375) );
  OR2_X1 U492 ( .A1(n736), .A2(n429), .ZN(n376) );
  OR2_X1 U493 ( .A1(n411), .A2(KEYINPUT76), .ZN(n377) );
  XOR2_X1 U494 ( .A(KEYINPUT87), .B(KEYINPUT39), .Z(n378) );
  OR2_X1 U495 ( .A1(n575), .A2(KEYINPUT85), .ZN(n379) );
  BUF_X1 U496 ( .A(n426), .Z(n381) );
  NAND2_X1 U497 ( .A1(n382), .A2(KEYINPUT48), .ZN(n630) );
  INV_X1 U498 ( .A(n628), .ZN(n382) );
  NAND2_X1 U499 ( .A1(n383), .A2(n435), .ZN(n628) );
  AND2_X1 U500 ( .A1(n374), .A2(n420), .ZN(n383) );
  NAND2_X1 U501 ( .A1(n390), .A2(n436), .ZN(n643) );
  NAND2_X1 U502 ( .A1(n395), .A2(n371), .ZN(n392) );
  NAND2_X1 U503 ( .A1(n367), .A2(KEYINPUT85), .ZN(n393) );
  NAND2_X1 U504 ( .A1(n380), .A2(n410), .ZN(n394) );
  XNOR2_X1 U505 ( .A(n568), .B(KEYINPUT88), .ZN(n404) );
  XNOR2_X1 U506 ( .A(KEYINPUT41), .B(n614), .ZN(n760) );
  XNOR2_X1 U507 ( .A(n616), .B(KEYINPUT42), .ZN(n790) );
  NAND2_X1 U508 ( .A1(n666), .A2(KEYINPUT44), .ZN(n568) );
  NAND2_X1 U509 ( .A1(n398), .A2(n397), .ZN(n550) );
  INV_X1 U510 ( .A(n701), .ZN(n397) );
  INV_X1 U511 ( .A(n715), .ZN(n398) );
  AND2_X2 U512 ( .A1(n405), .A2(n404), .ZN(n403) );
  AND2_X2 U513 ( .A1(n555), .A2(n556), .ZN(n405) );
  NAND2_X1 U514 ( .A1(n632), .A2(n407), .ZN(n406) );
  INV_X1 U515 ( .A(n411), .ZN(n409) );
  NAND2_X1 U516 ( .A1(n575), .A2(KEYINPUT85), .ZN(n410) );
  XNOR2_X2 U517 ( .A(G113), .B(KEYINPUT71), .ZN(n415) );
  XNOR2_X2 U518 ( .A(n418), .B(n417), .ZN(n782) );
  NAND2_X1 U519 ( .A1(n375), .A2(n419), .ZN(n593) );
  INV_X1 U520 ( .A(n381), .ZN(n419) );
  AND2_X2 U521 ( .A1(n690), .A2(n450), .ZN(n426) );
  XNOR2_X1 U522 ( .A(n617), .B(KEYINPUT46), .ZN(n420) );
  XNOR2_X2 U523 ( .A(n591), .B(KEYINPUT77), .ZN(n611) );
  INV_X1 U524 ( .A(n733), .ZN(n424) );
  OR2_X1 U525 ( .A1(n690), .A2(n431), .ZN(n430) );
  NOR2_X1 U526 ( .A1(n426), .A2(n376), .ZN(n425) );
  XNOR2_X2 U527 ( .A(G143), .B(G128), .ZN(n464) );
  XNOR2_X2 U528 ( .A(n428), .B(G469), .ZN(n604) );
  INV_X1 U529 ( .A(n433), .ZN(n429) );
  BUF_X1 U530 ( .A(n491), .Z(n500) );
  AND2_X1 U531 ( .A1(n626), .A2(n625), .ZN(n434) );
  NOR2_X1 U532 ( .A1(n718), .A2(n434), .ZN(n435) );
  INV_X1 U533 ( .A(n736), .ZN(n454) );
  OR2_X1 U534 ( .A1(n641), .A2(n640), .ZN(n436) );
  INV_X1 U535 ( .A(KEYINPUT80), .ZN(n597) );
  INV_X1 U536 ( .A(KEYINPUT101), .ZN(n495) );
  XNOR2_X1 U537 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U538 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U539 ( .A(G140), .B(G110), .Z(n513) );
  XNOR2_X1 U540 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U541 ( .A(n469), .B(n468), .ZN(n471) );
  NAND2_X1 U542 ( .A1(n689), .A2(G475), .ZN(n647) );
  XNOR2_X1 U543 ( .A(n772), .B(n771), .ZN(n773) );
  XNOR2_X1 U544 ( .A(n613), .B(n612), .ZN(n791) );
  INV_X1 U545 ( .A(KEYINPUT60), .ZN(n650) );
  BUF_X1 U546 ( .A(n666), .Z(n667) );
  XNOR2_X2 U547 ( .A(G101), .B(KEYINPUT94), .ZN(n437) );
  XNOR2_X2 U548 ( .A(KEYINPUT95), .B(KEYINPUT3), .ZN(n438) );
  XNOR2_X1 U549 ( .A(n439), .B(KEYINPUT75), .ZN(n440) );
  XNOR2_X1 U550 ( .A(n464), .B(n441), .ZN(n443) );
  XNOR2_X1 U551 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U552 ( .A(n489), .B(n478), .ZN(n444) );
  XNOR2_X1 U553 ( .A(n445), .B(n444), .ZN(n446) );
  INV_X1 U554 ( .A(n641), .ZN(n575) );
  NAND2_X1 U555 ( .A1(n523), .A2(n448), .ZN(n451) );
  NAND2_X1 U556 ( .A1(n451), .A2(G210), .ZN(n449) );
  XNOR2_X1 U557 ( .A(n449), .B(KEYINPUT78), .ZN(n450) );
  NAND2_X1 U558 ( .A1(n451), .A2(G214), .ZN(n453) );
  INV_X1 U559 ( .A(KEYINPUT96), .ZN(n452) );
  XNOR2_X1 U560 ( .A(n453), .B(n452), .ZN(n736) );
  INV_X1 U561 ( .A(KEYINPUT90), .ZN(n455) );
  XNOR2_X2 U562 ( .A(n456), .B(n455), .ZN(n621) );
  XNOR2_X1 U563 ( .A(G898), .B(KEYINPUT97), .ZN(n783) );
  INV_X1 U564 ( .A(n580), .ZN(n457) );
  NAND2_X1 U565 ( .A1(n783), .A2(n457), .ZN(n458) );
  NAND2_X1 U566 ( .A1(n465), .A2(G952), .ZN(n584) );
  NAND2_X1 U567 ( .A1(n458), .A2(n584), .ZN(n461) );
  INV_X1 U568 ( .A(KEYINPUT14), .ZN(n459) );
  XNOR2_X1 U569 ( .A(n460), .B(n459), .ZN(n765) );
  INV_X1 U570 ( .A(n765), .ZN(n582) );
  NAND2_X1 U571 ( .A1(n461), .A2(n582), .ZN(n462) );
  NAND2_X1 U572 ( .A1(G217), .A2(n518), .ZN(n469) );
  XNOR2_X1 U573 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U574 ( .A(n490), .B(n472), .ZN(n680) );
  NOR2_X1 U575 ( .A1(G902), .A2(n680), .ZN(n473) );
  XNOR2_X1 U576 ( .A(G478), .B(n473), .ZN(n549) );
  XNOR2_X1 U577 ( .A(G143), .B(n661), .ZN(n476) );
  XNOR2_X1 U578 ( .A(n478), .B(n477), .ZN(n519) );
  XNOR2_X1 U579 ( .A(n507), .B(n519), .ZN(n652) );
  XNOR2_X1 U580 ( .A(n479), .B(n652), .ZN(n645) );
  NAND2_X1 U581 ( .A1(n645), .A2(n523), .ZN(n481) );
  XNOR2_X1 U582 ( .A(KEYINPUT13), .B(G475), .ZN(n480) );
  XNOR2_X1 U583 ( .A(n481), .B(n480), .ZN(n563) );
  AND2_X1 U584 ( .A1(n549), .A2(n563), .ZN(n739) );
  NAND2_X1 U585 ( .A1(n641), .A2(G234), .ZN(n482) );
  XNOR2_X1 U586 ( .A(n482), .B(KEYINPUT20), .ZN(n524) );
  AND2_X1 U587 ( .A1(n524), .A2(G221), .ZN(n484) );
  INV_X1 U588 ( .A(KEYINPUT21), .ZN(n483) );
  XNOR2_X1 U589 ( .A(n484), .B(n483), .ZN(n744) );
  INV_X1 U590 ( .A(n744), .ZN(n539) );
  AND2_X1 U591 ( .A1(n739), .A2(n539), .ZN(n485) );
  NAND2_X1 U592 ( .A1(n543), .A2(n485), .ZN(n488) );
  XNOR2_X1 U593 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n486) );
  XNOR2_X1 U594 ( .A(n486), .B(KEYINPUT67), .ZN(n487) );
  XNOR2_X2 U595 ( .A(n488), .B(n487), .ZN(n535) );
  XNOR2_X1 U596 ( .A(n653), .B(G146), .ZN(n510) );
  NAND2_X1 U597 ( .A1(n492), .A2(G210), .ZN(n493) );
  XNOR2_X1 U598 ( .A(n494), .B(n493), .ZN(n498) );
  XNOR2_X1 U599 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U600 ( .A(n510), .B(n501), .ZN(n669) );
  INV_X1 U601 ( .A(KEYINPUT102), .ZN(n502) );
  XNOR2_X1 U602 ( .A(n502), .B(G472), .ZN(n503) );
  XNOR2_X2 U603 ( .A(n504), .B(n503), .ZN(n577) );
  XNOR2_X1 U604 ( .A(n577), .B(KEYINPUT6), .ZN(n618) );
  INV_X1 U605 ( .A(n618), .ZN(n505) );
  AND2_X2 U606 ( .A1(n535), .A2(n505), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n465), .A2(G227), .ZN(n506) );
  XNOR2_X1 U608 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U609 ( .A(n511), .B(n510), .ZN(n685) );
  XOR2_X1 U610 ( .A(n513), .B(n512), .Z(n517) );
  XOR2_X1 U611 ( .A(KEYINPUT99), .B(KEYINPUT24), .Z(n515) );
  XNOR2_X1 U612 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U613 ( .A(n517), .B(n516), .ZN(n522) );
  NAND2_X1 U614 ( .A1(G221), .A2(n518), .ZN(n520) );
  NAND2_X1 U615 ( .A1(n675), .A2(n523), .ZN(n527) );
  AND2_X1 U616 ( .A1(n524), .A2(G217), .ZN(n525) );
  XNOR2_X1 U617 ( .A(KEYINPUT25), .B(n525), .ZN(n526) );
  XNOR2_X1 U618 ( .A(n527), .B(n526), .ZN(n540) );
  BUF_X1 U619 ( .A(n540), .Z(n601) );
  INV_X1 U620 ( .A(n601), .ZN(n743) );
  NAND2_X1 U621 ( .A1(n364), .A2(n743), .ZN(n528) );
  XNOR2_X1 U622 ( .A(n528), .B(KEYINPUT107), .ZN(n529) );
  NAND2_X1 U623 ( .A1(n553), .A2(n529), .ZN(n532) );
  INV_X1 U624 ( .A(KEYINPUT66), .ZN(n530) );
  XNOR2_X1 U625 ( .A(n530), .B(KEYINPUT32), .ZN(n531) );
  XNOR2_X2 U626 ( .A(n532), .B(n531), .ZN(n665) );
  NAND2_X1 U627 ( .A1(n577), .A2(n743), .ZN(n533) );
  NOR2_X1 U628 ( .A1(n364), .A2(n533), .ZN(n534) );
  AND2_X1 U629 ( .A1(n535), .A2(n534), .ZN(n664) );
  NAND2_X1 U630 ( .A1(n540), .A2(n539), .ZN(n541) );
  INV_X1 U631 ( .A(n577), .ZN(n754) );
  NOR2_X1 U632 ( .A1(n588), .A2(n754), .ZN(n542) );
  AND2_X1 U633 ( .A1(n560), .A2(n542), .ZN(n701) );
  BUF_X1 U634 ( .A(n543), .Z(n545) );
  NAND2_X1 U635 ( .A1(n557), .A2(n754), .ZN(n756) );
  INV_X1 U636 ( .A(n756), .ZN(n544) );
  NAND2_X1 U637 ( .A1(n545), .A2(n544), .ZN(n548) );
  INV_X1 U638 ( .A(KEYINPUT103), .ZN(n546) );
  XNOR2_X1 U639 ( .A(n546), .B(KEYINPUT31), .ZN(n547) );
  INV_X1 U640 ( .A(n549), .ZN(n564) );
  AND2_X1 U641 ( .A1(n563), .A2(n564), .ZN(n714) );
  NAND2_X1 U642 ( .A1(n550), .A2(n576), .ZN(n551) );
  XNOR2_X1 U643 ( .A(n551), .B(KEYINPUT106), .ZN(n554) );
  NOR2_X1 U644 ( .A1(n364), .A2(n743), .ZN(n552) );
  NAND2_X1 U645 ( .A1(n553), .A2(n552), .ZN(n700) );
  AND2_X1 U646 ( .A1(n554), .A2(n700), .ZN(n555) );
  NAND2_X1 U647 ( .A1(n557), .A2(n618), .ZN(n559) );
  XNOR2_X1 U648 ( .A(KEYINPUT92), .B(KEYINPUT33), .ZN(n558) );
  NAND2_X1 U649 ( .A1(n560), .A2(n735), .ZN(n562) );
  XNOR2_X1 U650 ( .A(n562), .B(n561), .ZN(n566) );
  INV_X1 U651 ( .A(n563), .ZN(n565) );
  AND2_X1 U652 ( .A1(n565), .A2(n564), .ZN(n592) );
  NAND2_X1 U653 ( .A1(n566), .A2(n592), .ZN(n567) );
  INV_X1 U654 ( .A(KEYINPUT44), .ZN(n569) );
  NOR2_X1 U655 ( .A1(n665), .A2(n664), .ZN(n573) );
  NAND2_X1 U656 ( .A1(n737), .A2(KEYINPUT47), .ZN(n596) );
  XNOR2_X1 U657 ( .A(KEYINPUT30), .B(KEYINPUT112), .ZN(n578) );
  XNOR2_X1 U658 ( .A(n579), .B(n578), .ZN(n590) );
  NOR2_X1 U659 ( .A1(G900), .A2(n580), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U661 ( .A(KEYINPUT108), .B(n583), .Z(n586) );
  NOR2_X1 U662 ( .A1(n765), .A2(n584), .ZN(n585) );
  NOR2_X1 U663 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U664 ( .A(KEYINPUT79), .B(n587), .Z(n599) );
  NOR2_X1 U665 ( .A1(n588), .A2(n599), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U667 ( .A(n592), .ZN(n594) );
  NOR2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n611), .A2(n595), .ZN(n708) );
  NAND2_X1 U670 ( .A1(n596), .A2(n708), .ZN(n598) );
  XNOR2_X1 U671 ( .A(KEYINPUT113), .B(KEYINPUT28), .ZN(n603) );
  OR2_X1 U672 ( .A1(n744), .A2(n599), .ZN(n600) );
  NOR2_X1 U673 ( .A1(n601), .A2(n600), .ZN(n619) );
  AND2_X1 U674 ( .A1(n619), .A2(n754), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n603), .B(n602), .ZN(n606) );
  INV_X1 U676 ( .A(n604), .ZN(n605) );
  OR2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n615) );
  OR2_X1 U678 ( .A1(n615), .A2(n607), .ZN(n710) );
  NAND2_X1 U679 ( .A1(n710), .A2(KEYINPUT47), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U681 ( .A(KEYINPUT38), .B(n593), .Z(n733) );
  NAND2_X1 U682 ( .A1(n631), .A2(n712), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n739), .A2(n454), .ZN(n732) );
  NOR2_X1 U684 ( .A1(n733), .A2(n732), .ZN(n614) );
  NOR2_X1 U685 ( .A1(n760), .A2(n615), .ZN(n616) );
  INV_X1 U686 ( .A(n364), .ZN(n624) );
  NAND2_X1 U687 ( .A1(n619), .A2(n618), .ZN(n620) );
  INV_X1 U688 ( .A(n712), .ZN(n709) );
  NOR2_X1 U689 ( .A1(n620), .A2(n709), .ZN(n635) );
  NAND2_X1 U690 ( .A1(n621), .A2(n635), .ZN(n622) );
  XNOR2_X1 U691 ( .A(n622), .B(KEYINPUT36), .ZN(n623) );
  NOR2_X1 U692 ( .A1(n624), .A2(n623), .ZN(n718) );
  XOR2_X1 U693 ( .A(KEYINPUT47), .B(KEYINPUT70), .Z(n626) );
  NOR2_X1 U694 ( .A1(n710), .A2(n737), .ZN(n625) );
  INV_X1 U695 ( .A(KEYINPUT48), .ZN(n627) );
  NAND2_X1 U696 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U697 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U698 ( .A1(n631), .A2(n714), .ZN(n721) );
  XNOR2_X1 U699 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n633) );
  XNOR2_X1 U700 ( .A(n633), .B(KEYINPUT43), .ZN(n637) );
  NOR2_X1 U701 ( .A1(n736), .A2(n364), .ZN(n634) );
  NAND2_X1 U702 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U703 ( .A(n637), .B(n636), .Z(n638) );
  NAND2_X1 U704 ( .A1(n638), .A2(n593), .ZN(n639) );
  XNOR2_X1 U705 ( .A(n639), .B(KEYINPUT111), .ZN(n789) );
  INV_X1 U706 ( .A(KEYINPUT2), .ZN(n640) );
  NAND2_X1 U707 ( .A1(n372), .A2(KEYINPUT2), .ZN(n642) );
  INV_X1 U708 ( .A(n380), .ZN(n775) );
  AND2_X2 U709 ( .A1(n643), .A2(n727), .ZN(n689) );
  XNOR2_X1 U710 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n644) );
  XNOR2_X1 U711 ( .A(n647), .B(n646), .ZN(n649) );
  INV_X1 U712 ( .A(G952), .ZN(n648) );
  NAND2_X1 U713 ( .A1(n649), .A2(n696), .ZN(n651) );
  XNOR2_X1 U714 ( .A(n651), .B(n650), .ZN(G60) );
  XNOR2_X1 U715 ( .A(n653), .B(n652), .ZN(n654) );
  XOR2_X1 U716 ( .A(KEYINPUT127), .B(n654), .Z(n656) );
  XOR2_X1 U717 ( .A(n656), .B(n372), .Z(n655) );
  NAND2_X1 U718 ( .A1(n655), .A2(n465), .ZN(n660) );
  XNOR2_X1 U719 ( .A(G227), .B(n656), .ZN(n657) );
  NAND2_X1 U720 ( .A1(n657), .A2(G900), .ZN(n658) );
  NAND2_X1 U721 ( .A1(n658), .A2(G953), .ZN(n659) );
  NAND2_X1 U722 ( .A1(n660), .A2(n659), .ZN(G72) );
  NAND2_X1 U723 ( .A1(n701), .A2(n712), .ZN(n662) );
  XNOR2_X1 U724 ( .A(n662), .B(n661), .ZN(G6) );
  XNOR2_X1 U725 ( .A(n664), .B(n663), .ZN(G12) );
  XOR2_X1 U726 ( .A(n665), .B(G119), .Z(G21) );
  XOR2_X1 U727 ( .A(n667), .B(G122), .Z(G24) );
  NAND2_X1 U728 ( .A1(n689), .A2(G472), .ZN(n671) );
  XOR2_X1 U729 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n668) );
  XNOR2_X1 U730 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U731 ( .A1(n672), .A2(n696), .ZN(n674) );
  XOR2_X1 U732 ( .A(KEYINPUT93), .B(KEYINPUT63), .Z(n673) );
  XNOR2_X1 U733 ( .A(n674), .B(n673), .ZN(G57) );
  BUF_X2 U734 ( .A(n689), .Z(n683) );
  NAND2_X1 U735 ( .A1(n683), .A2(G217), .ZN(n677) );
  XNOR2_X1 U736 ( .A(n675), .B(KEYINPUT124), .ZN(n676) );
  XNOR2_X1 U737 ( .A(n677), .B(n676), .ZN(n678) );
  AND2_X1 U738 ( .A1(n678), .A2(n696), .ZN(G66) );
  NAND2_X1 U739 ( .A1(n683), .A2(G478), .ZN(n679) );
  XNOR2_X1 U740 ( .A(n680), .B(n679), .ZN(n682) );
  INV_X1 U741 ( .A(n696), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n682), .A2(n681), .ZN(G63) );
  NAND2_X1 U743 ( .A1(n683), .A2(G469), .ZN(n687) );
  XNOR2_X1 U744 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n684) );
  XNOR2_X1 U745 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U746 ( .A(n687), .B(n686), .ZN(n688) );
  AND2_X1 U747 ( .A1(n688), .A2(n696), .ZN(G54) );
  NAND2_X1 U748 ( .A1(n689), .A2(G210), .ZN(n695) );
  BUF_X1 U749 ( .A(n690), .Z(n693) );
  XNOR2_X1 U750 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n691) );
  XOR2_X1 U751 ( .A(n691), .B(KEYINPUT55), .Z(n692) );
  XNOR2_X1 U752 ( .A(n695), .B(n694), .ZN(n697) );
  NAND2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n699) );
  XOR2_X1 U754 ( .A(KEYINPUT86), .B(KEYINPUT56), .Z(n698) );
  XNOR2_X1 U755 ( .A(n699), .B(n698), .ZN(G51) );
  XNOR2_X1 U756 ( .A(G101), .B(n700), .ZN(G3) );
  NAND2_X1 U757 ( .A1(n701), .A2(n714), .ZN(n703) );
  XOR2_X1 U758 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n702) );
  XNOR2_X1 U759 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U760 ( .A(G107), .B(n704), .ZN(G9) );
  INV_X1 U761 ( .A(n714), .ZN(n705) );
  NOR2_X1 U762 ( .A1(n710), .A2(n705), .ZN(n707) );
  XNOR2_X1 U763 ( .A(G128), .B(KEYINPUT29), .ZN(n706) );
  XNOR2_X1 U764 ( .A(n707), .B(n706), .ZN(G30) );
  XNOR2_X1 U765 ( .A(G143), .B(n708), .ZN(G45) );
  NOR2_X1 U766 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U767 ( .A(G146), .B(n711), .Z(G48) );
  NAND2_X1 U768 ( .A1(n715), .A2(n712), .ZN(n713) );
  XNOR2_X1 U769 ( .A(n713), .B(G113), .ZN(G15) );
  XOR2_X1 U770 ( .A(G116), .B(KEYINPUT115), .Z(n717) );
  NAND2_X1 U771 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U772 ( .A(n717), .B(n716), .ZN(G18) );
  XNOR2_X1 U773 ( .A(n718), .B(KEYINPUT37), .ZN(n719) );
  XNOR2_X1 U774 ( .A(n719), .B(KEYINPUT116), .ZN(n720) );
  XNOR2_X1 U775 ( .A(G125), .B(n720), .ZN(G27) );
  XNOR2_X1 U776 ( .A(G134), .B(n721), .ZN(G36) );
  XNOR2_X1 U777 ( .A(KEYINPUT81), .B(KEYINPUT2), .ZN(n724) );
  INV_X1 U778 ( .A(n724), .ZN(n722) );
  NOR2_X1 U779 ( .A1(n372), .A2(n722), .ZN(n723) );
  XNOR2_X1 U780 ( .A(n723), .B(KEYINPUT83), .ZN(n726) );
  NAND2_X1 U781 ( .A1(n775), .A2(n724), .ZN(n725) );
  NAND2_X1 U782 ( .A1(n726), .A2(n725), .ZN(n729) );
  INV_X1 U783 ( .A(n727), .ZN(n728) );
  NOR2_X1 U784 ( .A1(n729), .A2(n728), .ZN(n770) );
  INV_X1 U785 ( .A(n735), .ZN(n730) );
  NOR2_X1 U786 ( .A1(n730), .A2(n760), .ZN(n731) );
  XNOR2_X1 U787 ( .A(n731), .B(KEYINPUT121), .ZN(n768) );
  NAND2_X1 U788 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U789 ( .A1(n735), .A2(n734), .ZN(n741) );
  NOR2_X1 U790 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U792 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U793 ( .A(n742), .B(KEYINPUT120), .ZN(n762) );
  NAND2_X1 U794 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U795 ( .A(n745), .B(KEYINPUT49), .ZN(n746) );
  XNOR2_X1 U796 ( .A(KEYINPUT117), .B(n746), .ZN(n752) );
  NOR2_X1 U797 ( .A1(n748), .A2(n364), .ZN(n749) );
  XOR2_X1 U798 ( .A(KEYINPUT50), .B(n749), .Z(n750) );
  XNOR2_X1 U799 ( .A(KEYINPUT118), .B(n750), .ZN(n751) );
  NAND2_X1 U800 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U801 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U802 ( .A(n755), .B(KEYINPUT119), .ZN(n757) );
  NAND2_X1 U803 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U804 ( .A(KEYINPUT51), .B(n758), .ZN(n759) );
  NOR2_X1 U805 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U806 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U807 ( .A(n763), .B(KEYINPUT52), .ZN(n764) );
  NOR2_X1 U808 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U809 ( .A1(n766), .A2(G952), .ZN(n767) );
  NAND2_X1 U810 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U811 ( .A1(n770), .A2(n769), .ZN(n772) );
  NOR2_X1 U812 ( .A1(G953), .A2(n773), .ZN(n774) );
  XNOR2_X1 U813 ( .A(KEYINPUT53), .B(n774), .ZN(G75) );
  NOR2_X1 U814 ( .A1(n775), .A2(G953), .ZN(n780) );
  NAND2_X1 U815 ( .A1(G224), .A2(G953), .ZN(n776) );
  XNOR2_X1 U816 ( .A(n776), .B(KEYINPUT61), .ZN(n777) );
  XNOR2_X1 U817 ( .A(n777), .B(KEYINPUT125), .ZN(n778) );
  NOR2_X1 U818 ( .A1(n783), .A2(n778), .ZN(n779) );
  NOR2_X1 U819 ( .A1(n780), .A2(n779), .ZN(n788) );
  XOR2_X1 U820 ( .A(n782), .B(n369), .Z(n785) );
  NAND2_X1 U821 ( .A1(n783), .A2(G953), .ZN(n784) );
  NAND2_X1 U822 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U823 ( .A(n786), .B(KEYINPUT126), .ZN(n787) );
  XNOR2_X1 U824 ( .A(n788), .B(n787), .ZN(G69) );
  XOR2_X1 U825 ( .A(G140), .B(n789), .Z(G42) );
  XOR2_X1 U826 ( .A(G137), .B(n790), .Z(G39) );
  BUF_X1 U827 ( .A(n791), .Z(n792) );
  XOR2_X1 U828 ( .A(G131), .B(n792), .Z(G33) );
endmodule

