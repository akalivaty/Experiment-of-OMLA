//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n581, new_n582, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n605, new_n606, new_n607, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n642, new_n643, new_n646,
    new_n648, new_n649, new_n650, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XNOR2_X1  g016(.A(KEYINPUT68), .B(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT69), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT71), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n469), .B2(G137), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n462), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  NOR3_X1   g048(.A1(new_n472), .A2(KEYINPUT71), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n464), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(G125), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n476), .A2(KEYINPUT70), .B1(G113), .B2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n471), .A2(new_n478), .A3(G125), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n462), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(G160));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n468), .A2(new_n462), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n469), .A2(G136), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n462), .B1(KEYINPUT73), .B2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n491), .A2(KEYINPUT73), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT72), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n471), .A2(new_n497), .A3(G126), .A4(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n494), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n466), .B2(new_n467), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT74), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n501), .B(new_n503), .C1(new_n467), .C2(new_n466), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT76), .ZN(new_n510));
  AND3_X1   g085(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(G543), .B1(KEYINPUT75), .B2(KEYINPUT5), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n510), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT75), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT6), .B(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n522), .A2(KEYINPUT76), .A3(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G88), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G62), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n513), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n515), .ZN(new_n530));
  NAND2_X1  g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n519), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n529), .A2(G651), .B1(G50), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n526), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  XNOR2_X1  g110(.A(KEYINPUT79), .B(G89), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n517), .A2(new_n524), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n532), .A2(G51), .ZN(new_n541));
  NAND2_X1  g116(.A1(G63), .A2(G651), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(KEYINPUT77), .B1(new_n522), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT77), .ZN(new_n545));
  AOI211_X1 g120(.A(new_n545), .B(new_n542), .C1(new_n520), .C2(new_n521), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n541), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(KEYINPUT78), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n545), .B1(new_n513), .B2(new_n542), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n522), .A2(KEYINPUT77), .A3(new_n543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT78), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n551), .A2(new_n552), .A3(new_n541), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n540), .B1(new_n548), .B2(new_n553), .ZN(G168));
  NAND3_X1  g129(.A1(new_n517), .A2(G90), .A3(new_n524), .ZN(new_n555));
  NAND2_X1  g130(.A1(G77), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G64), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n513), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  INV_X1    g134(.A(G52), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n523), .A2(G543), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n555), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(G301));
  INV_X1    g137(.A(G301), .ZN(G171));
  XNOR2_X1  g138(.A(KEYINPUT82), .B(G81), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n525), .A2(new_n564), .B1(G43), .B2(new_n532), .ZN(new_n565));
  INV_X1    g140(.A(G56), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n520), .B2(new_n521), .ZN(new_n567));
  NAND2_X1  g142(.A1(G68), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT80), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n571), .B(new_n568), .C1(new_n513), .C2(new_n566), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n570), .A2(new_n572), .A3(KEYINPUT81), .A4(G651), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(new_n572), .A3(G651), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n565), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G860), .ZN(G153));
  NAND4_X1  g154(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g155(.A1(G1), .A2(G3), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT8), .ZN(new_n582));
  NAND4_X1  g157(.A1(G319), .A2(G483), .A3(G661), .A4(new_n582), .ZN(G188));
  INV_X1    g158(.A(G65), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n585), .B1(new_n511), .B2(new_n512), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n520), .A2(KEYINPUT84), .A3(new_n521), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G78), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT83), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G53), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT9), .B1(new_n561), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT9), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n532), .A2(new_n592), .A3(new_n595), .A4(G53), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n517), .A2(G91), .A3(new_n524), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n591), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT85), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n591), .A2(new_n597), .A3(KEYINPUT85), .A4(new_n598), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G299));
  AND2_X1   g179(.A1(new_n537), .A2(new_n539), .ZN(new_n605));
  AOI221_X4 g180(.A(KEYINPUT78), .B1(G51), .B2(new_n532), .C1(new_n549), .C2(new_n550), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n552), .B1(new_n551), .B2(new_n541), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(G286));
  NAND2_X1  g183(.A1(new_n525), .A2(G87), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n522), .A2(G74), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n610), .A2(G651), .B1(G49), .B2(new_n532), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT86), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n609), .A2(KEYINPUT86), .A3(new_n611), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(G288));
  NAND2_X1  g192(.A1(G73), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G61), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n513), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n620), .A2(G651), .B1(G48), .B2(new_n532), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n517), .A2(G86), .A3(new_n524), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(G305));
  NAND2_X1  g198(.A1(new_n525), .A2(G85), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n532), .A2(G47), .ZN(new_n625));
  INV_X1    g200(.A(G651), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n627), .ZN(G290));
  NAND2_X1  g203(.A1(G301), .A2(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n532), .A2(G54), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n586), .A2(new_n587), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n631), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n630), .B1(new_n632), .B2(new_n626), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n517), .A2(G92), .A3(new_n524), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT10), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n634), .A2(new_n635), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n629), .B1(new_n639), .B2(G868), .ZN(G284));
  OAI21_X1  g215(.A(new_n629), .B1(new_n639), .B2(G868), .ZN(G321));
  INV_X1    g216(.A(G868), .ZN(new_n642));
  NOR2_X1   g217(.A1(G286), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n603), .ZN(G297));
  AOI21_X1  g219(.A(new_n643), .B1(new_n642), .B2(new_n603), .ZN(G280));
  INV_X1    g220(.A(G559), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n639), .B1(new_n646), .B2(G860), .ZN(G148));
  NAND2_X1  g222(.A1(new_n577), .A2(new_n642), .ZN(new_n648));
  INV_X1    g223(.A(new_n639), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n649), .A2(G559), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n648), .B1(new_n650), .B2(new_n642), .ZN(G323));
  XNOR2_X1  g226(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g227(.A1(new_n471), .A2(new_n463), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT13), .ZN(new_n656));
  INV_X1    g231(.A(G2100), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n469), .A2(G135), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n485), .A2(G123), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n462), .A2(G111), .ZN(new_n662));
  OAI21_X1  g237(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n660), .B(new_n661), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(G2096), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n658), .A2(new_n659), .A3(new_n666), .ZN(G156));
  XNOR2_X1  g242(.A(G2427), .B(G2438), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2430), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT15), .B(G2435), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(KEYINPUT14), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2451), .B(G2454), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT16), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2443), .B(G2446), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1341), .B(G1348), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(KEYINPUT88), .B1(new_n678), .B2(new_n680), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(G14), .B1(new_n678), .B2(new_n680), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(G401));
  XNOR2_X1  g262(.A(G2084), .B(G2090), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT89), .ZN(new_n689));
  XNOR2_X1  g264(.A(G2067), .B(G2678), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(KEYINPUT18), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G2072), .B(G2078), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT90), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(new_n657), .ZN(new_n696));
  OAI21_X1  g271(.A(KEYINPUT17), .B1(new_n689), .B2(new_n691), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n689), .B2(new_n691), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n698), .A2(KEYINPUT18), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(new_n665), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n696), .B(new_n700), .ZN(G227));
  XNOR2_X1  g276(.A(G1971), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT19), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1961), .B(G1966), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT91), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1956), .B(G2474), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n704), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT20), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n704), .B1(new_n706), .B2(new_n708), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n706), .A2(new_n708), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n710), .B(new_n713), .C1(new_n703), .C2(new_n712), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT92), .ZN(new_n715));
  XOR2_X1   g290(.A(G1981), .B(G1986), .Z(new_n716));
  XNOR2_X1  g291(.A(G1991), .B(G1996), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n715), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(G229));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G23), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n609), .A2(new_n611), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n723), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT33), .B(G1976), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(KEYINPUT94), .ZN(new_n729));
  NOR2_X1   g304(.A1(G6), .A2(G16), .ZN(new_n730));
  INV_X1    g305(.A(G305), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G16), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT32), .ZN(new_n733));
  INV_X1    g308(.A(G1981), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n728), .A2(KEYINPUT94), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n723), .A2(G22), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT95), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G303), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1971), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n729), .A2(new_n735), .A3(new_n736), .A4(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT34), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(KEYINPUT34), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n469), .A2(G131), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n485), .A2(G119), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n462), .A2(G107), .ZN(new_n746));
  OAI21_X1  g321(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  MUX2_X1   g323(.A(G25), .B(new_n748), .S(G29), .Z(new_n749));
  XOR2_X1   g324(.A(KEYINPUT35), .B(G1991), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G16), .A2(G24), .ZN(new_n752));
  XOR2_X1   g327(.A(G290), .B(KEYINPUT93), .Z(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G16), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G1986), .Z(new_n755));
  NAND4_X1  g330(.A1(new_n742), .A2(new_n743), .A3(new_n751), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT36), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT99), .B(KEYINPUT26), .Z(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n463), .A2(G105), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n485), .A2(G129), .ZN(new_n763));
  INV_X1    g338(.A(G141), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n472), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G29), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n767), .B2(G32), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT27), .B(G1996), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT100), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT30), .B(G28), .ZN(new_n773));
  OR2_X1    g348(.A1(KEYINPUT31), .A2(G11), .ZN(new_n774));
  NAND2_X1  g349(.A1(KEYINPUT31), .A2(G11), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n773), .A2(new_n767), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n664), .B2(new_n767), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n769), .B2(new_n771), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n767), .A2(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n767), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT29), .B(G2090), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n767), .A2(G26), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n469), .A2(G140), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n485), .A2(G128), .ZN(new_n787));
  OR2_X1    g362(.A1(G104), .A2(G2105), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n788), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n785), .B1(new_n791), .B2(new_n767), .ZN(new_n792));
  INV_X1    g367(.A(G2067), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AND4_X1   g369(.A1(new_n772), .A2(new_n778), .A3(new_n782), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n767), .A2(G33), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT97), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT25), .Z(new_n799));
  AOI22_X1  g374(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n800));
  INV_X1    g375(.A(G139), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n800), .A2(new_n462), .B1(new_n801), .B2(new_n472), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n796), .B1(new_n803), .B2(new_n767), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G2072), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n723), .A2(G5), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G171), .B2(new_n723), .ZN(new_n807));
  INV_X1    g382(.A(G1961), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n767), .A2(G27), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G164), .B2(new_n767), .ZN(new_n811));
  INV_X1    g386(.A(G2078), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n795), .A2(new_n805), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n723), .A2(G19), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n578), .B2(new_n723), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1341), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n723), .A2(G20), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT23), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n603), .B2(new_n723), .ZN(new_n820));
  INV_X1    g395(.A(G1956), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n639), .A2(new_n723), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G4), .B2(new_n723), .ZN(new_n825));
  INV_X1    g400(.A(G1348), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n723), .A2(G21), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G168), .B2(new_n723), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT101), .B(G1966), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n827), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G34), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n834), .A2(KEYINPUT24), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(KEYINPUT24), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n767), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G160), .B2(new_n767), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT98), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G2084), .ZN(new_n840));
  NOR4_X1   g415(.A1(new_n814), .A2(new_n823), .A3(new_n833), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n757), .A2(new_n841), .ZN(G150));
  INV_X1    g417(.A(G150), .ZN(G311));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  INV_X1    g419(.A(G67), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n513), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n846), .A2(G651), .B1(G55), .B2(new_n532), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n517), .A2(G93), .A3(new_n524), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n639), .A2(G559), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n577), .A2(new_n849), .ZN(new_n856));
  INV_X1    g431(.A(new_n849), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n857), .A2(new_n565), .A3(new_n573), .A4(new_n576), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n855), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  INV_X1    g437(.A(G860), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n861), .B2(KEYINPUT39), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n852), .B1(new_n862), .B2(new_n864), .ZN(G145));
  INV_X1    g440(.A(new_n803), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n505), .A2(new_n867), .A3(new_n506), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n505), .B2(new_n506), .ZN(new_n869));
  OAI211_X1 g444(.A(KEYINPUT105), .B(new_n499), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n506), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n503), .B1(new_n471), .B2(new_n501), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT104), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n505), .A2(new_n867), .A3(new_n506), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT105), .B1(new_n876), .B2(new_n499), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n791), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n766), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n499), .B1(new_n868), .B2(new_n869), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(new_n790), .A3(new_n870), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n878), .A2(new_n879), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n879), .B1(new_n878), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n866), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n748), .B(new_n655), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n485), .A2(G130), .ZN(new_n888));
  OR2_X1    g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n889), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(G142), .B2(new_n469), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n887), .B(new_n892), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n871), .A2(new_n877), .A3(new_n791), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n790), .B1(new_n882), .B2(new_n870), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n766), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n878), .A2(new_n879), .A3(new_n883), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n803), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n886), .A2(new_n893), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT106), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n886), .A2(new_n898), .A3(new_n901), .A4(new_n893), .ZN(new_n902));
  INV_X1    g477(.A(new_n893), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n884), .A2(new_n885), .A3(new_n866), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n803), .B1(new_n896), .B2(new_n897), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n664), .B(new_n488), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(G160), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n900), .A2(new_n902), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT107), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n893), .B1(new_n886), .B2(new_n898), .ZN(new_n911));
  INV_X1    g486(.A(new_n908), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n913), .A2(new_n914), .A3(new_n902), .A4(new_n900), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n899), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n912), .B1(new_n917), .B2(new_n911), .ZN(new_n918));
  INV_X1    g493(.A(G37), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT108), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n916), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(KEYINPUT40), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n927));
  AOI211_X1 g502(.A(KEYINPUT108), .B(new_n920), .C1(new_n910), .C2(new_n915), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n924), .B1(new_n916), .B2(new_n921), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n926), .A2(new_n930), .ZN(G395));
  NAND2_X1  g506(.A1(new_n856), .A2(new_n858), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n650), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n603), .A2(KEYINPUT109), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n601), .A2(new_n935), .A3(new_n602), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n649), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n603), .A2(KEYINPUT109), .A3(new_n639), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n937), .A2(KEYINPUT41), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT41), .B1(new_n937), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n933), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n859), .B(new_n650), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n938), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(G290), .B(new_n731), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n725), .B(G303), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n950), .B(new_n951), .Z(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n946), .A2(new_n952), .A3(new_n948), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(G868), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n857), .A2(G868), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(G295));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n957), .B2(new_n959), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n642), .B1(new_n954), .B2(new_n955), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n963), .A2(KEYINPUT110), .A3(new_n958), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n962), .A2(new_n964), .ZN(G331));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n939), .A2(new_n940), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT112), .B1(G168), .B2(G301), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n969));
  NAND3_X1  g544(.A1(G286), .A2(G171), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(G301), .B(new_n605), .C1(new_n607), .C2(new_n606), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT111), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n974));
  NAND3_X1  g549(.A1(G168), .A2(new_n974), .A3(G301), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n859), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n971), .A2(new_n976), .A3(new_n932), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n967), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n943), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(KEYINPUT113), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n971), .A2(new_n976), .A3(new_n932), .A4(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n982), .A2(new_n983), .A3(new_n978), .A4(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(new_n953), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n981), .A2(new_n986), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n919), .B1(new_n989), .B2(new_n952), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n966), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(G37), .B1(new_n987), .B2(new_n953), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n983), .A2(new_n978), .A3(new_n985), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n967), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n980), .B2(new_n943), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n982), .A2(new_n978), .A3(KEYINPUT114), .A4(new_n979), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n998), .A2(KEYINPUT115), .A3(new_n952), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT115), .B1(new_n998), .B2(new_n952), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n992), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n991), .B1(new_n1001), .B2(new_n966), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT44), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n966), .B(new_n992), .C1(new_n999), .C2(new_n1000), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT43), .B1(new_n988), .B2(new_n990), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1003), .A2(new_n1008), .ZN(G397));
  INV_X1    g584(.A(KEYINPUT126), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n880), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n476), .A2(KEYINPUT70), .ZN(new_n1013));
  NAND2_X1  g588(.A1(G113), .A2(G2104), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n479), .ZN(new_n1016));
  OAI21_X1  g591(.A(G2105), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n469), .A2(new_n465), .A3(G137), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT71), .B1(new_n472), .B2(new_n473), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1018), .A2(new_n1019), .B1(G101), .B2(new_n463), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(new_n1020), .A3(G40), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1012), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G305), .A2(G1981), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT119), .B(G1981), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1025), .B(KEYINPUT49), .C1(G305), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT49), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1025), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G305), .A2(new_n1026), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1024), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n1033));
  INV_X1    g608(.A(G40), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n475), .A2(new_n480), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n876), .B2(new_n499), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n725), .A2(G1976), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1037), .A2(new_n1038), .A3(G8), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1032), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1039), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1033), .B1(new_n616), .B2(G1976), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT118), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1042), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n1039), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1040), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G166), .A2(new_n1023), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n1049));
  OR2_X1    g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(KEYINPUT117), .B2(KEYINPUT55), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n508), .A2(new_n1011), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1035), .B1(KEYINPUT50), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1036), .A2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1055), .A2(G2090), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1021), .B1(new_n1059), .B2(new_n1054), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n882), .A2(KEYINPUT45), .A3(new_n1011), .A4(new_n870), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1971), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1053), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1021), .B1(KEYINPUT50), .B2(new_n1054), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1036), .A2(new_n1056), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(G2090), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1052), .B(G8), .C1(new_n1068), .C2(new_n1062), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1047), .A2(new_n1064), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1060), .A2(new_n1061), .A3(new_n812), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1071), .A2(new_n1072), .B1(new_n1067), .B2(new_n808), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n1011), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1035), .B(new_n1074), .C1(new_n1036), .C2(KEYINPUT45), .ZN(new_n1075));
  OR3_X1    g650(.A1(new_n1075), .A2(new_n1072), .A3(G2078), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1966), .ZN(new_n1080));
  NAND3_X1  g655(.A1(G160), .A2(new_n1074), .A3(G40), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT45), .B1(new_n880), .B2(new_n1011), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1075), .A2(KEYINPUT120), .A3(new_n1080), .ZN(new_n1086));
  INV_X1    g661(.A(G2084), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1065), .A2(new_n1087), .A3(new_n1066), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1085), .A2(G168), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1089), .A2(new_n1090), .A3(G8), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1085), .A2(new_n1088), .A3(new_n1086), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G286), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1093), .A2(G8), .A3(new_n1089), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1094), .B2(KEYINPUT51), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT62), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1070), .B(new_n1079), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(KEYINPUT51), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1091), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(KEYINPUT62), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1010), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT122), .B1(new_n1037), .B2(G2067), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1022), .A2(new_n1104), .A3(new_n793), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1348), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT123), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1067), .A2(new_n826), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1109), .A2(new_n1103), .A3(new_n1110), .A4(new_n1105), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n821), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1060), .A2(new_n1061), .A3(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n599), .B(KEYINPUT57), .Z(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1108), .A2(new_n1111), .A3(new_n639), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1115), .B(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(KEYINPUT60), .A3(new_n649), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1121), .A2(KEYINPUT61), .A3(new_n1116), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1116), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1115), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(G1996), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1060), .A2(new_n1061), .A3(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT58), .B(G1341), .Z(new_n1132));
  NAND2_X1  g707(.A1(new_n1037), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n577), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1124), .A2(new_n1125), .A3(new_n1129), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1108), .A2(new_n1111), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1139), .A2(new_n1140), .A3(new_n649), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1122), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1073), .A2(G301), .A3(new_n1076), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT54), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1072), .A2(G2078), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n882), .A2(new_n1011), .A3(new_n870), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1021), .B1(new_n1146), .B2(new_n1059), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1061), .B(new_n1145), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1073), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1144), .B1(G171), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1047), .A2(new_n1064), .A3(new_n1069), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1073), .B(G301), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT54), .B1(new_n1078), .B2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1142), .A2(new_n1156), .A3(new_n1100), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1100), .A2(KEYINPUT62), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1153), .A2(new_n1078), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1158), .A2(KEYINPUT126), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  AOI211_X1 g736(.A(G1976), .B(G288), .C1(new_n1027), .C2(new_n1031), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1024), .B1(new_n1162), .B2(new_n1030), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1040), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1163), .B1(new_n1166), .B2(new_n1069), .ZN(new_n1167));
  OAI21_X1  g742(.A(G8), .B1(new_n1068), .B2(new_n1062), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1053), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT121), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1069), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1092), .A2(G8), .A3(G168), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1047), .A2(new_n1176), .A3(new_n1169), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1171), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1174), .B1(new_n1153), .B2(new_n1173), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1167), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1102), .A2(new_n1157), .A3(new_n1161), .A4(new_n1180), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1146), .A2(new_n1059), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1035), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n1130), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1185), .A2(new_n879), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT116), .ZN(new_n1187));
  INV_X1    g762(.A(new_n750), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n748), .A2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n748), .A2(new_n1188), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1184), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n790), .B(new_n793), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1192), .B1(new_n1130), .B2(new_n766), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1184), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1187), .A2(new_n1191), .A3(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(G290), .A2(G1986), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(G290), .A2(G1986), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1183), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1181), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1187), .A2(new_n1190), .A3(new_n1194), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n791), .A2(new_n793), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1183), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1183), .B1(new_n766), .B2(new_n1192), .ZN(new_n1205));
  OR2_X1    g780(.A1(new_n1185), .A2(KEYINPUT46), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1185), .A2(KEYINPUT46), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT47), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1184), .A2(new_n1196), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT48), .ZN(new_n1211));
  AND4_X1   g786(.A1(new_n1191), .A2(new_n1187), .A3(new_n1194), .A4(new_n1211), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1204), .A2(new_n1209), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1201), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g789(.A1(new_n923), .A2(new_n925), .ZN(new_n1216));
  NOR2_X1   g790(.A1(G227), .A2(new_n460), .ZN(new_n1217));
  NAND2_X1  g791(.A1(new_n1217), .A2(new_n721), .ZN(new_n1218));
  NOR2_X1   g792(.A1(G401), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n1220));
  XNOR2_X1  g794(.A(new_n1219), .B(new_n1220), .ZN(new_n1221));
  AND3_X1   g795(.A1(new_n1216), .A2(new_n1006), .A3(new_n1221), .ZN(G308));
  NAND3_X1  g796(.A1(new_n1216), .A2(new_n1006), .A3(new_n1221), .ZN(G225));
endmodule


