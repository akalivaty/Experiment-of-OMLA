

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U322 ( .A(n383), .B(n382), .Z(n579) );
  AND2_X1 U323 ( .A1(G231GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U324 ( .A(KEYINPUT112), .B(KEYINPUT47), .ZN(n386) );
  XNOR2_X1 U325 ( .A(n439), .B(n290), .ZN(n377) );
  XNOR2_X1 U326 ( .A(n387), .B(n386), .ZN(n392) );
  XNOR2_X1 U327 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U328 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n393) );
  XNOR2_X1 U329 ( .A(n394), .B(n393), .ZN(n540) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n446) );
  XNOR2_X1 U331 ( .A(n446), .B(KEYINPUT58), .ZN(n447) );
  XNOR2_X1 U332 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(G50GAT), .B(G162GAT), .Z(n414) );
  XOR2_X1 U334 ( .A(G36GAT), .B(G190GAT), .Z(n395) );
  XOR2_X1 U335 ( .A(G99GAT), .B(G85GAT), .Z(n354) );
  INV_X1 U336 ( .A(n354), .ZN(n291) );
  NAND2_X1 U337 ( .A1(n395), .A2(n291), .ZN(n294) );
  INV_X1 U338 ( .A(n395), .ZN(n292) );
  NAND2_X1 U339 ( .A1(n292), .A2(n354), .ZN(n293) );
  NAND2_X1 U340 ( .A1(n294), .A2(n293), .ZN(n296) );
  NAND2_X1 U341 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n414), .B(n297), .ZN(n305) );
  XOR2_X1 U344 ( .A(KEYINPUT77), .B(KEYINPUT65), .Z(n299) );
  XNOR2_X1 U345 ( .A(G218GAT), .B(KEYINPUT76), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U347 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n301) );
  XNOR2_X1 U348 ( .A(KEYINPUT9), .B(KEYINPUT10), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U350 ( .A(n303), .B(n302), .Z(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U352 ( .A(KEYINPUT75), .B(G92GAT), .Z(n307) );
  XNOR2_X1 U353 ( .A(G134GAT), .B(G106GAT), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U356 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n311) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(G29GAT), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U359 ( .A(KEYINPUT68), .B(n312), .ZN(n347) );
  XOR2_X1 U360 ( .A(n313), .B(n347), .Z(n553) );
  INV_X1 U361 ( .A(KEYINPUT55), .ZN(n429) );
  XOR2_X1 U362 ( .A(G57GAT), .B(KEYINPUT4), .Z(n315) );
  XNOR2_X1 U363 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n334) );
  XOR2_X1 U365 ( .A(G148GAT), .B(G162GAT), .Z(n317) );
  XNOR2_X1 U366 ( .A(G127GAT), .B(G155GAT), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U368 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n319) );
  XNOR2_X1 U369 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U371 ( .A(n321), .B(n320), .Z(n327) );
  XNOR2_X1 U372 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n322) );
  XNOR2_X1 U373 ( .A(n322), .B(KEYINPUT2), .ZN(n423) );
  XOR2_X1 U374 ( .A(G85GAT), .B(n423), .Z(n324) );
  NAND2_X1 U375 ( .A1(G225GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U377 ( .A(G29GAT), .B(n325), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U379 ( .A(n328), .B(KEYINPUT1), .Z(n332) );
  XOR2_X1 U380 ( .A(G120GAT), .B(KEYINPUT0), .Z(n330) );
  XNOR2_X1 U381 ( .A(G113GAT), .B(G134GAT), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n436) );
  XNOR2_X1 U383 ( .A(n436), .B(KEYINPUT6), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n334), .B(n333), .ZN(n512) );
  XOR2_X1 U386 ( .A(G169GAT), .B(G8GAT), .Z(n396) );
  XOR2_X1 U387 ( .A(G113GAT), .B(G15GAT), .Z(n336) );
  XNOR2_X1 U388 ( .A(G36GAT), .B(G50GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U390 ( .A(n396), .B(n337), .Z(n339) );
  NAND2_X1 U391 ( .A1(G229GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U393 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n341) );
  XNOR2_X1 U394 ( .A(KEYINPUT29), .B(KEYINPUT69), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U396 ( .A(n343), .B(n342), .Z(n349) );
  XOR2_X1 U397 ( .A(G1GAT), .B(G22GAT), .Z(n345) );
  XNOR2_X1 U398 ( .A(G141GAT), .B(G197GAT), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U400 ( .A(n347), .B(n346), .Z(n348) );
  XOR2_X1 U401 ( .A(n349), .B(n348), .Z(n498) );
  INV_X1 U402 ( .A(n498), .ZN(n571) );
  XOR2_X1 U403 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n351) );
  XNOR2_X1 U404 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n367) );
  XOR2_X1 U406 ( .A(G64GAT), .B(G92GAT), .Z(n353) );
  XNOR2_X1 U407 ( .A(G176GAT), .B(G204GAT), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n409) );
  XOR2_X1 U409 ( .A(n409), .B(n354), .Z(n356) );
  NAND2_X1 U410 ( .A1(G230GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U412 ( .A(KEYINPUT73), .B(KEYINPUT71), .Z(n358) );
  XNOR2_X1 U413 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n357) );
  XOR2_X1 U414 ( .A(n358), .B(n357), .Z(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n365) );
  XNOR2_X1 U416 ( .A(G106GAT), .B(G78GAT), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n361), .B(G148GAT), .ZN(n415) );
  XOR2_X1 U418 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n363) );
  XNOR2_X1 U419 ( .A(G71GAT), .B(G57GAT), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n378) );
  XNOR2_X1 U421 ( .A(n415), .B(n378), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n574) );
  INV_X1 U424 ( .A(KEYINPUT41), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n574), .B(n368), .ZN(n544) );
  NOR2_X1 U426 ( .A1(n571), .A2(n544), .ZN(n370) );
  XNOR2_X1 U427 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n385) );
  XOR2_X1 U429 ( .A(KEYINPUT15), .B(G64GAT), .Z(n372) );
  XNOR2_X1 U430 ( .A(G1GAT), .B(G78GAT), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U432 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n374) );
  XNOR2_X1 U433 ( .A(G8GAT), .B(KEYINPUT14), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n376), .B(n375), .ZN(n383) );
  XOR2_X1 U436 ( .A(G15GAT), .B(G127GAT), .Z(n439) );
  XOR2_X1 U437 ( .A(G22GAT), .B(G155GAT), .Z(n412) );
  XOR2_X1 U438 ( .A(n379), .B(n412), .Z(n381) );
  XNOR2_X1 U439 ( .A(G183GAT), .B(G211GAT), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n382) );
  AND2_X1 U441 ( .A1(n553), .A2(n579), .ZN(n384) );
  NAND2_X1 U442 ( .A1(n385), .A2(n384), .ZN(n387) );
  INV_X1 U443 ( .A(n553), .ZN(n463) );
  XOR2_X1 U444 ( .A(KEYINPUT36), .B(n463), .Z(n581) );
  NOR2_X1 U445 ( .A1(n581), .A2(n579), .ZN(n388) );
  XNOR2_X1 U446 ( .A(KEYINPUT45), .B(n388), .ZN(n389) );
  NAND2_X1 U447 ( .A1(n389), .A2(n571), .ZN(n390) );
  INV_X1 U448 ( .A(n574), .ZN(n467) );
  NOR2_X1 U449 ( .A1(n390), .A2(n467), .ZN(n391) );
  NOR2_X1 U450 ( .A1(n392), .A2(n391), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n407) );
  XOR2_X1 U452 ( .A(KEYINPUT89), .B(KEYINPUT87), .Z(n398) );
  NAND2_X1 U453 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U455 ( .A(n399), .B(KEYINPUT88), .Z(n405) );
  XOR2_X1 U456 ( .A(G183GAT), .B(KEYINPUT17), .Z(n401) );
  XNOR2_X1 U457 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n434) );
  XOR2_X1 U459 ( .A(G211GAT), .B(KEYINPUT21), .Z(n403) );
  XNOR2_X1 U460 ( .A(G197GAT), .B(G218GAT), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n422) );
  XNOR2_X1 U462 ( .A(n434), .B(n422), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U465 ( .A(n409), .B(n408), .Z(n488) );
  INV_X1 U466 ( .A(n488), .ZN(n514) );
  NOR2_X1 U467 ( .A1(n540), .A2(n514), .ZN(n410) );
  XNOR2_X1 U468 ( .A(KEYINPUT54), .B(n410), .ZN(n411) );
  AND2_X1 U469 ( .A1(n512), .A2(n411), .ZN(n569) );
  XNOR2_X1 U470 ( .A(KEYINPUT23), .B(KEYINPUT82), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n427) );
  XOR2_X1 U472 ( .A(n415), .B(n414), .Z(n417) );
  NAND2_X1 U473 ( .A1(G228GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U475 ( .A(G204GAT), .B(KEYINPUT81), .Z(n419) );
  XNOR2_X1 U476 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U478 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n460) );
  NAND2_X1 U482 ( .A1(n569), .A2(n460), .ZN(n428) );
  XOR2_X1 U483 ( .A(n429), .B(n428), .Z(n445) );
  XOR2_X1 U484 ( .A(KEYINPUT80), .B(KEYINPUT20), .Z(n431) );
  XNOR2_X1 U485 ( .A(G190GAT), .B(KEYINPUT79), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n444) );
  XOR2_X1 U487 ( .A(G71GAT), .B(G176GAT), .Z(n433) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U490 ( .A(n435), .B(n434), .Z(n438) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U493 ( .A(n440), .B(n439), .Z(n442) );
  XNOR2_X1 U494 ( .A(G43GAT), .B(G99GAT), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n518) );
  INV_X1 U497 ( .A(n518), .ZN(n528) );
  NAND2_X1 U498 ( .A1(n445), .A2(n528), .ZN(n562) );
  NOR2_X1 U499 ( .A1(n553), .A2(n562), .ZN(n448) );
  NAND2_X1 U500 ( .A1(n488), .A2(n528), .ZN(n449) );
  NAND2_X1 U501 ( .A1(n449), .A2(n460), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n450), .B(KEYINPUT92), .ZN(n451) );
  XOR2_X1 U503 ( .A(KEYINPUT25), .B(n451), .Z(n455) );
  XOR2_X1 U504 ( .A(KEYINPUT27), .B(KEYINPUT90), .Z(n452) );
  XOR2_X1 U505 ( .A(n488), .B(n452), .Z(n458) );
  NOR2_X1 U506 ( .A1(n460), .A2(n528), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n453), .B(KEYINPUT26), .ZN(n568) );
  NAND2_X1 U508 ( .A1(n458), .A2(n568), .ZN(n454) );
  NAND2_X1 U509 ( .A1(n455), .A2(n454), .ZN(n456) );
  NAND2_X1 U510 ( .A1(n512), .A2(n456), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n457), .B(KEYINPUT93), .ZN(n462) );
  INV_X1 U512 ( .A(n512), .ZN(n485) );
  NAND2_X1 U513 ( .A1(n458), .A2(n485), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n459), .B(KEYINPUT91), .ZN(n539) );
  XOR2_X1 U515 ( .A(KEYINPUT28), .B(n460), .Z(n493) );
  INV_X1 U516 ( .A(n493), .ZN(n522) );
  NAND2_X1 U517 ( .A1(n539), .A2(n522), .ZN(n526) );
  NOR2_X1 U518 ( .A1(n526), .A2(n528), .ZN(n461) );
  NOR2_X1 U519 ( .A1(n462), .A2(n461), .ZN(n479) );
  NOR2_X1 U520 ( .A1(n463), .A2(n579), .ZN(n464) );
  XOR2_X1 U521 ( .A(KEYINPUT16), .B(n464), .Z(n465) );
  NOR2_X1 U522 ( .A1(n479), .A2(n465), .ZN(n466) );
  XNOR2_X1 U523 ( .A(KEYINPUT94), .B(n466), .ZN(n500) );
  NOR2_X1 U524 ( .A1(n571), .A2(n467), .ZN(n483) );
  NAND2_X1 U525 ( .A1(n500), .A2(n483), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n468), .B(KEYINPUT95), .ZN(n477) );
  NAND2_X1 U527 ( .A1(n477), .A2(n485), .ZN(n472) );
  XOR2_X1 U528 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n470) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U532 ( .A(KEYINPUT96), .B(n473), .ZN(G1324GAT) );
  NAND2_X1 U533 ( .A1(n477), .A2(n488), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U535 ( .A(G15GAT), .B(KEYINPUT35), .Z(n476) );
  NAND2_X1 U536 ( .A1(n477), .A2(n528), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(G1326GAT) );
  NAND2_X1 U538 ( .A1(n493), .A2(n477), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n478), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U540 ( .A(G29GAT), .B(KEYINPUT39), .Z(n487) );
  XOR2_X1 U541 ( .A(KEYINPUT37), .B(KEYINPUT99), .Z(n482) );
  NOR2_X1 U542 ( .A1(n479), .A2(n581), .ZN(n480) );
  NAND2_X1 U543 ( .A1(n480), .A2(n579), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n482), .B(n481), .ZN(n511) );
  NAND2_X1 U545 ( .A1(n511), .A2(n483), .ZN(n484) );
  XOR2_X1 U546 ( .A(KEYINPUT38), .B(n484), .Z(n494) );
  NAND2_X1 U547 ( .A1(n485), .A2(n494), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(G1328GAT) );
  NAND2_X1 U549 ( .A1(n494), .A2(n488), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT100), .B(KEYINPUT40), .Z(n491) );
  NAND2_X1 U552 ( .A1(n528), .A2(n494), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U554 ( .A(G43GAT), .B(n492), .Z(G1330GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n496) );
  NAND2_X1 U556 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U558 ( .A(G50GAT), .B(n497), .ZN(G1331GAT) );
  XNOR2_X1 U559 ( .A(KEYINPUT104), .B(n544), .ZN(n557) );
  NOR2_X1 U560 ( .A1(n557), .A2(n498), .ZN(n499) );
  XOR2_X1 U561 ( .A(KEYINPUT105), .B(n499), .Z(n510) );
  NAND2_X1 U562 ( .A1(n510), .A2(n500), .ZN(n506) );
  NOR2_X1 U563 ( .A1(n512), .A2(n506), .ZN(n502) );
  XNOR2_X1 U564 ( .A(KEYINPUT103), .B(KEYINPUT42), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U567 ( .A1(n514), .A2(n506), .ZN(n504) );
  XOR2_X1 U568 ( .A(G64GAT), .B(n504), .Z(G1333GAT) );
  NOR2_X1 U569 ( .A1(n518), .A2(n506), .ZN(n505) );
  XOR2_X1 U570 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  NOR2_X1 U571 ( .A1(n522), .A2(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n511), .A2(n510), .ZN(n521) );
  NOR2_X1 U576 ( .A1(n512), .A2(n521), .ZN(n513) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U578 ( .A1(n514), .A2(n521), .ZN(n516) );
  XNOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n521), .ZN(n520) );
  XNOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1338GAT) );
  NOR2_X1 U585 ( .A1(n522), .A2(n521), .ZN(n524) );
  XNOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U588 ( .A(G106GAT), .B(n525), .Z(G1339GAT) );
  NOR2_X1 U589 ( .A1(n540), .A2(n526), .ZN(n527) );
  NAND2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n535) );
  NOR2_X1 U591 ( .A1(n571), .A2(n535), .ZN(n530) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n530), .B(n529), .ZN(G1340GAT) );
  NOR2_X1 U594 ( .A1(n557), .A2(n535), .ZN(n532) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NOR2_X1 U597 ( .A1(n579), .A2(n535), .ZN(n533) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(n533), .Z(n534) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  NOR2_X1 U600 ( .A1(n553), .A2(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(KEYINPUT51), .B(KEYINPUT114), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n539), .A2(n568), .ZN(n541) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n542), .B(KEYINPUT115), .ZN(n552) );
  NOR2_X1 U607 ( .A1(n571), .A2(n552), .ZN(n543) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n543), .Z(G1344GAT) );
  NOR2_X1 U609 ( .A1(n544), .A2(n552), .ZN(n549) );
  XOR2_X1 U610 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n546) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(KEYINPUT116), .B(n547), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n579), .A2(n552), .ZN(n550) );
  XOR2_X1 U616 ( .A(KEYINPUT118), .B(n550), .Z(n551) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(n551), .ZN(G1346GAT) );
  NOR2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1347GAT) );
  NOR2_X1 U621 ( .A1(n571), .A2(n562), .ZN(n556) );
  XOR2_X1 U622 ( .A(G169GAT), .B(n556), .Z(G1348GAT) );
  XNOR2_X1 U623 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n561) );
  NOR2_X1 U624 ( .A1(n557), .A2(n562), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NOR2_X1 U628 ( .A1(n579), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1350GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n566) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(KEYINPUT123), .B(n567), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT122), .B(n570), .ZN(n582) );
  NOR2_X1 U637 ( .A1(n571), .A2(n582), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n582), .ZN(n578) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n582), .A2(n579), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

