//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n804, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT97), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  XOR2_X1   g004(.A(G15gat), .B(G22gat), .Z(new_n206));
  OAI22_X1  g005(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(KEYINPUT16), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n207), .B1(new_n205), .B2(new_n204), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(G8gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210));
  AND2_X1   g009(.A1(G71gat), .A2(G78gat), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n211), .A2(KEYINPUT9), .ZN(new_n212));
  XOR2_X1   g011(.A(G57gat), .B(G64gat), .Z(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G71gat), .B(G78gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n209), .B1(new_n210), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(new_n220), .B(G183gat), .Z(new_n221));
  XNOR2_X1  g020(.A(G127gat), .B(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n220), .B(G183gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n222), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n219), .A2(new_n210), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(KEYINPUT99), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT100), .B(G211gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n233));
  NAND2_X1  g032(.A1(G231gat), .A2(G233gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n231), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n224), .A2(new_n236), .A3(new_n226), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n232), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n235), .B1(new_n232), .B2(new_n237), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(G134gat), .B(G162gat), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT101), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n242), .B(new_n243), .Z(new_n244));
  NAND2_X1  g043(.A1(G99gat), .A2(G106gat), .ZN(new_n245));
  INV_X1    g044(.A(G85gat), .ZN(new_n246));
  INV_X1    g045(.A(G92gat), .ZN(new_n247));
  AOI22_X1  g046(.A1(KEYINPUT8), .A2(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(KEYINPUT102), .A2(G85gat), .A3(G92gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT7), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(KEYINPUT102), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(G99gat), .B(G106gat), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT17), .ZN(new_n256));
  XNOR2_X1  g055(.A(G43gat), .B(G50gat), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT94), .B1(new_n257), .B2(KEYINPUT15), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(KEYINPUT15), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n258), .B(new_n259), .Z(new_n260));
  NOR2_X1   g059(.A1(G29gat), .A2(G36gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT14), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n262), .A2(KEYINPUT95), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(KEYINPUT95), .ZN(new_n264));
  XOR2_X1   g063(.A(KEYINPUT93), .B(G29gat), .Z(new_n265));
  INV_X1    g064(.A(G36gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n263), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT96), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n260), .A2(new_n268), .A3(KEYINPUT96), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(KEYINPUT15), .B(new_n257), .C1(new_n267), .C2(new_n262), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n256), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n274), .ZN(new_n276));
  AOI211_X1 g075(.A(KEYINPUT17), .B(new_n276), .C1(new_n271), .C2(new_n272), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n255), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(new_n274), .ZN(new_n280));
  INV_X1    g079(.A(new_n255), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G190gat), .B(G218gat), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n284), .B(KEYINPUT103), .Z(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AOI211_X1 g085(.A(KEYINPUT104), .B(new_n244), .C1(new_n283), .C2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n286), .B2(new_n283), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n286), .A3(new_n244), .ZN(new_n289));
  INV_X1    g088(.A(new_n283), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n290), .B(new_n285), .C1(KEYINPUT104), .C2(new_n244), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n240), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G228gat), .A2(G233gat), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n295), .B(KEYINPUT83), .Z(new_n296));
  XNOR2_X1  g095(.A(G211gat), .B(G218gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT22), .ZN(new_n299));
  INV_X1    g098(.A(G211gat), .ZN(new_n300));
  INV_X1    g099(.A(G218gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n297), .A2(new_n298), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n297), .B1(new_n302), .B2(new_n298), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G148gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G141gat), .ZN(new_n308));
  INV_X1    g107(.A(G141gat), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n309), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT77), .B1(new_n309), .B2(G148gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT78), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(KEYINPUT78), .B(new_n308), .C1(new_n310), .C2(new_n311), .ZN(new_n315));
  NAND2_X1  g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  INV_X1    g115(.A(G155gat), .ZN(new_n317));
  INV_X1    g116(.A(G162gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(new_n319), .B2(KEYINPUT2), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n314), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  XNOR2_X1  g121(.A(G141gat), .B(G148gat), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n319), .B(new_n316), .C1(new_n323), .C2(KEYINPUT2), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n306), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n322), .B1(new_n305), .B2(KEYINPUT29), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n321), .A2(new_n324), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n296), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT84), .ZN(new_n332));
  OR3_X1    g131(.A1(new_n327), .A2(new_n330), .A3(new_n295), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT84), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n334), .B(new_n296), .C1(new_n327), .C2(new_n330), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G22gat), .ZN(new_n337));
  INV_X1    g136(.A(G22gat), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n332), .A2(new_n333), .A3(new_n338), .A4(new_n335), .ZN(new_n339));
  XOR2_X1   g138(.A(G78gat), .B(G106gat), .Z(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT31), .ZN(new_n341));
  INV_X1    g140(.A(G50gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n337), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT86), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT86), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n337), .A2(new_n346), .A3(new_n339), .A4(new_n343), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n337), .A2(new_n339), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n343), .B(KEYINPUT82), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT85), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT85), .ZN(new_n353));
  AOI211_X1 g152(.A(new_n353), .B(new_n350), .C1(new_n337), .C2(new_n339), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n348), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n359));
  NOR2_X1   g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT66), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT66), .ZN(new_n362));
  INV_X1    g161(.A(new_n360), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT65), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(KEYINPUT23), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT23), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT65), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n362), .B(new_n363), .C1(new_n365), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n360), .A2(KEYINPUT23), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n361), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(G183gat), .A2(G190gat), .ZN(new_n371));
  AND2_X1   g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(KEYINPUT24), .ZN(new_n373));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT24), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT64), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(KEYINPUT64), .A3(new_n375), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n373), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n358), .B1(new_n370), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT67), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(KEYINPUT67), .B(new_n358), .C1(new_n370), .C2(new_n382), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT69), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT24), .B1(new_n372), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n387), .B2(new_n372), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n358), .B1(new_n389), .B2(new_n373), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n361), .A2(new_n368), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n381), .B(KEYINPUT68), .Z(new_n392));
  NAND4_X1  g191(.A1(new_n390), .A2(new_n391), .A3(new_n369), .A4(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n385), .A2(new_n386), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT27), .B(G183gat), .ZN(new_n395));
  INV_X1    g194(.A(G190gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n397), .B(KEYINPUT28), .Z(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT71), .B(KEYINPUT26), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n381), .B1(new_n399), .B2(new_n363), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n363), .A2(KEYINPUT26), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT70), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n398), .B(new_n374), .C1(new_n400), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n394), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n357), .B1(new_n404), .B2(new_n326), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n356), .B1(new_n394), .B2(new_n403), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n305), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n357), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT29), .B1(new_n394), .B2(new_n403), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n408), .B(new_n306), .C1(new_n357), .C2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT89), .B(KEYINPUT37), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G8gat), .B(G36gat), .Z(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(G64gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(new_n247), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT89), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT37), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n407), .A2(new_n410), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT38), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT1), .ZN(new_n421));
  INV_X1    g220(.A(G113gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(G120gat), .ZN(new_n423));
  INV_X1    g222(.A(G120gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(G113gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n421), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT72), .B1(new_n423), .B2(new_n425), .ZN(new_n427));
  XNOR2_X1  g226(.A(G127gat), .B(G134gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XOR2_X1   g228(.A(G113gat), .B(G120gat), .Z(new_n430));
  XOR2_X1   g229(.A(G127gat), .B(G134gat), .Z(new_n431));
  OAI211_X1 g230(.A(new_n421), .B(new_n430), .C1(new_n431), .C2(KEYINPUT72), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n329), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n321), .A2(new_n433), .A3(new_n324), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438));
  OAI211_X1 g237(.A(KEYINPUT79), .B(KEYINPUT5), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT79), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n435), .B2(new_n436), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT5), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n322), .B1(new_n321), .B2(new_n324), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(new_n434), .A3(new_n325), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT4), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n436), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n321), .A2(new_n433), .A3(KEYINPUT4), .A4(new_n324), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n446), .A2(new_n438), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n439), .A2(new_n443), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT80), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n450), .B2(KEYINPUT5), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n325), .A2(new_n434), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n448), .B(new_n449), .C1(new_n454), .C2(new_n444), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n456), .A2(KEYINPUT80), .A3(new_n442), .A4(new_n438), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT0), .B(G57gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(G85gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(G1gat), .B(G29gat), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n459), .B(new_n460), .Z(new_n461));
  NAND4_X1  g260(.A1(new_n451), .A2(new_n453), .A3(new_n457), .A4(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n451), .A2(new_n453), .A3(new_n457), .ZN(new_n465));
  INV_X1    g264(.A(new_n461), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(KEYINPUT6), .A3(new_n466), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n420), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n407), .A2(new_n410), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n417), .A2(new_n418), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT38), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n415), .A4(new_n412), .ZN(new_n475));
  INV_X1    g274(.A(new_n415), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n407), .A2(new_n476), .A3(new_n410), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT76), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT76), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n407), .A2(new_n479), .A3(new_n410), .A4(new_n476), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n355), .B1(new_n470), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT30), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n478), .A2(new_n483), .A3(new_n480), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n476), .B1(new_n407), .B2(new_n410), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n407), .A2(new_n476), .A3(new_n410), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n486), .B2(KEYINPUT30), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT39), .ZN(new_n489));
  INV_X1    g288(.A(new_n438), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n455), .A2(KEYINPUT87), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT87), .B1(new_n455), .B2(new_n490), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n455), .A2(new_n490), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n455), .A2(KEYINPUT87), .A3(new_n490), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n489), .B1(new_n437), .B2(new_n438), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n493), .A2(new_n499), .A3(KEYINPUT40), .A4(new_n461), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n500), .A2(new_n467), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n493), .A2(new_n499), .A3(new_n461), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT40), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n503), .B1(new_n502), .B2(new_n504), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n488), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT90), .B1(new_n482), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n484), .A2(new_n487), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n510), .B(new_n501), .C1(new_n506), .C2(new_n505), .ZN(new_n511));
  INV_X1    g310(.A(new_n469), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n512), .B1(new_n467), .B2(new_n464), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n478), .A2(new_n480), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n513), .A2(new_n514), .A3(new_n475), .A4(new_n420), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT90), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n511), .A2(new_n515), .A3(new_n516), .A4(new_n355), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT34), .ZN(new_n519));
  INV_X1    g318(.A(G227gat), .ZN(new_n520));
  INV_X1    g319(.A(G233gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n434), .B1(new_n394), .B2(new_n403), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n394), .A2(new_n434), .A3(new_n403), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n519), .B1(new_n526), .B2(KEYINPUT75), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n394), .A2(new_n434), .A3(new_n403), .ZN(new_n528));
  INV_X1    g327(.A(new_n522), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n528), .A2(new_n523), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT73), .B1(new_n530), .B2(KEYINPUT33), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT74), .B(G15gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G43gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(G71gat), .B(G99gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n524), .A2(new_n522), .A3(new_n525), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(KEYINPUT32), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT73), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT33), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n531), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT75), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n536), .B(KEYINPUT32), .C1(new_n539), .C2(new_n535), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n542), .B1(new_n541), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n527), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n543), .ZN(new_n547));
  INV_X1    g346(.A(new_n542), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n550));
  INV_X1    g349(.A(new_n527), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n546), .A2(new_n552), .A3(KEYINPUT36), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT36), .B1(new_n546), .B2(new_n552), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n462), .A2(new_n463), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT81), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n467), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n469), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n355), .B1(new_n560), .B2(new_n488), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n518), .A2(new_n555), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT35), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n552), .ZN(new_n565));
  INV_X1    g364(.A(new_n513), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n565), .A2(new_n488), .A3(new_n355), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n349), .A2(new_n351), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n353), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n349), .A2(KEYINPUT85), .A3(new_n351), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n569), .A2(new_n570), .B1(new_n345), .B2(new_n347), .ZN(new_n571));
  AOI211_X1 g370(.A(new_n564), .B(new_n571), .C1(new_n546), .C2(new_n552), .ZN(new_n572));
  INV_X1    g371(.A(new_n560), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(new_n510), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n564), .A2(new_n567), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n294), .B1(new_n563), .B2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G113gat), .B(G141gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G169gat), .B(G197gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT12), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n209), .B1(new_n275), .B2(new_n277), .ZN(new_n584));
  INV_X1    g383(.A(new_n209), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n280), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT98), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(KEYINPUT18), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n280), .B(new_n585), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n587), .B(KEYINPUT13), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n590), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n584), .A2(new_n586), .A3(new_n587), .A4(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n583), .B1(new_n598), .B2(KEYINPUT92), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT92), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n600), .A3(new_n582), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT105), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n281), .A2(KEYINPUT10), .A3(new_n217), .A4(new_n218), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n255), .B(new_n219), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(KEYINPUT10), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n604), .A2(new_n603), .ZN(new_n607));
  INV_X1    g406(.A(G230gat), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n606), .B(new_n607), .C1(new_n608), .C2(new_n521), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n521), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(KEYINPUT106), .A3(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(KEYINPUT106), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615));
  INV_X1    g414(.A(G176gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(G204gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OR3_X1    g419(.A1(new_n614), .A2(KEYINPUT107), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n620), .B1(new_n614), .B2(KEYINPUT107), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n602), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n576), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(new_n560), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT108), .B(G1gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(G1324gat));
  INV_X1    g427(.A(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n510), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT16), .B(G8gat), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT42), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(new_n630), .B2(G8gat), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n631), .B1(KEYINPUT109), .B2(new_n633), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(KEYINPUT109), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n632), .A2(new_n634), .B1(new_n636), .B2(new_n637), .ZN(G1325gat));
  NOR3_X1   g437(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT110), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT110), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n544), .A2(new_n545), .A3(new_n527), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n551), .B1(new_n549), .B2(new_n550), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n546), .A2(new_n552), .A3(KEYINPUT36), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n629), .A2(G15gat), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(G15gat), .B1(new_n629), .B2(new_n565), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(G1326gat));
  NOR2_X1   g450(.A1(new_n625), .A2(new_n355), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT43), .B(G22gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  NAND2_X1  g453(.A1(new_n563), .A2(new_n575), .ZN(new_n655));
  INV_X1    g454(.A(new_n292), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n655), .A2(new_n624), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n240), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n265), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n659), .A2(new_n560), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT45), .Z(new_n662));
  INV_X1    g461(.A(KEYINPUT112), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n561), .B1(new_n509), .B2(new_n517), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(new_n639), .B2(new_n646), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n575), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n667), .A3(new_n656), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n292), .B1(new_n563), .B2(new_n575), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n623), .B(KEYINPUT111), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n671), .A2(new_n602), .A3(new_n240), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n663), .B1(new_n673), .B2(new_n560), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n670), .A2(KEYINPUT112), .A3(new_n573), .A4(new_n672), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n660), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n662), .A2(new_n676), .ZN(G1328gat));
  NOR3_X1   g476(.A1(new_n659), .A2(G36gat), .A3(new_n488), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT46), .ZN(new_n679));
  OAI21_X1  g478(.A(G36gat), .B1(new_n673), .B2(new_n488), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(G1329gat));
  NAND3_X1  g480(.A1(new_n670), .A2(G43gat), .A3(new_n672), .ZN(new_n682));
  INV_X1    g481(.A(new_n565), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n659), .A2(new_n683), .ZN(new_n684));
  OAI22_X1  g483(.A1(new_n682), .A2(new_n647), .B1(new_n684), .B2(G43gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT47), .ZN(G1330gat));
  AOI211_X1 g485(.A(KEYINPUT44), .B(new_n292), .C1(new_n665), .C2(new_n575), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n667), .B1(new_n655), .B2(new_n656), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n571), .B(new_n672), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT113), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n689), .A2(new_n690), .A3(G50gat), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n689), .B2(G50gat), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n657), .A2(new_n342), .A3(new_n658), .A4(new_n571), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT114), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n689), .A2(G50gat), .ZN(new_n697));
  AND4_X1   g496(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT48), .A4(new_n693), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT48), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n689), .B2(G50gat), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n696), .B1(new_n700), .B2(new_n693), .ZN(new_n701));
  OAI22_X1  g500(.A1(new_n695), .A2(KEYINPUT48), .B1(new_n698), .B2(new_n701), .ZN(G1331gat));
  INV_X1    g501(.A(new_n671), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n665), .B2(new_n575), .ZN(new_n704));
  INV_X1    g503(.A(new_n602), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n294), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n560), .B(KEYINPUT115), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT116), .B(G57gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1332gat));
  NOR2_X1   g510(.A1(new_n707), .A2(new_n488), .ZN(new_n712));
  NOR2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  AND2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n712), .B2(new_n713), .ZN(G1333gat));
  OAI21_X1  g515(.A(G71gat), .B1(new_n707), .B2(new_n647), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n565), .B(KEYINPUT117), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(G71gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n707), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g520(.A1(new_n707), .A2(new_n355), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g522(.A1(new_n705), .A2(new_n240), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n666), .A2(new_n656), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n727), .A2(new_n246), .A3(new_n573), .A4(new_n623), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n623), .B(new_n724), .C1(new_n687), .C2(new_n688), .ZN(new_n729));
  OAI21_X1  g528(.A(G85gat), .B1(new_n729), .B2(new_n560), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1336gat));
  NOR3_X1   g530(.A1(new_n703), .A2(G92gat), .A3(new_n488), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT52), .ZN(new_n734));
  OAI21_X1  g533(.A(G92gat), .B1(new_n729), .B2(new_n488), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n729), .A2(new_n488), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n725), .A2(new_n726), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n725), .A2(new_n726), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n738), .A2(new_n739), .B1(KEYINPUT118), .B2(new_n732), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n732), .A2(KEYINPUT118), .ZN(new_n741));
  AOI22_X1  g540(.A1(G92gat), .A2(new_n737), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n736), .B1(new_n742), .B2(new_n734), .ZN(G1337gat));
  NOR2_X1   g542(.A1(new_n683), .A2(G99gat), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n623), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G99gat), .B1(new_n729), .B2(new_n647), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(G1338gat));
  NOR2_X1   g546(.A1(new_n703), .A2(G106gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n727), .A2(new_n571), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G106gat), .B1(new_n729), .B2(new_n355), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT53), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n749), .A2(new_n753), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1339gat));
  NAND2_X1  g554(.A1(new_n614), .A2(new_n620), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n619), .B1(new_n609), .B2(KEYINPUT54), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT54), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n606), .A2(new_n607), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(new_n610), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n757), .B1(new_n609), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n756), .B1(new_n761), .B2(KEYINPUT55), .ZN(new_n762));
  INV_X1    g561(.A(new_n757), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n609), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(KEYINPUT55), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT119), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n761), .A2(KEYINPUT119), .A3(KEYINPUT55), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n762), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(new_n599), .A3(new_n601), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n598), .A2(new_n582), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n592), .A2(new_n593), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n587), .B1(new_n584), .B2(new_n586), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n581), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(new_n623), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n770), .A2(new_n292), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n769), .A2(new_n771), .A3(new_n774), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n656), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n658), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n623), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n293), .A2(new_n602), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT120), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT120), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n779), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n683), .A2(new_n571), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n560), .A2(new_n510), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G113gat), .B1(new_n790), .B2(new_n602), .ZN(new_n791));
  INV_X1    g590(.A(new_n708), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(KEYINPUT121), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n786), .A2(new_n787), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n708), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n797), .A2(new_n422), .A3(new_n488), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n791), .B1(new_n798), .B2(new_n602), .ZN(G1340gat));
  OAI21_X1  g598(.A(G120gat), .B1(new_n790), .B2(new_n703), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n488), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n623), .A2(new_n424), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(G1341gat));
  INV_X1    g602(.A(G127gat), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n790), .A2(new_n804), .A3(new_n658), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n797), .A2(new_n240), .A3(new_n488), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n804), .ZN(G1342gat));
  INV_X1    g606(.A(G134gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n656), .A2(new_n488), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT122), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n797), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT56), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n813), .A3(new_n808), .A4(new_n810), .ZN(new_n814));
  OAI21_X1  g613(.A(G134gat), .B1(new_n790), .B2(new_n292), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(G1343gat));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n355), .B1(new_n783), .B2(new_n785), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n648), .A2(new_n708), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n705), .A3(new_n488), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n821), .A2(new_n309), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n782), .A2(new_n571), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT57), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n647), .A2(new_n789), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n824), .A2(G141gat), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n602), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n817), .B1(new_n822), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n821), .A2(new_n309), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n831), .B(KEYINPUT58), .C1(new_n602), .C2(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1344gat));
  NAND3_X1  g632(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n780), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n835), .A2(KEYINPUT59), .A3(new_n307), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837));
  INV_X1    g636(.A(new_n785), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n784), .B1(new_n779), .B2(new_n781), .ZN(new_n839));
  OAI211_X1 g638(.A(KEYINPUT57), .B(new_n571), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n823), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT123), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n827), .A2(KEYINPUT123), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n842), .A2(new_n843), .A3(new_n623), .A4(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n837), .B1(new_n845), .B2(G148gat), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n820), .A2(new_n488), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n623), .A2(new_n307), .ZN(new_n848));
  OAI22_X1  g647(.A1(new_n836), .A2(new_n846), .B1(new_n847), .B2(new_n848), .ZN(G1345gat));
  NOR3_X1   g648(.A1(new_n834), .A2(new_n317), .A3(new_n658), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n820), .A2(new_n240), .A3(new_n488), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n317), .B2(new_n851), .ZN(G1346gat));
  OAI21_X1  g651(.A(G162gat), .B1(new_n834), .B2(new_n292), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n820), .A2(new_n318), .A3(new_n810), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1347gat));
  NOR2_X1   g654(.A1(new_n573), .A2(new_n488), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n786), .A2(new_n787), .A3(new_n856), .ZN(new_n857));
  OR3_X1    g656(.A1(new_n857), .A2(G169gat), .A3(new_n602), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n708), .A2(new_n510), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n718), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n786), .A2(new_n355), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G169gat), .B1(new_n861), .B2(new_n602), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n862), .ZN(G1348gat));
  INV_X1    g662(.A(new_n857), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n616), .A3(new_n623), .ZN(new_n865));
  OAI21_X1  g664(.A(G176gat), .B1(new_n861), .B2(new_n703), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT124), .ZN(G1349gat));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n240), .A3(new_n395), .ZN(new_n869));
  OAI21_X1  g668(.A(G183gat), .B1(new_n861), .B2(new_n658), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g671(.A1(new_n864), .A2(new_n396), .A3(new_n656), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT125), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n786), .A2(new_n656), .A3(new_n355), .A4(new_n860), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT126), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n876), .A3(G190gat), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n876), .B1(new_n875), .B2(G190gat), .ZN(new_n880));
  OR3_X1    g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n879), .B1(new_n878), .B2(new_n880), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n874), .A2(new_n881), .A3(new_n882), .ZN(G1351gat));
  AND3_X1   g682(.A1(new_n818), .A2(new_n647), .A3(new_n856), .ZN(new_n884));
  INV_X1    g683(.A(G197gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(new_n705), .ZN(new_n886));
  INV_X1    g685(.A(new_n842), .ZN(new_n887));
  INV_X1    g686(.A(new_n859), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n647), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n887), .A2(new_n602), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n890), .B2(new_n885), .ZN(G1352gat));
  NAND3_X1  g690(.A1(new_n884), .A2(new_n618), .A3(new_n623), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n892), .A2(KEYINPUT62), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(KEYINPUT62), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n887), .A2(new_n703), .A3(new_n889), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n893), .B(new_n894), .C1(new_n618), .C2(new_n895), .ZN(G1353gat));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n897));
  AOI211_X1 g696(.A(new_n658), .B(new_n889), .C1(new_n840), .C2(new_n841), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(new_n300), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n842), .A2(new_n240), .A3(new_n647), .A4(new_n888), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n901), .A3(KEYINPUT127), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n300), .A3(new_n240), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT127), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n904), .B(new_n897), .C1(new_n898), .C2(new_n300), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(G1354gat));
  NAND3_X1  g705(.A1(new_n884), .A2(new_n301), .A3(new_n656), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n887), .A2(new_n292), .A3(new_n889), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n301), .ZN(G1355gat));
endmodule


