//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT65), .B(G50), .ZN(new_n208));
  AND3_X1   g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT66), .B(G77), .Z(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G50), .ZN(new_n224));
  INV_X1    g0024(.A(G226), .ZN(new_n225));
  INV_X1    g0025(.A(G116), .ZN(new_n226));
  INV_X1    g0026(.A(G270), .ZN(new_n227));
  OAI22_X1  g0027(.A1(new_n224), .A2(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(G68), .B2(G238), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n221), .A2(new_n223), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n214), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT68), .Z(new_n234));
  NOR2_X1   g0034(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n206), .A2(new_n224), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(G1), .A2(G13), .ZN(new_n238));
  NOR3_X1   g0038(.A1(new_n237), .A2(new_n212), .A3(new_n238), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n214), .A2(G13), .ZN(new_n240));
  OAI211_X1 g0040(.A(new_n240), .B(G250), .C1(G257), .C2(G264), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(KEYINPUT0), .Z(new_n242));
  NOR4_X1   g0042(.A1(new_n234), .A2(new_n235), .A3(new_n239), .A4(new_n242), .ZN(G361));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  INV_X1    g0044(.A(G232), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT2), .B(G226), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G264), .B(G270), .Z(new_n249));
  XNOR2_X1  g0049(.A(G250), .B(G257), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G358));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT69), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(G68), .B(G77), .Z(new_n257));
  XNOR2_X1  g0057(.A(G50), .B(G58), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n256), .B(new_n259), .ZN(G351));
  INV_X1    g0060(.A(G200), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(G1), .B(G13), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G87), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT77), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT74), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n267), .A2(KEYINPUT74), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n225), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n266), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n273), .A2(G223), .A3(new_n274), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n264), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(new_n264), .A3(G274), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n264), .A2(new_n279), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(new_n245), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n261), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n238), .B1(G33), .B2(G41), .ZN(new_n285));
  INV_X1    g0085(.A(new_n266), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n267), .A2(KEYINPUT74), .A3(G33), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(new_n270), .ZN(new_n289));
  INV_X1    g0089(.A(new_n275), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n286), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G223), .ZN(new_n292));
  AOI211_X1 g0092(.A(new_n292), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n285), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  INV_X1    g0095(.A(new_n283), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n284), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n238), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n268), .A2(new_n269), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT7), .B1(new_n302), .B2(new_n212), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT7), .ZN(new_n304));
  AOI211_X1 g0104(.A(new_n304), .B(G20), .C1(new_n268), .C2(new_n269), .ZN(new_n305));
  OAI21_X1  g0105(.A(G68), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G58), .A2(G68), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n204), .A2(new_n205), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT75), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n212), .A2(new_n262), .ZN(new_n310));
  INV_X1    g0110(.A(G159), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G20), .A2(G33), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(KEYINPUT75), .A3(G159), .ZN(new_n314));
  AOI22_X1  g0114(.A1(G20), .A2(new_n308), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n306), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT16), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n301), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n271), .A2(new_n212), .A3(new_n272), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT7), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n271), .A2(new_n304), .A3(new_n212), .A4(new_n272), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(G68), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n308), .A2(G20), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n312), .A2(new_n314), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT76), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT76), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n322), .B(KEYINPUT16), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n318), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n300), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT8), .B(G58), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n211), .A2(G20), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n332), .A2(new_n336), .B1(new_n329), .B2(new_n334), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n298), .A2(new_n328), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT17), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n328), .A2(new_n338), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT18), .ZN(new_n343));
  OAI21_X1  g0143(.A(G169), .B1(new_n278), .B2(new_n283), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n294), .A2(G179), .A3(new_n296), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n344), .A2(new_n345), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n337), .B1(new_n318), .B2(new_n327), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT18), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(KEYINPUT17), .A3(new_n298), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n341), .A2(new_n347), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n212), .B1(new_n206), .B2(new_n208), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n262), .A2(G20), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G150), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n333), .A2(new_n356), .B1(new_n357), .B2(new_n310), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n300), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n224), .B1(new_n211), .B2(G20), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n331), .A2(new_n360), .B1(new_n224), .B2(new_n330), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT70), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n363), .B(KEYINPUT9), .ZN(new_n364));
  INV_X1    g0164(.A(G274), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n285), .A2(new_n365), .A3(new_n279), .ZN(new_n366));
  INV_X1    g0166(.A(new_n282), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n366), .B1(G226), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(G222), .A2(G1698), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n274), .A2(G223), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n288), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n371), .B(new_n285), .C1(new_n222), .C2(new_n288), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(new_n295), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(G200), .B2(new_n373), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n364), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT10), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT10), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n364), .A2(new_n378), .A3(new_n375), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n313), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n356), .B2(new_n207), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n300), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n383), .A2(KEYINPUT11), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(KEYINPUT11), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n331), .A2(G68), .A3(new_n335), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n329), .A2(G68), .B1(KEYINPUT73), .B2(KEYINPUT12), .ZN(new_n388));
  NAND2_X1  g0188(.A1(KEYINPUT73), .A2(KEYINPUT12), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n386), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n245), .A2(G1698), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n288), .B(new_n392), .C1(G226), .C2(G1698), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G97), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT71), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(KEYINPUT71), .A2(G33), .A3(G97), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n285), .ZN(new_n400));
  INV_X1    g0200(.A(G238), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n281), .B1(new_n282), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT13), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n400), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n264), .B1(new_n393), .B2(new_n398), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT13), .B1(new_n406), .B2(new_n402), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT14), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(G169), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(G179), .A3(new_n407), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n409), .B1(new_n408), .B2(G169), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n391), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n261), .B1(new_n405), .B2(new_n407), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT72), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n408), .B2(new_n295), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT72), .A4(G190), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n391), .B(new_n416), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n288), .A2(G232), .A3(new_n274), .ZN(new_n422));
  INV_X1    g0222(.A(G107), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n288), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n302), .A2(new_n401), .A3(new_n274), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n285), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n366), .B1(G244), .B2(new_n367), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G169), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XOR2_X1   g0230(.A(KEYINPUT15), .B(G87), .Z(new_n431));
  AOI22_X1  g0231(.A1(G20), .A2(new_n222), .B1(new_n431), .B2(new_n355), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n334), .A2(new_n313), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n301), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n331), .A2(G77), .A3(new_n335), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n222), .B2(new_n329), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n430), .B(new_n438), .C1(G179), .C2(new_n428), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n428), .A2(G200), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n440), .B(new_n437), .C1(new_n295), .C2(new_n428), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n373), .A2(new_n429), .ZN(new_n442));
  INV_X1    g0242(.A(G179), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n368), .A2(new_n443), .A3(new_n372), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n362), .A3(new_n444), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n439), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  AND4_X1   g0246(.A1(new_n353), .A2(new_n380), .A3(new_n421), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT23), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n212), .B2(G107), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n423), .A2(KEYINPUT23), .A3(G20), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G116), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT83), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(new_n212), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT83), .B1(new_n452), .B2(G20), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT84), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n451), .A2(new_n455), .A3(KEYINPUT84), .A4(new_n456), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT24), .ZN(new_n462));
  AOI21_X1  g0262(.A(G20), .B1(new_n271), .B2(new_n272), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT22), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(new_n216), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n288), .A2(new_n212), .A3(G87), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n463), .A2(new_n465), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n461), .A2(new_n462), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n462), .B1(new_n461), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n300), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT25), .B1(new_n330), .B2(new_n423), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n330), .A2(KEYINPUT25), .A3(new_n423), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n262), .A2(G1), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n330), .A2(new_n300), .A3(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n473), .A2(new_n474), .B1(new_n476), .B2(G107), .ZN(new_n477));
  INV_X1    g0277(.A(G45), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G1), .ZN(new_n479));
  AND2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  NOR2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G264), .A3(new_n264), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT85), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n482), .A2(KEYINPUT85), .A3(G264), .A4(new_n264), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n482), .A2(new_n285), .A3(new_n365), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n217), .A2(new_n274), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n219), .A2(G1698), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n271), .B2(new_n272), .ZN(new_n493));
  INV_X1    g0293(.A(G294), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n262), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n285), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n487), .A2(new_n489), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G190), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(G200), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n471), .A2(new_n477), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT81), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT19), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n503), .B(new_n212), .C1(new_n398), .C2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n396), .B2(new_n397), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT81), .B1(new_n506), .B2(G20), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n216), .A2(new_n218), .A3(new_n423), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT19), .B1(new_n355), .B2(G97), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n463), .B2(G68), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n300), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n431), .A2(new_n329), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n476), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n513), .B(new_n515), .C1(new_n216), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n401), .A2(new_n274), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(G244), .B2(new_n274), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n272), .B2(new_n271), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n285), .B1(new_n520), .B2(new_n453), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n285), .A2(new_n217), .A3(new_n479), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n285), .A2(new_n365), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n479), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n261), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(new_n524), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n295), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n301), .B1(new_n509), .B2(new_n511), .ZN(new_n529));
  INV_X1    g0329(.A(new_n431), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n516), .A2(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n529), .A2(new_n514), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n527), .A2(new_n429), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(G179), .B2(new_n527), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n517), .A2(new_n528), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n502), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n482), .A2(new_n264), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n489), .B1(new_n219), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n274), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n288), .A2(G250), .A3(G1698), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G283), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT79), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n273), .A2(new_n543), .A3(G244), .A4(new_n274), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT4), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(G1698), .B1(new_n271), .B2(new_n272), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n547), .B2(G244), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n542), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n538), .B1(new_n549), .B2(new_n285), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT80), .B1(new_n550), .B2(G190), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n303), .A2(new_n305), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(new_n423), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n313), .A2(G77), .ZN(new_n555));
  XNOR2_X1  g0355(.A(G97), .B(G107), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT78), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(KEYINPUT6), .ZN(new_n558));
  MUX2_X1   g0358(.A(new_n557), .B(G97), .S(KEYINPUT6), .Z(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n555), .B1(new_n560), .B2(new_n212), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n300), .B1(new_n554), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n329), .A2(G97), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n476), .B2(G97), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n550), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(G200), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n550), .A2(KEYINPUT80), .A3(G190), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n552), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n550), .A2(new_n443), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n570), .B(new_n565), .C1(G169), .C2(new_n550), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n536), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n498), .A2(new_n443), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n497), .A2(new_n429), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n471), .B2(new_n477), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT82), .B1(new_n537), .B2(new_n227), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT82), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n482), .A2(new_n578), .A3(G270), .A4(new_n264), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n219), .A2(new_n274), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(G264), .B2(new_n274), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n272), .B2(new_n271), .ZN(new_n583));
  INV_X1    g0383(.A(G303), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n288), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n285), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n580), .A2(new_n489), .A3(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n541), .B(new_n212), .C1(G33), .C2(new_n218), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(new_n300), .C1(new_n212), .C2(G116), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT20), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n329), .A2(G116), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n476), .B2(G116), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n587), .A2(new_n594), .A3(G169), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n587), .A2(new_n594), .A3(KEYINPUT21), .A4(G169), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n580), .A2(new_n586), .A3(G179), .A4(new_n489), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n594), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n597), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n576), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n594), .B1(new_n587), .B2(G200), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n295), .B2(new_n587), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n447), .A2(new_n572), .A3(new_n606), .ZN(G372));
  NOR2_X1   g0407(.A1(new_n532), .A2(new_n534), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT26), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n571), .B2(new_n535), .ZN(new_n610));
  INV_X1    g0410(.A(new_n534), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n513), .B(new_n515), .C1(new_n516), .C2(new_n530), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n516), .A2(new_n216), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n529), .A2(new_n514), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n527), .A2(new_n295), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(new_n525), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n611), .A2(new_n612), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n562), .A2(new_n564), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n566), .B2(new_n429), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n617), .A2(new_n619), .A3(KEYINPUT26), .A4(new_n570), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n608), .B1(new_n610), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n536), .A2(new_n569), .A3(new_n571), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT86), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n576), .B2(new_n602), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n597), .A2(new_n598), .A3(new_n601), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n461), .A2(new_n467), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT24), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n301), .B1(new_n627), .B2(new_n468), .ZN(new_n628));
  INV_X1    g0428(.A(new_n477), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n574), .B(new_n573), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n625), .A2(new_n630), .A3(KEYINPUT86), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n621), .B1(new_n622), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n447), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n445), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT88), .ZN(new_n636));
  INV_X1    g0436(.A(new_n379), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n378), .B1(new_n364), .B2(new_n375), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n377), .A2(new_n379), .A3(KEYINPUT88), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n414), .B1(new_n420), .B2(new_n439), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n341), .A2(new_n351), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n347), .A2(new_n350), .A3(KEYINPUT87), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT87), .B1(new_n347), .B2(new_n350), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n635), .B1(new_n641), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n634), .A2(new_n649), .ZN(G369));
  NAND3_X1  g0450(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n594), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n625), .B(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(new_n605), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n630), .A2(new_n656), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n656), .B1(new_n628), .B2(new_n629), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n501), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n660), .B1(new_n630), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n659), .A2(G330), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n625), .A2(new_n656), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n660), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g0467(.A(new_n667), .B(KEYINPUT89), .Z(G399));
  INV_X1    g0468(.A(new_n240), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(G41), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n508), .A2(G116), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G1), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n237), .B2(new_n671), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT28), .ZN(new_n675));
  INV_X1    g0475(.A(new_n656), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n633), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT29), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(KEYINPUT92), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT92), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n618), .B1(new_n261), .B2(new_n550), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n551), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n682), .A2(new_n568), .B1(new_n570), .B2(new_n619), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n536), .A3(new_n624), .A4(new_n631), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n656), .B1(new_n684), .B2(new_n621), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n680), .B1(new_n685), .B2(KEYINPUT29), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n621), .B1(new_n622), .B2(new_n603), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .A3(new_n676), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n679), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n587), .A2(new_n443), .A3(new_n527), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT91), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n550), .B2(new_n498), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n273), .A2(G244), .A3(new_n274), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT79), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(new_n545), .A3(new_n544), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n264), .B1(new_n696), .B2(new_n542), .ZN(new_n697));
  OAI211_X1 g0497(.A(KEYINPUT91), .B(new_n497), .C1(new_n697), .C2(new_n538), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n691), .B1(new_n693), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n487), .A2(new_n521), .A3(new_n524), .A4(new_n496), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n599), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n550), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT90), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI211_X1 g0505(.A(KEYINPUT90), .B(KEYINPUT30), .C1(new_n550), .C2(new_n702), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n699), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT31), .B1(new_n707), .B2(new_n676), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT90), .B1(new_n550), .B2(new_n702), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(new_n700), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n709), .B(new_n656), .C1(new_n711), .C2(new_n699), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n572), .A2(new_n606), .A3(new_n676), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n690), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n689), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n675), .B1(new_n718), .B2(G1), .ZN(G364));
  AND2_X1   g0519(.A1(new_n212), .A2(G13), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n211), .B1(new_n720), .B2(G45), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n670), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n659), .B2(G330), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(G330), .B2(new_n659), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT93), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n238), .B1(G20), .B2(new_n429), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n295), .A2(G200), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n212), .B1(new_n729), .B2(new_n443), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n218), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n212), .A2(new_n443), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G200), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n295), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n288), .B1(new_n735), .B2(new_n224), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n733), .A2(G190), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n731), .B(new_n736), .C1(G68), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n732), .B(KEYINPUT96), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n729), .ZN(new_n740));
  INV_X1    g0540(.A(new_n222), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G190), .A2(G200), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI221_X1 g0544(.A(new_n738), .B1(new_n202), .B2(new_n740), .C1(new_n741), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n212), .A2(G179), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n742), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n311), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT32), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n746), .A2(G190), .A3(G200), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n746), .A2(new_n295), .A3(G200), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n749), .B1(new_n216), .B2(new_n750), .C1(new_n423), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n740), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G322), .A2(new_n753), .B1(new_n743), .B2(G311), .ZN(new_n754));
  INV_X1    g0554(.A(new_n737), .ZN(new_n755));
  XOR2_X1   g0555(.A(KEYINPUT33), .B(G317), .Z(new_n756));
  INV_X1    g0556(.A(G283), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n755), .A2(new_n756), .B1(new_n751), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n747), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n288), .B1(new_n759), .B2(G329), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(new_n584), .B2(new_n750), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n754), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n730), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n734), .A2(G326), .B1(new_n764), .B2(G294), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT97), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n745), .A2(new_n752), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n728), .B1(new_n767), .B2(KEYINPUT98), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(KEYINPUT98), .B2(new_n767), .ZN(new_n769));
  INV_X1    g0569(.A(new_n723), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n240), .A2(G355), .A3(new_n288), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n669), .A2(new_n273), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n478), .B2(new_n236), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n775), .A2(KEYINPUT94), .B1(new_n478), .B2(new_n259), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n775), .A2(KEYINPUT94), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n771), .B1(G116), .B2(new_n240), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n727), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT95), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n770), .B1(new_n778), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n781), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n769), .B(new_n785), .C1(new_n659), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n726), .A2(new_n787), .ZN(G396));
  NAND2_X1  g0588(.A1(new_n438), .A2(new_n656), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n439), .A2(new_n441), .A3(new_n789), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n790), .A2(KEYINPUT102), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(KEYINPUT102), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n439), .A2(new_n676), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  OR3_X1    g0594(.A1(new_n685), .A2(KEYINPUT103), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(KEYINPUT103), .B1(new_n685), .B2(new_n794), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n791), .A2(new_n792), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n685), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(new_n716), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n723), .B1(new_n799), .B2(new_n716), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n794), .A2(new_n780), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n728), .A2(new_n780), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT99), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n723), .B1(new_n804), .B2(G77), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n753), .A2(G143), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G137), .A2(new_n734), .B1(new_n737), .B2(G150), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(new_n311), .C2(new_n744), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n289), .B1(G132), .B2(new_n759), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT101), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n730), .A2(new_n202), .B1(new_n750), .B2(new_n224), .ZN(new_n813));
  INV_X1    g0613(.A(new_n751), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(G68), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n810), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n808), .A2(new_n809), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n302), .B1(new_n747), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n731), .B(new_n819), .C1(new_n743), .C2(G116), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n494), .B2(new_n740), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n751), .A2(new_n216), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G303), .B2(new_n734), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n755), .A2(KEYINPUT100), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n755), .A2(KEYINPUT100), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n823), .B1(new_n423), .B2(new_n750), .C1(new_n826), .C2(new_n757), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n816), .A2(new_n817), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n805), .B1(new_n828), .B2(new_n727), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G384));
  NOR3_X1   g0631(.A1(new_n238), .A2(new_n212), .A3(new_n226), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n560), .B(KEYINPUT104), .Z(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT35), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT36), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n236), .A2(new_n222), .A3(new_n307), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n208), .A2(G68), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n211), .B(G13), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n415), .A2(new_n676), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT107), .Z(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n349), .A2(new_n298), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n349), .A2(new_n654), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n328), .A2(new_n338), .B1(new_n344), .B2(new_n345), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n322), .B1(new_n326), .B2(new_n325), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n317), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(new_n300), .A3(new_n327), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n348), .B1(new_n338), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n654), .B1(new_n855), .B2(new_n338), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n856), .A2(new_n857), .A3(new_n846), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n852), .B1(new_n858), .B2(new_n849), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT106), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n352), .A2(new_n860), .A3(new_n857), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n860), .B1(new_n352), .B2(new_n857), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n859), .B(KEYINPUT38), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT87), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT18), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n343), .B1(new_n342), .B2(new_n346), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n347), .A2(new_n350), .A3(KEYINPUT87), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n643), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n847), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n339), .B(KEYINPUT87), .C1(new_n349), .C2(new_n654), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n851), .A2(new_n848), .B1(new_n872), .B2(KEYINPUT37), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n339), .B1(new_n349), .B2(new_n654), .ZN(new_n874));
  NOR4_X1   g0674(.A1(new_n874), .A2(KEYINPUT87), .A3(new_n849), .A4(new_n850), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT38), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g0677(.A(KEYINPUT108), .B(KEYINPUT39), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n864), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT39), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n881), .B1(new_n884), .B2(new_n863), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT109), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n352), .A2(new_n857), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT106), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n352), .A2(new_n860), .A3(new_n857), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n891), .B2(new_n859), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT39), .B1(new_n892), .B2(new_n864), .ZN(new_n893));
  INV_X1    g0693(.A(new_n847), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n647), .B2(new_n643), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n850), .B2(new_n874), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n848), .A2(new_n865), .A3(KEYINPUT37), .A4(new_n851), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n883), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(new_n863), .A3(new_n878), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT109), .B1(new_n893), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n845), .B1(new_n887), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n439), .A2(new_n656), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n685), .B2(new_n797), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n391), .A2(new_n656), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n413), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n411), .A3(new_n410), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n420), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n418), .A2(new_n419), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n391), .B1(G200), .B2(new_n408), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n414), .A2(new_n913), .A3(new_n906), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n910), .A2(KEYINPUT105), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT105), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n916), .B(new_n907), .C1(new_n420), .C2(new_n909), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n905), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n884), .A2(new_n863), .ZN(new_n920));
  INV_X1    g0720(.A(new_n647), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n919), .A2(new_n920), .B1(new_n921), .B2(new_n654), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n903), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n679), .A2(new_n686), .A3(new_n447), .A4(new_n688), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n649), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n923), .B(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n915), .A2(new_n794), .A3(new_n917), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n713), .B2(new_n714), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n892), .B2(new_n864), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n900), .B2(new_n863), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n929), .A2(new_n930), .B1(new_n931), .B2(new_n928), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n713), .A2(new_n714), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n933), .A2(new_n447), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n690), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n934), .B2(new_n932), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n926), .A2(new_n936), .B1(new_n211), .B2(new_n720), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT110), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n926), .A2(new_n936), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n937), .A2(KEYINPUT110), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n842), .B1(new_n940), .B2(new_n941), .ZN(G367));
  OAI221_X1 g0742(.A(new_n782), .B1(new_n240), .B2(new_n530), .C1(new_n773), .C2(new_n251), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT112), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n770), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n944), .B2(new_n943), .ZN(new_n946));
  INV_X1    g0746(.A(new_n750), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT46), .B1(new_n947), .B2(G116), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n743), .A2(G283), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n948), .B(new_n950), .C1(G303), .C2(new_n753), .ZN(new_n951));
  INV_X1    g0751(.A(new_n826), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(G294), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n735), .A2(new_n818), .B1(new_n423), .B2(new_n730), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G97), .B2(new_n814), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n947), .A2(KEYINPUT46), .A3(G116), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n273), .B(new_n956), .C1(G317), .C2(new_n759), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n951), .A2(new_n953), .A3(new_n955), .A4(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(G137), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n288), .B1(new_n747), .B2(new_n959), .C1(new_n202), .C2(new_n750), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(new_n753), .B2(G150), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n208), .B2(new_n744), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n764), .A2(G68), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n734), .A2(G143), .B1(new_n814), .B2(new_n222), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n826), .C2(new_n311), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n958), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n946), .B1(new_n967), .B2(new_n727), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n614), .A2(new_n676), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n535), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n608), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n781), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n569), .B(new_n571), .C1(new_n618), .C2(new_n676), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n619), .A2(new_n570), .A3(new_n656), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n666), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(KEYINPUT44), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n666), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n666), .A2(new_n976), .A3(KEYINPUT45), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT45), .B1(new_n666), .B2(new_n976), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n978), .A2(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(new_n664), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n659), .A2(G330), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT111), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n659), .A2(KEYINPUT111), .A3(G330), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n663), .A2(new_n665), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n663), .A2(new_n665), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n987), .A2(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n986), .B2(new_n985), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n717), .B1(new_n984), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n670), .B(KEYINPUT41), .Z(new_n997));
  OAI21_X1  g0797(.A(new_n721), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n974), .A2(new_n630), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n656), .B1(new_n1000), .B2(new_n571), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n976), .A2(new_n663), .A3(new_n665), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1001), .B1(new_n1002), .B2(KEYINPUT42), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1002), .A2(KEYINPUT42), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n971), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1003), .A2(new_n1004), .B1(KEYINPUT43), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(KEYINPUT43), .B2(new_n1005), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT43), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1003), .A2(new_n1008), .A3(new_n971), .A4(new_n1004), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n976), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1010), .B1(new_n664), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n664), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1007), .A2(new_n1013), .A3(new_n976), .A4(new_n1009), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n973), .B1(new_n999), .B2(new_n1015), .ZN(G387));
  AOI22_X1  g0816(.A1(new_n743), .A2(G303), .B1(G322), .B2(new_n734), .ZN(new_n1017));
  INV_X1    g0817(.A(G317), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1017), .B1(new_n1018), .B2(new_n740), .C1(new_n826), .C2(new_n818), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT48), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n764), .A2(G283), .B1(new_n947), .B2(G294), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT49), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n751), .A2(new_n226), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n273), .B(new_n1028), .C1(G326), .C2(new_n759), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n530), .A2(new_n730), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n755), .A2(new_n333), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(G159), .C2(new_n734), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n289), .B1(G150), .B2(new_n759), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n947), .A2(new_n222), .B1(new_n814), .B2(G97), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G50), .A2(new_n753), .B1(new_n743), .B2(G68), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n728), .B1(new_n1030), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n672), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1039), .A2(new_n240), .A3(new_n288), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(G107), .B2(new_n240), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n248), .A2(G45), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT113), .ZN(new_n1043));
  AOI211_X1 g0843(.A(G45), .B(new_n1039), .C1(G68), .C2(G77), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n333), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n773), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1041), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n723), .B1(new_n1048), .B2(new_n783), .ZN(new_n1049));
  OR3_X1    g0849(.A1(new_n1038), .A2(KEYINPUT114), .A3(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(KEYINPUT114), .B1(new_n1038), .B2(new_n1049), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n663), .C2(new_n786), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n670), .B1(new_n994), .B2(new_n717), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n994), .A2(new_n717), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1052), .B1(new_n721), .B2(new_n994), .C1(new_n1053), .C2(new_n1055), .ZN(G393));
  NAND2_X1  g0856(.A1(new_n1011), .A2(new_n781), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n256), .A2(new_n773), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n782), .B1(new_n218), .B2(new_n240), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n723), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n208), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n952), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n750), .A2(new_n203), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n822), .B(new_n1063), .C1(G77), .C2(new_n764), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n743), .A2(new_n334), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n289), .B1(G143), .B2(new_n759), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n740), .A2(new_n311), .B1(new_n357), .B2(new_n735), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT51), .Z(new_n1069));
  OAI22_X1  g0869(.A1(new_n730), .A2(new_n226), .B1(new_n750), .B2(new_n757), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n288), .B1(new_n759), .B2(G322), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n423), .B2(new_n751), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(G294), .C2(new_n743), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n584), .B2(new_n826), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n740), .A2(new_n818), .B1(new_n1018), .B2(new_n735), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1067), .A2(new_n1069), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1060), .B1(new_n1078), .B2(new_n727), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n984), .A2(new_n722), .B1(new_n1057), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n994), .A2(new_n717), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n984), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n670), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1081), .A2(new_n984), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1080), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT116), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(KEYINPUT116), .B(new_n1080), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(G390));
  INV_X1    g0889(.A(new_n918), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n715), .A2(new_n794), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1090), .B1(new_n715), .B2(new_n794), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n798), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n1091), .A2(new_n1092), .B1(new_n1093), .B2(new_n904), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n715), .A2(new_n794), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n918), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n715), .A2(new_n794), .A3(new_n1090), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n687), .A2(new_n676), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n904), .B1(new_n1098), .B2(new_n797), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1094), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n715), .A2(new_n447), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n924), .A2(new_n649), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n886), .B1(new_n880), .B2(new_n885), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n893), .A2(new_n901), .A3(KEYINPUT109), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n844), .B1(new_n905), .B2(new_n918), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n844), .B1(new_n864), .B2(new_n877), .C1(new_n1099), .C2(new_n918), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1108), .A2(new_n1097), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1097), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1104), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1091), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1108), .A2(new_n1097), .A3(new_n1109), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n924), .A2(new_n649), .A3(new_n1102), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n1094), .B2(new_n1100), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1112), .A2(new_n1118), .A3(new_n670), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1105), .A2(new_n779), .A3(new_n1106), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n723), .B1(new_n804), .B2(new_n334), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT53), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n750), .B2(new_n357), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n947), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n952), .A2(G137), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT54), .B(G143), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G132), .A2(new_n753), .B1(new_n743), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n302), .B1(new_n759), .B2(G125), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n208), .B2(new_n751), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n734), .A2(G128), .B1(new_n764), .B2(G159), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1125), .A2(new_n1128), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT117), .Z(new_n1134));
  AOI22_X1  g0934(.A1(new_n743), .A2(G97), .B1(G283), .B2(new_n734), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n826), .B2(new_n423), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT118), .Z(new_n1137));
  OAI21_X1  g0937(.A(new_n302), .B1(new_n747), .B2(new_n494), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G87), .B2(new_n947), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n764), .A2(G77), .B1(new_n814), .B2(G68), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(new_n226), .C2(new_n740), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1134), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1121), .B1(new_n1142), .B2(new_n727), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1120), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n722), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1119), .A2(new_n1146), .ZN(G378));
  AOI21_X1  g0947(.A(new_n1116), .B1(new_n1145), .B2(new_n1101), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n929), .A2(new_n930), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n931), .A2(new_n928), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(G330), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n641), .A2(new_n445), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n362), .B(KEYINPUT70), .Z(new_n1153));
  NOR2_X1   g0953(.A1(new_n1153), .A2(new_n654), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1154), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n641), .A2(new_n445), .A3(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1158), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1156), .B1(new_n641), .B2(new_n445), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n635), .B(new_n1154), .C1(new_n639), .C2(new_n640), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1151), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n932), .A2(G330), .A3(new_n1166), .ZN(new_n1167));
  AND4_X1   g0967(.A1(new_n903), .A2(new_n1165), .A3(new_n922), .A4(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1167), .A2(new_n1165), .B1(new_n903), .B2(new_n922), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT57), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n670), .B1(new_n1148), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1118), .A2(new_n1103), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n923), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1165), .A2(new_n903), .A3(new_n1167), .A4(new_n922), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT57), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1171), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n721), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n751), .A2(new_n202), .B1(new_n747), .B2(new_n757), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n273), .A2(G41), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n741), .B2(new_n750), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1180), .B1(new_n1182), .B2(KEYINPUT119), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(KEYINPUT119), .B2(new_n1182), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT120), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n963), .B1(new_n755), .B2(new_n218), .C1(new_n226), .C2(new_n735), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n744), .A2(new_n530), .B1(new_n423), .B2(new_n740), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT58), .Z(new_n1189));
  AOI211_X1 g0989(.A(G50), .B(new_n1181), .C1(new_n262), .C2(new_n263), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G128), .A2(new_n753), .B1(new_n743), .B2(G137), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n750), .A2(new_n1126), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT121), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n734), .A2(G125), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n737), .A2(G132), .B1(new_n764), .B2(G150), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G33), .B(G41), .C1(new_n759), .C2(G124), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n311), .B2(new_n751), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1196), .B2(KEYINPUT59), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1190), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n728), .B1(new_n1189), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n723), .B1(new_n1061), .B2(new_n803), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(new_n1164), .C2(new_n779), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1178), .A2(new_n1179), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(G375));
  NAND2_X1  g1006(.A1(new_n1101), .A2(new_n722), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n723), .B1(new_n804), .B2(G68), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n734), .A2(G294), .B1(new_n947), .B2(G97), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n207), .B2(new_n751), .C1(new_n826), .C2(new_n226), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n302), .B1(new_n747), .B2(new_n584), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1031), .B(new_n1211), .C1(new_n743), .C2(G107), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n757), .B2(new_n740), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n289), .B1(G128), .B2(new_n759), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n959), .B2(new_n740), .C1(new_n744), .C2(new_n357), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n764), .A2(G50), .B1(new_n814), .B2(G58), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n734), .A2(G132), .B1(new_n947), .B2(G159), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n826), .C2(new_n1126), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1210), .A2(new_n1213), .B1(new_n1215), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1208), .B1(new_n1219), .B2(new_n727), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT122), .Z(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1090), .B2(new_n780), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1207), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n997), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1116), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1104), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1224), .A2(new_n1227), .ZN(G381));
  NOR2_X1   g1028(.A1(G393), .A2(G396), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n830), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(G390), .A2(new_n1230), .A3(G387), .A4(G381), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT123), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G378), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1119), .A2(new_n1146), .A3(KEYINPUT123), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1205), .A2(new_n1231), .A3(new_n1236), .ZN(G407));
  NAND2_X1  g1037(.A1(new_n1205), .A2(new_n1236), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G407), .B(G213), .C1(new_n1238), .C2(G343), .ZN(G409));
  AND2_X1   g1039(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1240), .A2(new_n998), .B1(new_n972), .B2(new_n968), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(G390), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(G387), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1243));
  AND2_X1   g1043(.A1(G393), .A2(G396), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(new_n1229), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1245), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1247), .A2(new_n1248), .A3(KEYINPUT127), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT127), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1245), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1250), .B1(new_n1253), .B2(new_n1246), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1249), .A2(new_n1254), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1110), .A2(new_n1111), .A3(new_n1104), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1176), .B(new_n1225), .C1(new_n1256), .C2(new_n1116), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1204), .B1(new_n1176), .B2(new_n722), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1233), .A2(new_n1234), .A3(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G378), .B(new_n1258), .C1(new_n1171), .C2(new_n1177), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n655), .A2(G213), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1104), .B2(new_n1226), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1226), .A2(new_n1264), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n670), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1224), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n830), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1226), .ZN(new_n1270));
  OAI21_X1  g1070(.A(KEYINPUT60), .B1(new_n1270), .B2(new_n1117), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n671), .B1(new_n1226), .B2(new_n1264), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(G384), .A3(new_n1224), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1269), .A2(new_n1274), .A3(KEYINPUT124), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT124), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  XOR2_X1   g1077(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1278));
  NAND4_X1  g1078(.A1(new_n1262), .A2(new_n1263), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT61), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1260), .A2(new_n1261), .B1(G213), .B2(new_n655), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT124), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G384), .B1(new_n1273), .B2(new_n1224), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n830), .B(new_n1223), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1269), .A2(new_n1274), .A3(KEYINPUT124), .ZN(new_n1286));
  INV_X1    g1086(.A(G2897), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1285), .B(new_n1286), .C1(new_n1287), .C2(new_n1263), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1269), .A2(new_n1274), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1289), .A2(G213), .A3(new_n655), .A4(G2897), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1279), .B(new_n1280), .C1(new_n1281), .C2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1293), .B1(new_n1281), .B2(new_n1277), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1255), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT61), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1281), .A2(new_n1277), .ZN(new_n1299));
  XOR2_X1   g1099(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1281), .A2(KEYINPUT63), .A3(new_n1277), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1298), .A2(new_n1301), .A3(new_n1302), .A4(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1295), .A2(new_n1304), .ZN(G405));
  OAI21_X1  g1105(.A(new_n1261), .B1(new_n1205), .B2(new_n1235), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1277), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1303), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1261), .B(new_n1289), .C1(new_n1205), .C2(new_n1235), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1308), .B1(new_n1307), .B2(new_n1309), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(G402));
endmodule


