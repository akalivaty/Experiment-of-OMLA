//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(G2106), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT68), .B(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n462), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(KEYINPUT3), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n470), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  AND4_X1   g049(.A1(KEYINPUT69), .A2(new_n472), .A3(new_n474), .A4(KEYINPUT3), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n463), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n467), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n472), .A2(new_n474), .A3(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(new_n470), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n472), .A2(new_n474), .A3(KEYINPUT69), .A4(KEYINPUT3), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(KEYINPUT70), .A3(G137), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n466), .B1(new_n478), .B2(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n483), .A2(G136), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n463), .B1(new_n481), .B2(new_n482), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT71), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n463), .A2(KEYINPUT72), .A3(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT73), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(new_n495), .C1(new_n498), .C2(new_n499), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n487), .A2(G126), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n505), .B1(new_n483), .B2(G138), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n505), .A2(KEYINPUT74), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(KEYINPUT74), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n463), .A2(G138), .ZN(new_n509));
  AND4_X1   g084(.A1(new_n464), .A2(new_n507), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  AND2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT75), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(new_n516), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n514), .B2(new_n513), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT76), .B(G88), .Z(new_n527));
  OAI22_X1  g102(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n519), .A2(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n513), .A2(new_n514), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n521), .A2(new_n522), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(G63), .A2(G651), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n535), .A2(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n533), .A2(new_n542), .B1(new_n526), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n525), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(G171));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n533), .A2(new_n548), .B1(new_n526), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n525), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT79), .ZN(new_n559));
  XNOR2_X1  g134(.A(KEYINPUT78), .B(KEYINPUT8), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n555), .A2(new_n561), .ZN(G188));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n533), .A2(KEYINPUT9), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n533), .B2(new_n563), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n536), .A2(new_n515), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n564), .A2(new_n565), .B1(G91), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n536), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n571), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(G651), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n567), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND2_X1  g152(.A1(new_n517), .A2(G49), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n532), .A2(G87), .A3(new_n523), .ZN(new_n579));
  INV_X1    g154(.A(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n521), .A2(new_n580), .A3(new_n522), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n581), .A2(KEYINPUT81), .A3(G651), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT81), .B1(new_n581), .B2(G651), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n578), .B(new_n579), .C1(new_n582), .C2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(new_n566), .A2(G86), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n521), .B2(new_n522), .ZN(new_n587));
  AND2_X1   g162(.A1(G73), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n532), .A2(G48), .A3(G543), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n566), .A2(G85), .B1(G47), .B2(new_n517), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n525), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT82), .ZN(G290));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(G301), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G54), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n598), .A2(new_n525), .B1(new_n533), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT83), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n566), .A2(G92), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT10), .Z(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT84), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n597), .B1(new_n606), .B2(new_n596), .ZN(G284));
  AOI21_X1  g182(.A(new_n597), .B1(new_n606), .B2(new_n596), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT85), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(G868), .B2(new_n611), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(G868), .B2(new_n611), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n606), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n606), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n461), .A2(new_n464), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n483), .A2(G135), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n487), .A2(G123), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT86), .B(G2096), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n623), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT88), .ZN(G401));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT89), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n649), .A3(new_n651), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n650), .A2(new_n651), .ZN(new_n659));
  INV_X1    g234(.A(new_n649), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n653), .B1(new_n660), .B2(new_n652), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT90), .B(G2096), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT91), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT93), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n673), .A2(new_n678), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT20), .Z(new_n681));
  NOR2_X1   g256(.A1(new_n674), .A2(new_n678), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT92), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n679), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT95), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT94), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1981), .B(G1986), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n685), .B(new_n691), .ZN(G229));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G22), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G166), .B2(new_n693), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(G1971), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(G1971), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT99), .ZN(new_n699));
  MUX2_X1   g274(.A(G6), .B(G305), .S(G16), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT32), .ZN(new_n701));
  INV_X1    g276(.A(G1981), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(G23), .B(G288), .S(G16), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT33), .B(G1976), .Z(new_n705));
  XOR2_X1   g280(.A(new_n704), .B(new_n705), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n698), .A2(KEYINPUT99), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n699), .A2(new_n703), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT34), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(KEYINPUT100), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  OR2_X1    g289(.A1(G95), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT96), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G119), .B2(new_n487), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n483), .A2(G131), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n714), .B1(new_n721), .B2(new_n713), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT97), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  MUX2_X1   g301(.A(G24), .B(G290), .S(G16), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT98), .ZN(new_n728));
  INV_X1    g303(.A(G1986), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n723), .A2(new_n725), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n729), .ZN(new_n732));
  AND4_X1   g307(.A1(new_n726), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n710), .A2(new_n712), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n693), .A2(G21), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G168), .B2(new_n693), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G1966), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT107), .Z(new_n738));
  INV_X1    g313(.A(G1956), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n693), .A2(G20), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT23), .Z(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G299), .B2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n738), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G5), .A2(G16), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT108), .Z(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G301), .B2(new_n693), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT109), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n742), .A2(new_n739), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n736), .A2(G1966), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n553), .A2(G16), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G16), .B2(G19), .ZN(new_n755));
  INV_X1    g330(.A(G1341), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n628), .A2(new_n713), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(G28), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n713), .B1(new_n759), .B2(G28), .ZN(new_n761));
  AND2_X1   g336(.A1(KEYINPUT31), .A2(G11), .ZN(new_n762));
  NOR2_X1   g337(.A1(KEYINPUT31), .A2(G11), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n755), .B2(new_n756), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n753), .A2(new_n757), .A3(new_n758), .A4(new_n765), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n743), .A2(new_n752), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G164), .A2(new_n713), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G27), .B2(new_n713), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n713), .B1(KEYINPUT24), .B2(G34), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(KEYINPUT24), .B2(G34), .ZN(new_n772));
  INV_X1    g347(.A(G160), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(G29), .ZN(new_n774));
  INV_X1    g349(.A(G2084), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n769), .A2(new_n770), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n767), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n713), .A2(G32), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n483), .A2(G141), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n487), .A2(G129), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT26), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n461), .A2(G105), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n779), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT105), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n778), .B1(new_n787), .B2(new_n713), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT27), .B(G1996), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT106), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n788), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n769), .A2(new_n770), .ZN(new_n792));
  INV_X1    g367(.A(G33), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n483), .A2(G139), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT102), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n464), .A2(G127), .ZN(new_n796));
  INV_X1    g371(.A(G115), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n469), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT101), .B(KEYINPUT25), .Z(new_n799));
  NAND3_X1  g374(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n798), .A2(G2105), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n795), .A2(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(new_n793), .B(new_n804), .S(G29), .Z(new_n805));
  INV_X1    g380(.A(G2072), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n792), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n713), .A2(G35), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT110), .Z(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n492), .B2(G29), .ZN(new_n810));
  INV_X1    g385(.A(G2090), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT111), .B(KEYINPUT29), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n713), .A2(G26), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT28), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n483), .A2(G140), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n487), .A2(G128), .ZN(new_n818));
  OR2_X1    g393(.A1(G104), .A2(G2105), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n819), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n816), .B1(new_n821), .B2(G29), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G2067), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n807), .A2(new_n814), .A3(new_n823), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n777), .A2(new_n791), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n774), .A2(new_n775), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT103), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n805), .A2(new_n806), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT104), .Z(new_n829));
  NOR2_X1   g404(.A1(G4), .A2(G16), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n606), .B2(G16), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G1348), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n825), .A2(new_n827), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n712), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n711), .A2(KEYINPUT100), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n710), .B2(new_n733), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n734), .A2(new_n834), .A3(new_n838), .ZN(G311));
  INV_X1    g414(.A(new_n838), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n825), .A2(new_n827), .A3(new_n833), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n710), .A2(new_n712), .A3(new_n733), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(G150));
  INV_X1    g418(.A(G55), .ZN(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n533), .A2(new_n844), .B1(new_n526), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT112), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(new_n525), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT114), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n606), .A2(G559), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n847), .A2(new_n553), .A3(new_n849), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n553), .B1(new_n847), .B2(new_n849), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n854), .B(KEYINPUT38), .ZN(new_n862));
  INV_X1    g437(.A(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n866));
  AOI21_X1  g441(.A(G860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT39), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n867), .A2(KEYINPUT113), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT113), .B1(new_n867), .B2(new_n868), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n853), .B1(new_n869), .B2(new_n870), .ZN(G145));
  NOR2_X1   g446(.A1(new_n804), .A2(new_n786), .ZN(new_n872));
  INV_X1    g447(.A(new_n787), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n804), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n720), .B(new_n621), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n483), .A2(G142), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n487), .A2(G130), .ZN(new_n877));
  OR2_X1    g452(.A1(G106), .A2(G2105), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n878), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g455(.A(G138), .B(new_n463), .C1(new_n471), .C2(new_n475), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n510), .B1(new_n881), .B2(KEYINPUT4), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n501), .A2(new_n503), .ZN(new_n883));
  OAI211_X1 g458(.A(G126), .B(G2105), .C1(new_n471), .C2(new_n475), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT115), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT115), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n504), .B(new_n887), .C1(new_n506), .C2(new_n510), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(new_n821), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n821), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n880), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n880), .A3(new_n891), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n875), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  INV_X1    g471(.A(new_n875), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n896), .A2(new_n897), .A3(new_n892), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n874), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n896), .B2(new_n892), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n893), .A2(new_n875), .A3(new_n894), .ZN(new_n901));
  INV_X1    g476(.A(new_n874), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(G162), .B(G160), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(new_n628), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n899), .A2(new_n906), .A3(new_n903), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g487(.A(KEYINPUT116), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n860), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT116), .B1(new_n858), .B2(new_n859), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n616), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n914), .A2(new_n614), .A3(new_n606), .A4(new_n915), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n605), .A2(new_n611), .ZN(new_n920));
  NAND3_X1  g495(.A1(G299), .A2(new_n602), .A3(new_n604), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(KEYINPUT117), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT117), .ZN(new_n923));
  NAND4_X1  g498(.A1(G299), .A2(new_n923), .A3(new_n602), .A4(new_n604), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n919), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(KEYINPUT41), .A3(new_n924), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n920), .A2(new_n929), .A3(new_n921), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n917), .A2(new_n931), .A3(new_n918), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n926), .A2(new_n927), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n927), .B1(new_n926), .B2(new_n932), .ZN(new_n935));
  XNOR2_X1  g510(.A(G290), .B(G305), .ZN(new_n936));
  XNOR2_X1  g511(.A(G166), .B(G288), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n936), .B(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n934), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n926), .A2(new_n932), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n938), .B1(new_n942), .B2(new_n933), .ZN(new_n943));
  OAI21_X1  g518(.A(G868), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n850), .A2(new_n596), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(G295));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n945), .ZN(G331));
  INV_X1    g522(.A(KEYINPUT118), .ZN(new_n948));
  OAI21_X1  g523(.A(G286), .B1(new_n948), .B2(G171), .ZN(new_n949));
  NAND2_X1  g524(.A1(G171), .A2(new_n948), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n858), .A2(new_n859), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n553), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n850), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n950), .B1(new_n954), .B2(new_n857), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n949), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n951), .B1(new_n858), .B2(new_n859), .ZN(new_n957));
  INV_X1    g532(.A(new_n949), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n857), .A3(new_n950), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n931), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n956), .A2(new_n925), .A3(new_n960), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n964), .B2(new_n939), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n929), .B1(new_n956), .B2(new_n960), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n920), .A2(new_n921), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n925), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n968), .B(new_n938), .C1(new_n969), .C2(new_n966), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n965), .A2(KEYINPUT43), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n963), .ZN(new_n972));
  AOI22_X1  g547(.A1(new_n956), .A2(new_n960), .B1(new_n928), .B2(new_n930), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT119), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT119), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n962), .A2(new_n975), .A3(new_n963), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n974), .A2(new_n976), .A3(new_n938), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT43), .B1(new_n977), .B2(new_n965), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT44), .B1(new_n971), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n965), .A2(new_n981), .A3(new_n970), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(new_n977), .B2(new_n965), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n984), .ZN(G397));
  INV_X1    g560(.A(G2067), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n821), .B(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n786), .A2(G1996), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n987), .B(new_n988), .C1(new_n873), .C2(G1996), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n720), .B(new_n725), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(G290), .B(new_n729), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n886), .A2(new_n888), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n466), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n476), .A2(new_n467), .A3(new_n477), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT70), .B1(new_n483), .B2(G137), .ZN(new_n1000));
  OAI211_X1 g575(.A(G40), .B(new_n998), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n993), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G286), .A2(G8), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT51), .B1(new_n1004), .B2(KEYINPUT124), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n994), .B1(new_n882), .B2(new_n885), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT50), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n511), .A2(new_n1009), .A3(new_n994), .ZN(new_n1010));
  INV_X1    g585(.A(G40), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n1011), .B(new_n466), .C1(new_n478), .C2(new_n484), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1008), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1007), .A2(new_n996), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n996), .A2(G1384), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n511), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1966), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1013), .A2(new_n775), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1004), .B(new_n1006), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1008), .A2(new_n1010), .A3(new_n775), .A4(new_n1012), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(G8), .B(new_n1005), .C1(new_n1024), .C2(G286), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(G8), .A3(G286), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1021), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT62), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(G160), .A2(new_n511), .A3(G40), .A4(new_n994), .ZN(new_n1033));
  OR2_X1    g608(.A1(G288), .A2(new_n1029), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(G8), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G305), .A2(G1981), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n585), .A2(new_n702), .A3(new_n589), .A4(new_n590), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1036), .A2(KEYINPUT49), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT49), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(new_n1033), .A3(G8), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1034), .B(G8), .C1(new_n1001), .C2(new_n1007), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1035), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n886), .A2(new_n888), .A3(new_n1015), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1046));
  INV_X1    g621(.A(G1971), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1008), .A2(new_n1010), .A3(new_n811), .A4(new_n1012), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1020), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(G8), .B1(new_n519), .B2(new_n528), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT55), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1044), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1001), .B1(new_n996), .B2(new_n1007), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1971), .B1(new_n1055), .B2(new_n1045), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1049), .ZN(new_n1057));
  OAI211_X1 g632(.A(G8), .B(new_n1053), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1061), .A2(KEYINPUT120), .A3(G8), .A4(new_n1053), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1054), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1045), .A2(new_n770), .A3(new_n1014), .A4(new_n1012), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1008), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n748), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1055), .A2(KEYINPUT53), .A3(new_n770), .A4(new_n1016), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT125), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT125), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1073), .A3(G171), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1021), .A2(new_n1025), .A3(new_n1076), .A4(new_n1026), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1028), .A2(new_n1063), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1060), .A2(new_n1062), .A3(new_n1044), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1033), .A2(G8), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AOI211_X1 g656(.A(G1976), .B(G288), .C1(new_n1081), .C2(new_n1040), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1037), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1079), .A2(new_n1084), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1019), .A2(new_n1020), .A3(G286), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT63), .B1(new_n1063), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1035), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1061), .A2(G8), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n1052), .ZN(new_n1091));
  AND4_X1   g666(.A1(KEYINPUT63), .A2(new_n1088), .A3(new_n1091), .A4(new_n1086), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1078), .B(new_n1085), .C1(new_n1087), .C2(new_n1092), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1001), .A2(new_n1065), .A3(G2078), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n997), .A2(new_n1045), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1066), .A2(new_n1068), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G171), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1066), .A2(G301), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(KEYINPUT54), .A3(new_n1098), .ZN(new_n1099));
  AND4_X1   g674(.A1(new_n1027), .A2(new_n1099), .A3(new_n1088), .A4(new_n1091), .ZN(new_n1100));
  INV_X1    g675(.A(G1348), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1067), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1033), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n986), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n606), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1067), .A2(new_n1101), .B1(new_n1103), .B2(new_n986), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1107), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1996), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1045), .A2(new_n1114), .A3(new_n1014), .A4(new_n1012), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(G1341), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1033), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1119), .A2(new_n553), .B1(KEYINPUT123), .B2(KEYINPUT59), .ZN(new_n1120));
  NAND2_X1  g695(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n953), .B(new_n1121), .C1(new_n1115), .C2(new_n1118), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1067), .A2(new_n739), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1055), .A2(new_n1045), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n1128));
  XNOR2_X1  g703(.A(G299), .B(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1129), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1124), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1129), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(KEYINPUT61), .A3(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1113), .A2(new_n1123), .A3(new_n1132), .A4(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1136), .B1(new_n1139), .B2(new_n1131), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1096), .A2(G171), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1072), .A2(new_n1074), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1100), .A2(new_n1141), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1003), .B1(new_n1093), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n721), .A2(new_n724), .ZN(new_n1148));
  OAI22_X1  g723(.A1(new_n989), .A2(new_n1148), .B1(G2067), .B2(new_n821), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1002), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1002), .ZN(new_n1151));
  OR3_X1    g726(.A1(new_n1151), .A2(G1986), .A3(G290), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT48), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1152), .A2(new_n1153), .B1(new_n1151), .B2(new_n991), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1150), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT46), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1151), .B2(G1996), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1158), .A2(KEYINPUT126), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(KEYINPUT126), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n786), .B1(KEYINPUT46), .B2(new_n1114), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n987), .A2(new_n1161), .ZN(new_n1162));
  OAI22_X1  g737(.A1(new_n1159), .A2(new_n1160), .B1(new_n1151), .B2(new_n1162), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1163), .A2(KEYINPUT47), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(KEYINPUT47), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1156), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1147), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g742(.A1(new_n667), .A2(new_n668), .A3(G319), .ZN(new_n1169));
  OR3_X1    g743(.A1(G401), .A2(KEYINPUT127), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g744(.A(KEYINPUT127), .B1(G401), .B2(new_n1169), .ZN(new_n1171));
  AOI21_X1  g745(.A(G229), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g746(.A(new_n911), .B(new_n1172), .C1(new_n982), .C2(new_n983), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


