//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  AND2_X1   g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n211), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n210), .B1(new_n220), .B2(KEYINPUT0), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n221), .B1(KEYINPUT0), .B2(new_n220), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT64), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G87), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n211), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  INV_X1    g0029(.A(G77), .ZN(new_n230));
  INV_X1    g0030(.A(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G107), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n229), .B1(new_n230), .B2(new_n231), .C1(new_n232), .C2(new_n219), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n215), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT1), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n223), .A2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT65), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  INV_X1    g0041(.A(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n240), .B(new_n245), .Z(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  INV_X1    g0047(.A(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT66), .B(G50), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  OR2_X1    g0055(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G97), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n262), .B1(new_n267), .B2(G232), .ZN(new_n268));
  OR2_X1    g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G226), .A3(new_n266), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n259), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(new_n259), .A3(G274), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n275), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n212), .A2(new_n278), .B1(new_n208), .B2(new_n258), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n280), .B2(new_n226), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n256), .B(new_n257), .C1(new_n273), .C2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n262), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n271), .A2(G1698), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n272), .B(new_n283), .C1(new_n284), .C2(new_n242), .ZN(new_n285));
  INV_X1    g0085(.A(new_n259), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n281), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n287), .A2(new_n288), .A3(KEYINPUT74), .A4(KEYINPUT13), .ZN(new_n289));
  AND2_X1   g0089(.A1(KEYINPUT76), .A2(G169), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n282), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT14), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT14), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n282), .A2(new_n293), .A3(new_n289), .A4(new_n290), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT13), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(KEYINPUT75), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n287), .A2(new_n288), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n296), .B1(new_n287), .B2(new_n288), .ZN(new_n298));
  OAI21_X1  g0098(.A(G179), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n292), .A2(new_n294), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n225), .A2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n213), .A2(G33), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G20), .A2(G33), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n301), .B1(new_n302), .B2(new_n230), .C1(new_n304), .C2(new_n202), .ZN(new_n305));
  NAND3_X1  g0105(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G1), .A2(G13), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT11), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT71), .ZN(new_n311));
  INV_X1    g0111(.A(G13), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(G1), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n311), .B1(new_n313), .B2(G20), .ZN(new_n314));
  NOR4_X1   g0114(.A1(new_n312), .A2(new_n213), .A3(KEYINPUT71), .A4(G1), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(new_n308), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n212), .A2(G20), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(G68), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n313), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n321), .A2(KEYINPUT12), .A3(new_n301), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n316), .A2(new_n225), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(KEYINPUT12), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n300), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n282), .A2(G200), .A3(new_n289), .ZN(new_n329));
  OAI21_X1  g0129(.A(G190), .B1(new_n297), .B2(new_n298), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n325), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT72), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n317), .A2(G77), .A3(new_n318), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n316), .A2(new_n230), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT15), .B(G87), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n302), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n339), .A2(new_n340), .B1(G20), .B2(G77), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT8), .B(G58), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT69), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n341), .B1(new_n343), .B2(new_n304), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT70), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n344), .A2(new_n345), .A3(new_n308), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n344), .B2(new_n308), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n337), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n271), .A2(new_n266), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT68), .B1(new_n349), .B2(new_n242), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n265), .A2(G1698), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT68), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(G232), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n284), .A2(new_n226), .B1(new_n232), .B2(new_n271), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n259), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n277), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(G244), .B2(new_n279), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G179), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n357), .B2(new_n360), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n348), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n355), .B1(new_n353), .B2(new_n350), .ZN(new_n367));
  OAI211_X1 g0167(.A(G190), .B(new_n359), .C1(new_n367), .C2(new_n259), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n337), .C1(new_n346), .C2(new_n347), .ZN(new_n369));
  OAI21_X1  g0169(.A(G200), .B1(new_n357), .B2(new_n360), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n334), .B1(new_n366), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n351), .A2(G222), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G223), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n284), .A2(new_n376), .B1(new_n230), .B2(new_n271), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n286), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n358), .B1(G226), .B2(new_n279), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(G169), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n362), .ZN(new_n382));
  INV_X1    g0182(.A(new_n308), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n248), .A2(KEYINPUT8), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT8), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G58), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(new_n340), .B1(G150), .B2(new_n303), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n203), .A2(G20), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n383), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(KEYINPUT67), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(KEYINPUT67), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n312), .A2(new_n213), .A3(G1), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n308), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n202), .B1(new_n212), .B2(G20), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n395), .A2(new_n396), .B1(new_n202), .B2(new_n394), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n381), .A2(new_n382), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n373), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n335), .A2(new_n336), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n344), .A2(new_n308), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT70), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n344), .A2(new_n345), .A3(new_n308), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(new_n370), .A3(new_n368), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n348), .A2(new_n363), .A3(new_n365), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n407), .A3(KEYINPUT72), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT10), .ZN(new_n409));
  INV_X1    g0209(.A(G200), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n378), .B2(new_n379), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(G190), .B2(new_n380), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n393), .A2(new_n397), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT9), .B1(new_n413), .B2(new_n391), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT9), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n392), .A2(new_n415), .A3(new_n393), .A4(new_n397), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n409), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n412), .A2(new_n417), .A3(new_n409), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n408), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT73), .B1(new_n400), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n399), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n406), .A2(new_n407), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n334), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n412), .A2(new_n417), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT10), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n412), .A2(new_n417), .A3(new_n409), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT73), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n424), .A2(new_n428), .A3(new_n429), .A4(new_n408), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT16), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n269), .A2(new_n213), .A3(new_n270), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT7), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n213), .A4(new_n270), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n225), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n248), .A2(new_n225), .ZN(new_n437));
  OAI21_X1  g0237(.A(G20), .B1(new_n437), .B2(new_n201), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n303), .A2(G159), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n431), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT7), .B1(new_n265), .B2(new_n213), .ZN(new_n442));
  NOR4_X1   g0242(.A1(new_n263), .A2(new_n264), .A3(new_n433), .A4(G20), .ZN(new_n443));
  OAI21_X1  g0243(.A(G68), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n440), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(KEYINPUT16), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n441), .A2(new_n446), .A3(new_n308), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n387), .A2(new_n318), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n448), .A2(new_n395), .B1(new_n394), .B2(new_n342), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n376), .A2(new_n266), .ZN(new_n451));
  INV_X1    g0251(.A(G226), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G1698), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n451), .B(new_n453), .C1(new_n263), .C2(new_n264), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G87), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n286), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT77), .ZN(new_n458));
  INV_X1    g0258(.A(G274), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n208), .B2(new_n258), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n279), .A2(G232), .B1(new_n460), .B2(new_n276), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n259), .B1(new_n454), .B2(new_n455), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n259), .A2(G232), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n277), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT77), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(G200), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n463), .A2(new_n466), .A3(G190), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n450), .A2(new_n470), .A3(KEYINPUT17), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n447), .B(new_n449), .C1(new_n468), .C2(new_n469), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT17), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n447), .A2(new_n449), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n463), .A2(new_n466), .A3(G179), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n462), .A2(new_n467), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(new_n364), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n476), .A2(KEYINPUT18), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT78), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n476), .A2(new_n479), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT18), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n481), .A3(new_n484), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n475), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND4_X1   g0288(.A1(new_n333), .A2(new_n421), .A3(new_n430), .A4(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT21), .ZN(new_n490));
  INV_X1    g0290(.A(new_n314), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n394), .A2(new_n311), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(new_n212), .B2(G33), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n383), .B(new_n495), .C1(new_n314), .C2(new_n315), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G283), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n498), .B(new_n213), .C1(G33), .C2(new_n261), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT84), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n493), .A2(G20), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n308), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(new_n308), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT20), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(KEYINPUT20), .B(new_n499), .C1(new_n502), .C2(new_n503), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n497), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n509));
  OAI211_X1 g0309(.A(G257), .B(new_n266), .C1(new_n263), .C2(new_n264), .ZN(new_n510));
  XOR2_X1   g0310(.A(KEYINPUT83), .B(G303), .Z(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(new_n510), .C1(new_n511), .C2(new_n271), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n512), .A2(new_n286), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n212), .A2(G45), .ZN(new_n514));
  OR2_X1    g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  NAND2_X1  g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n460), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n275), .A2(G1), .ZN(new_n519));
  INV_X1    g0319(.A(new_n516), .ZN(new_n520));
  NOR2_X1   g0320(.A1(KEYINPUT5), .A2(G41), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n259), .ZN(new_n523));
  INV_X1    g0323(.A(G270), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(G169), .B1(new_n513), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n490), .B1(new_n508), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n506), .A2(new_n507), .ZN(new_n528));
  INV_X1    g0328(.A(new_n497), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n517), .A2(new_n286), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(G270), .B1(new_n460), .B2(new_n517), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n512), .A2(new_n286), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n364), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(KEYINPUT21), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G200), .ZN(new_n537));
  INV_X1    g0337(.A(G190), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n508), .C1(new_n538), .C2(new_n536), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n513), .A2(new_n362), .A3(new_n525), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n530), .A2(new_n540), .ZN(new_n541));
  AND4_X1   g0341(.A1(new_n527), .A2(new_n535), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n259), .A2(G274), .A3(new_n519), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT80), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n460), .A2(KEYINPUT80), .A3(new_n519), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n259), .A2(G250), .A3(new_n514), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n260), .A2(new_n493), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G238), .A2(G1698), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n231), .B2(G1698), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n550), .B1(new_n552), .B2(new_n271), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n549), .B1(new_n553), .B2(new_n259), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n364), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n549), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n231), .A2(G1698), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(G238), .B2(G1698), .ZN(new_n558));
  OAI22_X1  g0358(.A1(new_n558), .A2(new_n265), .B1(new_n260), .B2(new_n493), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n556), .B1(new_n559), .B2(new_n286), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(new_n362), .A3(new_n547), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  AOI211_X1 g0362(.A(new_n308), .B(new_n394), .C1(new_n212), .C2(G33), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n339), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n213), .B(G68), .C1(new_n263), .C2(new_n264), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n302), .B2(new_n261), .ZN(new_n567));
  NAND3_X1  g0367(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G97), .A2(G107), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n213), .A2(new_n568), .B1(new_n569), .B2(new_n227), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT81), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n565), .B(new_n567), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n213), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n569), .A2(new_n227), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(KEYINPUT81), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n308), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n316), .A2(new_n338), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n564), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT82), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n575), .A2(KEYINPUT81), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n570), .A2(new_n571), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n565), .A4(new_n567), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(new_n308), .B1(new_n316), .B2(new_n338), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT82), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n564), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n562), .B1(new_n580), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n563), .A2(G87), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(new_n577), .A3(new_n578), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n560), .A2(G190), .A3(new_n547), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n410), .B1(new_n560), .B2(new_n547), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n594));
  OAI211_X1 g0394(.A(G250), .B(new_n266), .C1(new_n263), .C2(new_n264), .ZN(new_n595));
  INV_X1    g0395(.A(G294), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n594), .B(new_n595), .C1(new_n260), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n286), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT88), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n597), .A2(KEYINPUT88), .A3(new_n286), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n522), .A2(G264), .A3(new_n259), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n518), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n600), .A2(new_n538), .A3(new_n601), .A4(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n598), .A2(new_n518), .A3(new_n602), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n410), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT23), .B1(new_n213), .B2(G107), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT86), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(KEYINPUT86), .B(KEYINPUT23), .C1(new_n213), .C2(G107), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n611), .A2(new_n612), .B1(new_n213), .B2(new_n550), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n213), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT22), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(KEYINPUT85), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT23), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n232), .A3(G20), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT87), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT87), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n620), .A2(new_n617), .A3(new_n232), .A4(G20), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g0422(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n271), .A2(new_n623), .A3(new_n213), .A4(G87), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n613), .A2(new_n616), .A3(new_n622), .A4(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n625), .A2(KEYINPUT24), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(KEYINPUT24), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n308), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n563), .A2(G107), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n394), .A2(new_n232), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n630), .B(KEYINPUT25), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n608), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n616), .A2(new_n624), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT24), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(new_n622), .A4(new_n613), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n625), .A2(KEYINPUT24), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n383), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n629), .A2(new_n631), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n603), .B1(new_n598), .B2(new_n599), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n364), .B1(new_n640), .B2(new_n601), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n606), .A2(new_n362), .ZN(new_n642));
  OAI22_X1  g0442(.A1(new_n638), .A2(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(G244), .B(new_n266), .C1(new_n263), .C2(new_n264), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT79), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT4), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n271), .A2(G244), .A3(new_n266), .A4(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n647), .A2(new_n498), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n286), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n518), .B1(new_n523), .B2(new_n218), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n362), .A3(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n232), .A2(KEYINPUT6), .A3(G97), .ZN(new_n656));
  XNOR2_X1  g0456(.A(G97), .B(G107), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT6), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n659), .A2(new_n213), .B1(new_n230), .B2(new_n304), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n232), .B1(new_n434), .B2(new_n435), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n308), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n394), .A2(new_n261), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n563), .B2(G97), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n653), .B1(new_n651), .B2(new_n286), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n655), .B(new_n665), .C1(G169), .C2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n665), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n666), .A2(G200), .ZN(new_n669));
  AOI211_X1 g0469(.A(G190), .B(new_n653), .C1(new_n286), .C2(new_n651), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND4_X1   g0471(.A1(new_n633), .A2(new_n643), .A3(new_n667), .A4(new_n671), .ZN(new_n672));
  AND4_X1   g0472(.A1(new_n489), .A2(new_n542), .A3(new_n593), .A4(new_n672), .ZN(G372));
  NAND2_X1  g0473(.A1(new_n485), .A2(new_n480), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n328), .B1(new_n331), .B2(new_n366), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n475), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT91), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n428), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n426), .A2(KEYINPUT91), .A3(new_n427), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n422), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n489), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT26), .ZN(new_n683));
  NOR4_X1   g0483(.A1(new_n587), .A2(new_n667), .A3(new_n592), .A4(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT90), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n667), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n562), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n579), .A2(KEYINPUT82), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n585), .B1(new_n584), .B2(new_n564), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n590), .A2(new_n591), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT89), .B1(new_n584), .B2(new_n588), .ZN(new_n692));
  AND4_X1   g0492(.A1(KEYINPUT89), .A2(new_n588), .A3(new_n577), .A4(new_n578), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n362), .A2(new_n666), .B1(new_n662), .B2(new_n664), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n652), .A2(new_n654), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n364), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(KEYINPUT90), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n686), .A2(new_n690), .A3(new_n694), .A4(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n684), .B1(new_n683), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n652), .A2(new_n538), .A3(new_n654), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(G200), .B2(new_n666), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n702), .A2(new_n668), .B1(new_n695), .B2(new_n697), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n703), .A2(new_n690), .A3(new_n633), .A4(new_n694), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n600), .A2(new_n601), .A3(new_n604), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G169), .ZN(new_n706));
  INV_X1    g0506(.A(new_n606), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G179), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n628), .A2(new_n632), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n535), .A2(new_n527), .A3(new_n541), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n690), .B1(new_n704), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n700), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n681), .B1(new_n682), .B2(new_n713), .ZN(G369));
  OR3_X1    g0514(.A1(new_n321), .A2(KEYINPUT27), .A3(G20), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT27), .B1(new_n321), .B2(G20), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G213), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G343), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n530), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n542), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n710), .A2(new_n530), .A3(new_n719), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT92), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT92), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n721), .A2(new_n725), .A3(new_n722), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n719), .B1(new_n638), .B2(new_n639), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n709), .B1(new_n633), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n643), .A2(new_n719), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n724), .A2(G330), .A3(new_n726), .A4(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n729), .ZN(new_n733));
  INV_X1    g0533(.A(new_n719), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n710), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n733), .B1(new_n728), .B2(new_n735), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n732), .A2(new_n736), .ZN(G399));
  NOR2_X1   g0537(.A1(new_n217), .A2(G41), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n574), .A2(G116), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n739), .A2(G1), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n207), .B2(new_n739), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n734), .B1(new_n700), .B2(new_n712), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT94), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT94), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n747), .B(new_n734), .C1(new_n700), .C2(new_n712), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT95), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n704), .B2(new_n711), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n633), .A2(new_n667), .A3(new_n671), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n690), .A2(new_n694), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n643), .A2(new_n527), .A3(new_n541), .A4(new_n535), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n753), .A2(new_n755), .A3(new_n756), .A4(KEYINPUT95), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n699), .A2(KEYINPUT26), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n587), .A2(new_n592), .A3(new_n667), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n587), .B1(new_n759), .B2(new_n683), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n751), .A2(new_n757), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(KEYINPUT29), .A3(new_n734), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n672), .A2(new_n542), .A3(new_n593), .A4(new_n734), .ZN(new_n763));
  AND4_X1   g0563(.A1(new_n547), .A2(new_n560), .A3(new_n598), .A4(new_n602), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(new_n540), .A3(new_n666), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT30), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n764), .A2(new_n540), .A3(KEYINPUT30), .A4(new_n666), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n560), .A2(new_n547), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n536), .A2(new_n770), .A3(new_n362), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT93), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n707), .B2(new_n666), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n696), .A2(KEYINPUT93), .A3(new_n606), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n719), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT31), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g0578(.A(KEYINPUT31), .B(new_n719), .C1(new_n769), .C2(new_n775), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n763), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n749), .A2(new_n762), .B1(G330), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n743), .B1(new_n781), .B2(G1), .ZN(G364));
  AND2_X1   g0582(.A1(new_n724), .A2(new_n726), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(G330), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n312), .A2(G20), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n212), .B1(new_n785), .B2(G45), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n738), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n724), .A2(G330), .A3(new_n726), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(KEYINPUT96), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT96), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n724), .A2(new_n792), .A3(G330), .A4(new_n726), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n784), .A2(new_n789), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n307), .B1(G20), .B2(new_n364), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n362), .A2(G200), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT97), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n213), .B1(new_n796), .B2(KEYINPUT97), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n538), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G107), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n799), .A2(G190), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n271), .B1(new_n803), .B2(new_n227), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT98), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n805), .B2(new_n804), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT99), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n213), .A2(new_n362), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G190), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n410), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n213), .A2(G190), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n813), .A2(G179), .A3(new_n410), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n812), .A2(new_n202), .B1(new_n230), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n810), .A2(G200), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n809), .A2(new_n538), .A3(G200), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G58), .A2(new_n816), .B1(new_n818), .B2(G68), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n813), .A2(new_n362), .A3(new_n410), .ZN(new_n820));
  INV_X1    g0620(.A(G159), .ZN(new_n821));
  OAI21_X1  g0621(.A(KEYINPUT32), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OR3_X1    g0622(.A1(new_n820), .A2(KEYINPUT32), .A3(new_n821), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n819), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n538), .A2(G179), .A3(G200), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n213), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n815), .B(new_n824), .C1(G97), .C2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n808), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT100), .ZN(new_n830));
  INV_X1    g0630(.A(G317), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(KEYINPUT33), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n831), .A2(KEYINPUT33), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n818), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n816), .ZN(new_n835));
  INV_X1    g0635(.A(G322), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT101), .ZN(new_n838));
  INV_X1    g0638(.A(new_n814), .ZN(new_n839));
  INV_X1    g0639(.A(new_n820), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n839), .A2(G311), .B1(new_n840), .B2(G329), .ZN(new_n841));
  INV_X1    g0641(.A(G326), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n842), .B2(new_n812), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n271), .B(new_n843), .C1(G294), .C2(new_n827), .ZN(new_n844));
  INV_X1    g0644(.A(G283), .ZN(new_n845));
  INV_X1    g0645(.A(G303), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n844), .B1(new_n845), .B2(new_n800), .C1(new_n846), .C2(new_n803), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n829), .A2(new_n830), .B1(new_n838), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n829), .A2(new_n830), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n795), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n217), .A2(new_n271), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n207), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n852), .B1(new_n275), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n275), .B2(new_n251), .ZN(new_n855));
  INV_X1    g0655(.A(G355), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n216), .A2(new_n271), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n855), .B1(G116), .B2(new_n216), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(G13), .A2(G33), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(G20), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(new_n795), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n789), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n850), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT102), .ZN(new_n865));
  INV_X1    g0665(.A(new_n861), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n783), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n794), .B1(new_n865), .B2(new_n867), .ZN(G396));
  OAI22_X1  g0668(.A1(new_n369), .A2(new_n371), .B1(new_n405), .B2(new_n734), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n407), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n366), .A2(new_n734), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n745), .A2(new_n748), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n872), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n874), .B(new_n734), .C1(new_n700), .C2(new_n712), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n780), .A2(G330), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n788), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n877), .B2(new_n876), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n795), .A2(new_n859), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n789), .B1(new_n230), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n795), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n801), .A2(G87), .ZN(new_n883));
  INV_X1    g0683(.A(G311), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n883), .B1(new_n884), .B2(new_n820), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT104), .ZN(new_n886));
  XNOR2_X1  g0686(.A(KEYINPUT103), .B(G283), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n265), .B1(new_n817), .B2(new_n887), .C1(new_n261), .C2(new_n826), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n811), .A2(G303), .B1(new_n839), .B2(G116), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n596), .B2(new_n835), .ZN(new_n890));
  INV_X1    g0690(.A(new_n803), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n888), .B(new_n890), .C1(G107), .C2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n265), .B1(new_n840), .B2(G132), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n248), .B2(new_n826), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n800), .A2(new_n225), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n894), .B(new_n895), .C1(G50), .C2(new_n891), .ZN(new_n896));
  AOI22_X1  g0696(.A1(G143), .A2(new_n816), .B1(new_n818), .B2(G150), .ZN(new_n897));
  INV_X1    g0697(.A(G137), .ZN(new_n898));
  OAI221_X1 g0698(.A(new_n897), .B1(new_n898), .B2(new_n812), .C1(new_n821), .C2(new_n814), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT34), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n886), .A2(new_n892), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n881), .B1(new_n882), .B2(new_n901), .C1(new_n874), .C2(new_n860), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n879), .A2(new_n902), .ZN(G384));
  NOR2_X1   g0703(.A1(new_n209), .A2(new_n493), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n659), .B(KEYINPUT105), .Z(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT35), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n907), .B2(new_n906), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT36), .ZN(new_n910));
  OR3_X1    g0710(.A1(new_n207), .A2(new_n230), .A3(new_n437), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n202), .A2(G68), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n212), .B(G13), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n327), .A2(new_n719), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n717), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n476), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n483), .A2(new_n918), .A3(new_n472), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT37), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT37), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n483), .A2(new_n918), .A3(new_n921), .A4(new_n472), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n488), .B2(new_n918), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(KEYINPUT38), .B(new_n923), .C1(new_n488), .C2(new_n918), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(KEYINPUT106), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT106), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n924), .A2(new_n929), .A3(new_n925), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(KEYINPUT39), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n923), .ZN(new_n932));
  INV_X1    g0732(.A(new_n475), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n918), .B1(new_n933), .B2(new_n674), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n925), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n935), .A2(new_n927), .ZN(new_n936));
  XOR2_X1   g0736(.A(KEYINPUT107), .B(KEYINPUT39), .Z(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n916), .B1(new_n931), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n928), .A2(new_n930), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n875), .A2(new_n871), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n326), .A2(new_n719), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n327), .A2(new_n331), .A3(new_n942), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n326), .B(new_n719), .C1(new_n332), .C2(new_n300), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n940), .A2(new_n946), .B1(new_n674), .B2(new_n917), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n939), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n749), .A2(new_n489), .A3(new_n762), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n949), .A2(new_n681), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n948), .B(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(G330), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n779), .A2(KEYINPUT108), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n773), .A2(new_n774), .ZN(new_n954));
  INV_X1    g0754(.A(new_n771), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(new_n767), .A3(new_n768), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT108), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n957), .A2(new_n958), .A3(KEYINPUT31), .A4(new_n719), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n763), .A2(new_n953), .A3(new_n959), .A4(new_n778), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n872), .B1(new_n943), .B2(new_n944), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n928), .A2(new_n930), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT40), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n935), .B2(new_n927), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n963), .A2(new_n964), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n489), .A2(new_n960), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n952), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n966), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n951), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n212), .B2(new_n785), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n951), .A2(new_n969), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n914), .B1(new_n971), .B2(new_n972), .ZN(G367));
  NOR2_X1   g0773(.A1(new_n240), .A2(new_n852), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n862), .B1(new_n216), .B2(new_n338), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n826), .A2(new_n225), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n816), .A2(G150), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n898), .B2(new_n820), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n976), .B(new_n978), .C1(G143), .C2(new_n811), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n271), .B1(new_n817), .B2(new_n821), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(G50), .B2(new_n839), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n801), .A2(G77), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n891), .A2(G58), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n979), .A2(new_n981), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n800), .A2(new_n261), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n511), .A2(new_n835), .B1(new_n812), .B2(new_n884), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n265), .B1(new_n814), .B2(new_n887), .C1(new_n596), .C2(new_n817), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n826), .A2(new_n232), .B1(new_n820), .B2(new_n831), .ZN(new_n988));
  OR4_X1    g0788(.A1(new_n985), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n803), .A2(new_n493), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT46), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n984), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT47), .Z(new_n993));
  OAI221_X1 g0793(.A(new_n788), .B1(new_n974), .B2(new_n975), .C1(new_n993), .C2(new_n882), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT114), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n692), .A2(new_n693), .A3(new_n734), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT109), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n587), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n754), .B2(new_n997), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n995), .B1(new_n866), .B2(new_n999), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n671), .B(new_n667), .C1(new_n668), .C2(new_n734), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n695), .A2(new_n697), .A3(new_n719), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1003), .B(new_n733), .C1(new_n728), .C2(new_n735), .ZN(new_n1004));
  XOR2_X1   g0804(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1003), .ZN(new_n1007));
  AOI21_X1  g0807(.A(KEYINPUT44), .B1(new_n736), .B2(new_n1007), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n736), .A2(KEYINPUT44), .A3(new_n1007), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT113), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n731), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n735), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n730), .B(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n791), .A2(new_n1014), .A3(new_n793), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n790), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1010), .A2(KEYINPUT113), .A3(new_n732), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1012), .A2(new_n1017), .A3(new_n1018), .A4(new_n781), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n781), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n738), .B(KEYINPUT41), .Z(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n787), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT111), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(KEYINPUT111), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n730), .A2(new_n1013), .A3(new_n1003), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT42), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n667), .B1(new_n1001), .B2(new_n643), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1028), .A2(KEYINPUT42), .B1(new_n734), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT110), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n732), .A2(new_n1035), .A3(new_n1003), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1037));
  OAI21_X1  g0837(.A(KEYINPUT110), .B1(new_n731), .B2(new_n1007), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1037), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1034), .B(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1000), .B1(new_n1023), .B2(new_n1042), .ZN(G387));
  OAI21_X1  g0843(.A(new_n861), .B1(new_n728), .B2(new_n729), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n857), .A2(new_n740), .B1(G107), .B2(new_n216), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n343), .A2(G50), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT50), .ZN(new_n1047));
  AOI21_X1  g0847(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n740), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n852), .B1(new_n245), .B2(G45), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1045), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n862), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n788), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n803), .A2(new_n230), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n985), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n271), .B1(new_n817), .B2(new_n342), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G150), .B2(new_n840), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n826), .A2(new_n338), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G50), .B2(new_n816), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n811), .A2(G159), .B1(new_n839), .B2(G68), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1055), .A2(new_n1057), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G322), .A2(new_n811), .B1(new_n818), .B2(G311), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n831), .B2(new_n835), .C1(new_n511), .C2(new_n814), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n887), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n891), .A2(G294), .B1(new_n827), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT49), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n265), .B1(new_n842), .B2(new_n820), .C1(new_n800), .C2(new_n493), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1061), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1053), .B1(new_n1075), .B2(new_n795), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1017), .A2(new_n787), .B1(new_n1044), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1017), .A2(new_n781), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n738), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1017), .A2(new_n781), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(G393));
  NAND2_X1  g0881(.A1(new_n1019), .A2(new_n738), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1010), .B(new_n732), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n1078), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT115), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT115), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1083), .A2(new_n1078), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1082), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n862), .B1(new_n261), .B2(new_n216), .C1(new_n852), .C2(new_n254), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n788), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n826), .A2(new_n230), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n271), .B1(new_n817), .B2(new_n202), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(G143), .C2(new_n840), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n891), .A2(G68), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n343), .A2(new_n814), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1093), .A2(new_n883), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G150), .A2(new_n811), .B1(new_n816), .B2(G159), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT51), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n891), .A2(new_n1067), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n265), .B1(new_n817), .B2(new_n511), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G294), .B2(new_n839), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n827), .A2(G116), .B1(new_n840), .B2(G322), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n802), .A2(new_n1099), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G311), .A2(new_n816), .B1(new_n811), .B2(G317), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT52), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1096), .A2(new_n1098), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1090), .B1(new_n1106), .B2(new_n795), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n1003), .B2(new_n866), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1083), .B2(new_n786), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1088), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(G390));
  AND2_X1   g0911(.A1(new_n960), .A2(G330), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n780), .A2(G330), .A3(new_n874), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n945), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1112), .A2(new_n961), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n752), .A2(new_n754), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n587), .B1(new_n1116), .B2(new_n756), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n699), .A2(new_n683), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n759), .A2(KEYINPUT26), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n719), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1121), .A2(new_n870), .B1(new_n366), .B2(new_n734), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n960), .A2(G330), .A3(new_n874), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1123), .A2(new_n1114), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n780), .A2(G330), .A3(new_n945), .A4(new_n874), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n761), .A2(new_n734), .A3(new_n870), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n1126), .A3(new_n871), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1115), .A2(new_n1122), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n489), .A2(new_n1112), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n950), .A2(KEYINPUT116), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT116), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1123), .A2(new_n1114), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1125), .A2(new_n1126), .A3(new_n871), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n960), .A2(new_n961), .A3(G330), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1132), .A2(new_n1133), .B1(new_n1136), .B2(new_n941), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n949), .A2(new_n681), .A3(new_n1129), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1131), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n916), .B1(new_n1122), .B2(new_n1114), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(new_n931), .A3(new_n938), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n936), .A2(new_n915), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1126), .A2(new_n871), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1142), .B1(new_n1143), .B2(new_n1114), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1141), .A2(new_n1144), .A3(new_n1125), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1135), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1130), .B(new_n1139), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1135), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1141), .A2(new_n1144), .A3(new_n1125), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1147), .A2(new_n738), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT117), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT117), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1147), .A2(new_n1156), .A3(new_n738), .A4(new_n1153), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n931), .A2(new_n859), .A3(new_n938), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n880), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n788), .B1(new_n387), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n265), .B1(new_n803), .B2(new_n227), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT118), .Z(new_n1164));
  INV_X1    g0964(.A(new_n895), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1091), .B1(G107), .B2(new_n818), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n811), .A2(G283), .B1(new_n840), .B2(G294), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n816), .A2(G116), .B1(new_n839), .B2(G97), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n891), .A2(G150), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT53), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n816), .A2(G132), .ZN(new_n1172));
  INV_X1    g0972(.A(G128), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1172), .B1(new_n812), .B2(new_n1173), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n271), .B1(new_n817), .B2(new_n898), .C1(new_n821), .C2(new_n826), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT54), .B(G143), .ZN(new_n1176));
  INV_X1    g0976(.A(G125), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1176), .A2(new_n814), .B1(new_n820), .B2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1174), .A2(new_n1175), .A3(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n202), .B2(new_n800), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n1164), .A2(new_n1169), .B1(new_n1171), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1162), .B1(new_n1181), .B2(new_n795), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1159), .A2(new_n787), .B1(new_n1160), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1158), .A2(new_n1183), .ZN(G378));
  OR2_X1    g0984(.A1(new_n939), .A2(new_n947), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n398), .A2(new_n917), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n680), .B2(new_n399), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1186), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n422), .B(new_n1188), .C1(new_n678), .C2(new_n679), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1191), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n963), .A2(new_n964), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n952), .B1(new_n965), .B2(new_n962), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1185), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1204), .A2(new_n948), .A3(new_n1198), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1203), .A2(new_n859), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n788), .B1(G50), .B2(new_n1161), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n801), .A2(G58), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT119), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n820), .A2(new_n845), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n835), .A2(new_n232), .B1(new_n338), .B2(new_n814), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G116), .C2(new_n811), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n271), .A2(G41), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n976), .B(new_n1216), .C1(G97), .C2(new_n818), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1211), .A2(new_n1054), .A3(new_n1218), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1219), .A2(KEYINPUT58), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n835), .A2(new_n1173), .B1(new_n812), .B2(new_n1177), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G137), .B2(new_n839), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G150), .A2(new_n827), .B1(new_n818), .B2(G132), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n803), .C2(new_n1176), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n801), .A2(G159), .ZN(new_n1227));
  AOI211_X1 g1027(.A(G33), .B(G41), .C1(new_n840), .C2(G124), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1219), .A2(KEYINPUT58), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1216), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1220), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1208), .B1(new_n1232), .B2(new_n795), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1206), .A2(new_n787), .B1(new_n1207), .B2(new_n1233), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1204), .A2(new_n948), .A3(new_n1198), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n948), .B1(new_n1204), .B2(new_n1198), .ZN(new_n1236));
  OAI21_X1  g1036(.A(KEYINPUT57), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1138), .A2(KEYINPUT120), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT120), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n949), .A2(new_n1239), .A3(new_n681), .A4(new_n1129), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1159), .B2(new_n1151), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n738), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1241), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1153), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT57), .B1(new_n1245), .B2(new_n1206), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1234), .B1(new_n1243), .B2(new_n1246), .ZN(G375));
  NAND2_X1  g1047(.A1(new_n1128), .A2(new_n787), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT121), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n788), .B1(G68), .B2(new_n1161), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n835), .A2(new_n845), .B1(new_n812), .B2(new_n596), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n820), .A2(new_n846), .B1(new_n814), .B2(new_n232), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n271), .B(new_n1058), .C1(G116), .C2(new_n818), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n891), .A2(G97), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1254), .A2(new_n982), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n891), .A2(G159), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n271), .B1(new_n817), .B2(new_n1176), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G137), .B2(new_n816), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n839), .A2(G150), .B1(new_n840), .B2(G128), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G50), .A2(new_n827), .B1(new_n811), .B2(G132), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1258), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1257), .B1(new_n1211), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1251), .B1(new_n1264), .B2(new_n795), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n945), .B2(new_n860), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1250), .A2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT122), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1268), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT122), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1270), .A2(new_n1271), .A3(new_n1266), .A4(new_n1250), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1130), .A2(new_n1139), .A3(new_n1022), .A4(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(G381));
  OR2_X1    g1076(.A1(G393), .A2(G396), .ZN(new_n1277));
  OR4_X1    g1077(.A1(G384), .A2(G390), .A3(G387), .A4(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1154), .A2(new_n1183), .ZN(new_n1279));
  OR4_X1    g1079(.A1(G375), .A2(new_n1278), .A3(G381), .A4(new_n1279), .ZN(G407));
  OAI21_X1  g1080(.A(new_n787), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1207), .A2(new_n1233), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1245), .A2(new_n1206), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT57), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n739), .B1(new_n1287), .B2(new_n1245), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1283), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1279), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n718), .A2(G213), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1289), .A2(new_n1290), .A3(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(G407), .A2(G213), .A3(new_n1293), .ZN(G409));
  NAND3_X1  g1094(.A1(new_n1245), .A2(new_n1206), .A3(new_n1022), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1234), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1290), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1183), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(G375), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1137), .A2(KEYINPUT60), .A3(new_n1138), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT60), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT123), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n1274), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1302), .B2(new_n1274), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n738), .B(new_n1301), .C1(new_n1304), .C2(new_n1305), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1273), .A2(G384), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G384), .B1(new_n1273), .B2(new_n1306), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1300), .A2(new_n1291), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(KEYINPUT62), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT62), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1300), .A2(new_n1309), .A3(new_n1312), .A4(new_n1291), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1308), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1273), .A2(G384), .A3(new_n1306), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1292), .A2(G2897), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1314), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  OAI211_X1 g1117(.A(G2897), .B(new_n1292), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1279), .B1(new_n1234), .B2(new_n1295), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1319), .B1(G378), .B2(new_n1289), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1317), .B(new_n1318), .C1(new_n1320), .C2(new_n1292), .ZN(new_n1321));
  XOR2_X1   g1121(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1322));
  NAND4_X1  g1122(.A1(new_n1311), .A2(new_n1313), .A3(new_n1321), .A4(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT126), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1041), .B(new_n1033), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1021), .B1(new_n1019), .B2(new_n781), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1325), .B1(new_n1326), .B2(new_n787), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1327), .B(new_n1000), .C1(new_n1088), .C2(new_n1109), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G387), .A2(new_n1110), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(G393), .B(G396), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1328), .A2(new_n1329), .A3(KEYINPUT124), .A4(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT124), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1333), .B1(G387), .B2(new_n1110), .ZN(new_n1334));
  AOI22_X1  g1134(.A1(new_n1334), .A2(new_n1330), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1324), .B1(new_n1332), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1334), .A2(new_n1330), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1339), .A2(KEYINPUT126), .A3(new_n1331), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1336), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1323), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT63), .ZN(new_n1343));
  OR2_X1    g1143(.A1(new_n1310), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1310), .A2(new_n1343), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT61), .B1(new_n1339), .B2(new_n1331), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1344), .A2(new_n1321), .A3(new_n1345), .A4(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1342), .A2(new_n1347), .ZN(G405));
  OR3_X1    g1148(.A1(new_n1289), .A2(KEYINPUT127), .A3(new_n1279), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(G378), .A2(new_n1289), .ZN(new_n1350));
  OAI21_X1  g1150(.A(KEYINPUT127), .B1(new_n1289), .B2(new_n1279), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1349), .A2(new_n1350), .A3(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1309), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1336), .A2(new_n1340), .A3(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1353), .B1(new_n1336), .B2(new_n1340), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1352), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1341), .A2(new_n1309), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1352), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1336), .A2(new_n1340), .A3(new_n1353), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1357), .A2(new_n1358), .A3(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1356), .A2(new_n1360), .ZN(G402));
endmodule


