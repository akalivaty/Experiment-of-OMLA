//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n211), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(KEYINPUT9), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n246), .A2(new_n217), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n208), .A2(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G50), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G50), .ZN(new_n252));
  INV_X1    g0052(.A(new_n246), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT71), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n247), .A2(new_n217), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n209), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n257), .A2(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n209), .B1(new_n201), .B2(new_n252), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n256), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n254), .A2(new_n255), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n255), .B1(new_n254), .B2(new_n264), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n245), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n254), .A2(new_n264), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(new_n265), .A3(KEYINPUT9), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT65), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n274), .B1(new_n273), .B2(new_n275), .ZN(new_n277));
  OAI21_X1  g0077(.A(G226), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n273), .A2(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(new_n275), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1698), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G222), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n286), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(G223), .A3(G1698), .ZN(new_n290));
  AND2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G77), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n288), .A2(new_n290), .A3(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n217), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n282), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g0099(.A(KEYINPUT70), .B(G200), .Z(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n268), .A2(new_n271), .A3(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n298), .A2(G190), .A3(new_n281), .A4(new_n278), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT72), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n282), .A2(KEYINPUT72), .A3(G190), .A4(new_n298), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT10), .B1(new_n303), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n270), .A2(new_n265), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n311), .A2(new_n245), .B1(new_n299), .B2(new_n301), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(new_n308), .A4(new_n271), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G1698), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n293), .A2(new_n316), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n317), .A2(G238), .B1(G107), .B2(new_n293), .ZN(new_n318));
  NOR4_X1   g0118(.A1(new_n293), .A2(KEYINPUT67), .A3(new_n230), .A4(G1698), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT67), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n287), .B2(G232), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n318), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n297), .ZN(new_n323));
  OAI21_X1  g0123(.A(G244), .B1(new_n276), .B2(new_n277), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(KEYINPUT66), .A3(new_n281), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n281), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT66), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n323), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n301), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n249), .A2(G77), .ZN(new_n331));
  OAI22_X1  g0131(.A1(new_n248), .A2(new_n331), .B1(G77), .B2(new_n246), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT69), .ZN(new_n333));
  INV_X1    g0133(.A(G77), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n257), .A2(new_n261), .B1(new_n209), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT15), .B(G87), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT68), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n336), .A2(KEYINPUT68), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n258), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n335), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n256), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n333), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n339), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(new_n341), .A3(new_n337), .ZN(new_n346));
  INV_X1    g0146(.A(new_n335), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(KEYINPUT69), .A3(new_n256), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n332), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n323), .A2(G190), .A3(new_n325), .A4(new_n328), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n330), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G169), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n329), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n332), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT69), .B1(new_n348), .B2(new_n256), .ZN(new_n356));
  AOI211_X1 g0156(.A(new_n333), .B(new_n343), .C1(new_n346), .C2(new_n347), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G179), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n323), .A2(new_n359), .A3(new_n325), .A4(new_n328), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n352), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n299), .A2(new_n353), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n282), .A2(new_n359), .A3(new_n298), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n269), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n315), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n316), .A2(G226), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n289), .B(new_n367), .C1(G223), .C2(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G87), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n297), .ZN(new_n371));
  NOR2_X1   g0171(.A1(G41), .A2(G45), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n296), .A2(new_n217), .B1(new_n372), .B2(G1), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n280), .B1(G232), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G169), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n359), .B2(new_n376), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n257), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n249), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(KEYINPUT77), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n248), .B1(new_n381), .B2(KEYINPUT77), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n382), .A2(new_n383), .B1(new_n253), .B2(new_n257), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AND2_X1   g0185(.A1(G58), .A2(G68), .ZN(new_n386));
  OAI21_X1  g0186(.A(G20), .B1(new_n386), .B2(new_n201), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n260), .A2(G159), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n286), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT76), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n293), .A2(KEYINPUT76), .A3(KEYINPUT7), .A4(new_n209), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n285), .A2(new_n209), .A3(new_n286), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n392), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n389), .B1(new_n397), .B2(G68), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n343), .B1(new_n398), .B2(KEYINPUT16), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT16), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n396), .A2(new_n390), .ZN(new_n401));
  INV_X1    g0201(.A(G68), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n400), .B1(new_n403), .B2(new_n389), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n385), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT18), .B1(new_n379), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n399), .A2(new_n404), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n384), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n378), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n371), .A2(new_n375), .A3(G190), .ZN(new_n411));
  INV_X1    g0211(.A(G200), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n371), .B2(new_n375), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n407), .A2(new_n414), .A3(new_n384), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n405), .A2(KEYINPUT17), .A3(new_n414), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n406), .A2(new_n410), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n366), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n253), .A2(new_n402), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT12), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n402), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n334), .B2(new_n258), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(KEYINPUT11), .A3(new_n256), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n249), .A2(G68), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n422), .B(new_n425), .C1(new_n248), .C2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT11), .B1(new_n424), .B2(new_n256), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT14), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT73), .B1(new_n276), .B2(new_n277), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n373), .A2(KEYINPUT65), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT73), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(new_n436), .A3(G238), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT13), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G97), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n230), .A2(G1698), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(G226), .B2(G1698), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n441), .B2(new_n293), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n280), .B1(new_n442), .B2(new_n297), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n437), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n438), .B1(new_n437), .B2(new_n443), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n431), .B(G169), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT74), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n437), .A2(new_n443), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT13), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n437), .A2(new_n438), .A3(new_n443), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT74), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(new_n431), .A4(G169), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT75), .ZN(new_n455));
  OAI21_X1  g0255(.A(G169), .B1(new_n444), .B2(new_n445), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n444), .A2(new_n445), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n456), .A2(KEYINPUT14), .B1(new_n457), .B2(G179), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n454), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n455), .B1(new_n454), .B2(new_n458), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n430), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(G190), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n451), .A2(G200), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(new_n429), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n420), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT19), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n209), .B1(new_n439), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(G87), .B2(new_n206), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n209), .B(G68), .C1(new_n291), .C2(new_n292), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n466), .B1(new_n258), .B2(new_n204), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n256), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n253), .B1(new_n338), .B2(new_n339), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n208), .A2(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n246), .A2(new_n474), .A3(new_n217), .A4(new_n247), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G87), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n472), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(G1), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n279), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT80), .ZN(new_n483));
  INV_X1    g0283(.A(G250), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n208), .B2(G45), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(new_n273), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n273), .A3(new_n483), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n482), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(G244), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G116), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n287), .A2(KEYINPUT81), .A3(G238), .ZN(new_n493));
  OAI211_X1 g0293(.A(G238), .B(new_n316), .C1(new_n291), .C2(new_n292), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT81), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n492), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n489), .B(G190), .C1(new_n497), .C2(new_n273), .ZN(new_n498));
  INV_X1    g0298(.A(new_n488), .ZN(new_n499));
  OAI22_X1  g0299(.A1(new_n499), .A2(new_n486), .B1(new_n279), .B2(new_n481), .ZN(new_n500));
  INV_X1    g0300(.A(new_n492), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT81), .B1(new_n287), .B2(G238), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n494), .A2(new_n495), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n500), .B1(new_n504), .B2(new_n297), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n478), .B(new_n498), .C1(new_n505), .C2(new_n300), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n345), .A2(new_n337), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n472), .B(new_n473), .C1(new_n507), .C2(new_n475), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n489), .B(new_n359), .C1(new_n497), .C2(new_n273), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n508), .B(new_n509), .C1(new_n505), .C2(G169), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT79), .ZN(new_n512));
  OAI211_X1 g0312(.A(G244), .B(new_n316), .C1(new_n291), .C2(new_n292), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT4), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n289), .A2(KEYINPUT4), .A3(G244), .A4(new_n316), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G283), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n289), .A2(G250), .A3(G1698), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n515), .A2(new_n516), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n297), .ZN(new_n520));
  AND2_X1   g0320(.A1(KEYINPUT5), .A2(G41), .ZN(new_n521));
  NOR2_X1   g0321(.A1(KEYINPUT5), .A2(G41), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n480), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(G257), .A3(new_n273), .ZN(new_n524));
  XNOR2_X1  g0324(.A(KEYINPUT5), .B(G41), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n525), .A2(G274), .A3(new_n273), .A4(new_n480), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT78), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT78), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n524), .A2(new_n529), .A3(new_n526), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n520), .A2(new_n359), .A3(new_n528), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n260), .A2(G77), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n205), .A2(KEYINPUT6), .A3(G97), .ZN(new_n533));
  XNOR2_X1  g0333(.A(G97), .B(G107), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT6), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n532), .B1(new_n536), .B2(new_n209), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n205), .B1(new_n396), .B2(new_n390), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n256), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n246), .A2(G97), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n476), .B2(G97), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n531), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n527), .B1(new_n519), .B2(new_n297), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(G169), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n512), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n544), .A2(G169), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n547), .A2(KEYINPUT79), .A3(new_n531), .A4(new_n542), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n520), .A2(new_n528), .A3(new_n530), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n544), .A2(G190), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n550), .A2(new_n539), .A3(new_n541), .A4(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n511), .A2(new_n546), .A3(new_n548), .A4(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(G257), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n554));
  OAI211_X1 g0354(.A(G250), .B(new_n316), .C1(new_n291), .C2(new_n292), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G294), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n297), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n297), .B1(new_n480), .B2(new_n525), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G264), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n560), .A3(new_n526), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n353), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n558), .A2(new_n560), .A3(new_n359), .A4(new_n526), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n209), .B(G87), .C1(new_n291), .C2(new_n292), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT22), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT22), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n289), .A2(new_n567), .A3(new_n209), .A4(G87), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT24), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n491), .A2(G20), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT23), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n209), .B2(G107), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n569), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n570), .B1(new_n569), .B2(new_n575), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n256), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n253), .A2(KEYINPUT25), .A3(new_n205), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT25), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n246), .B2(G107), .ZN(new_n581));
  AOI22_X1  g0381(.A1(G107), .A2(new_n476), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n564), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n558), .A2(new_n560), .A3(G190), .A4(new_n526), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n561), .A2(G200), .ZN(new_n585));
  AND4_X1   g0385(.A1(new_n578), .A2(new_n582), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G116), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n247), .A2(new_n217), .B1(G20), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n517), .B(new_n209), .C1(G33), .C2(new_n204), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n589), .A2(KEYINPUT20), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT20), .B1(new_n589), .B2(new_n590), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n475), .A2(G116), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(G116), .B2(new_n253), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n353), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(G264), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT82), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT82), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n289), .A2(new_n599), .A3(G264), .A4(G1698), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n293), .A2(G303), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n289), .A2(G257), .A3(new_n316), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n598), .A2(new_n600), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n297), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n523), .A2(new_n273), .ZN(new_n605));
  INV_X1    g0405(.A(G270), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n526), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n596), .A2(new_n609), .A3(KEYINPUT21), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n607), .B1(new_n603), .B2(new_n297), .ZN(new_n611));
  INV_X1    g0411(.A(new_n594), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n253), .A2(G116), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n612), .A2(new_n613), .B1(new_n591), .B2(new_n592), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(G179), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n596), .A2(new_n609), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n616), .A2(KEYINPUT83), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT83), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n610), .A2(new_n620), .A3(new_n615), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n611), .A2(G190), .ZN(new_n622));
  INV_X1    g0422(.A(new_n614), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n622), .B(new_n623), .C1(new_n412), .C2(new_n611), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n587), .A2(new_n619), .A3(new_n621), .A4(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n465), .A2(new_n553), .A3(new_n625), .ZN(G372));
  INV_X1    g0426(.A(KEYINPUT84), .ZN(new_n627));
  INV_X1    g0427(.A(new_n315), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n417), .A2(new_n418), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n353), .B1(new_n449), .B2(new_n450), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n452), .B1(new_n631), .B2(new_n431), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n446), .A2(KEYINPUT74), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n458), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT75), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n454), .A2(new_n455), .A3(new_n458), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n429), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n464), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(new_n361), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n630), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n406), .A2(new_n410), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n628), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n365), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n627), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n639), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n461), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n641), .B1(new_n647), .B2(new_n630), .ZN(new_n648));
  OAI211_X1 g0448(.A(KEYINPUT84), .B(new_n365), .C1(new_n648), .C2(new_n628), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n465), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n546), .A2(new_n548), .A3(new_n552), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n578), .A2(new_n582), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(new_n562), .A3(new_n563), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n618), .A2(new_n617), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n654), .A2(new_n615), .A3(new_n610), .A4(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n578), .A2(new_n582), .A3(new_n584), .A4(new_n585), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n652), .A2(new_n656), .A3(new_n511), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n546), .A2(new_n548), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n511), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT26), .ZN(new_n661));
  INV_X1    g0461(.A(new_n510), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n506), .A2(new_n510), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n663), .A2(new_n545), .A3(new_n543), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n658), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n651), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n650), .A2(new_n668), .ZN(G369));
  NAND3_X1  g0469(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n623), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n655), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(new_n616), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n614), .A2(G169), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n680), .A2(new_n611), .A3(new_n617), .ZN(new_n681));
  AND4_X1   g0481(.A1(G179), .A2(new_n604), .A3(new_n614), .A4(new_n608), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT83), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n621), .A3(new_n655), .A4(new_n624), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n679), .B1(new_n684), .B2(new_n677), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n653), .A2(new_n675), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n587), .B1(new_n688), .B2(KEYINPUT85), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n688), .A2(KEYINPUT85), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n583), .A2(new_n675), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(KEYINPUT86), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(KEYINPUT86), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n689), .A2(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n654), .A2(new_n675), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n675), .B1(new_n619), .B2(new_n621), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n695), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(G41), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n212), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n208), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n703), .A2(new_n704), .B1(new_n216), .B2(new_n702), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT28), .Z(new_n706));
  AND2_X1   g0506(.A1(new_n611), .A2(G179), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n558), .A2(new_n560), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n505), .A3(new_n544), .A4(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n505), .A2(new_n708), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(KEYINPUT30), .A3(new_n707), .A4(new_n544), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n505), .A2(G179), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n549), .A3(new_n561), .A4(new_n609), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n711), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT31), .B1(new_n716), .B2(new_n675), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n546), .A2(new_n548), .A3(new_n552), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n720), .A2(new_n663), .A3(new_n675), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n654), .A2(new_n657), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n684), .A2(new_n722), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n721), .A2(new_n723), .A3(KEYINPUT87), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT87), .B1(new_n721), .B2(new_n723), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n719), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT29), .B1(new_n667), .B2(new_n676), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AND4_X1   g0530(.A1(new_n654), .A2(new_n683), .A3(new_n621), .A4(new_n655), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n731), .A2(new_n553), .A3(new_n586), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n543), .A2(new_n545), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n510), .A3(new_n506), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n662), .B1(new_n734), .B2(KEYINPUT26), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n659), .A2(new_n665), .A3(new_n511), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT29), .B(new_n676), .C1(new_n732), .C2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT88), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n652), .A2(new_n511), .A3(new_n657), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n736), .B(new_n735), .C1(new_n741), .C2(new_n731), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(KEYINPUT88), .A3(KEYINPUT29), .A4(new_n676), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n728), .B1(new_n730), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n706), .B1(new_n745), .B2(G1), .ZN(G364));
  AND2_X1   g0546(.A1(new_n209), .A2(G13), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G45), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT89), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n702), .A2(new_n749), .A3(new_n208), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n212), .A2(new_n289), .ZN(new_n751));
  INV_X1    g0551(.A(G355), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n751), .A2(new_n752), .B1(G116), .B2(new_n212), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n240), .A2(new_n479), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n212), .A2(new_n293), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n479), .B2(new_n216), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n217), .B1(G20), .B2(new_n353), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n750), .B1(new_n757), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n209), .A2(new_n359), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n412), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(KEYINPUT92), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(KEYINPUT92), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n766), .A2(G200), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT90), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n773), .A2(G50), .B1(G58), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n209), .A2(G179), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n301), .A2(G190), .A3(new_n778), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT93), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT93), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G87), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G179), .A2(G200), .ZN(new_n785));
  INV_X1    g0585(.A(G190), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n785), .A2(G20), .A3(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G159), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT32), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n209), .B1(new_n785), .B2(G190), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n204), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n765), .A2(new_n786), .A3(G200), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n289), .B1(new_n793), .B2(new_n402), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n790), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n301), .A2(new_n786), .A3(new_n778), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n205), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n765), .A2(new_n786), .A3(new_n412), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT91), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n798), .A2(new_n799), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n797), .B1(new_n804), .B2(G77), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n777), .A2(new_n784), .A3(new_n795), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n773), .A2(G326), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n783), .A2(G303), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n804), .A2(G311), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n289), .B1(new_n788), .B2(G329), .ZN(new_n810));
  INV_X1    g0610(.A(G294), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n791), .ZN(new_n812));
  INV_X1    g0612(.A(new_n796), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(G283), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT33), .B(G317), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(KEYINPUT94), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n793), .B1(new_n817), .B2(KEYINPUT94), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n818), .A2(new_n819), .B1(G322), .B2(new_n774), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT95), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n806), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n764), .B1(new_n822), .B2(new_n761), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT96), .ZN(new_n824));
  INV_X1    g0624(.A(new_n760), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n685), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n687), .A2(new_n750), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(G330), .B2(new_n685), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G396));
  NAND2_X1  g0630(.A1(new_n667), .A2(new_n676), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n352), .B1(new_n350), .B2(new_n676), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n361), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n361), .A2(new_n675), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n835), .A2(new_n667), .A3(new_n676), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n750), .B1(new_n839), .B2(new_n727), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n727), .B2(new_n839), .ZN(new_n841));
  INV_X1    g0641(.A(new_n793), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n804), .A2(G159), .B1(G150), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n776), .A2(G143), .ZN(new_n844));
  INV_X1    g0644(.A(G137), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n772), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT34), .Z(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n289), .B1(new_n787), .B2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT98), .Z(new_n850));
  INV_X1    g0650(.A(new_n791), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n813), .A2(G68), .B1(G58), .B2(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n850), .B(new_n852), .C1(new_n782), .C2(new_n252), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT97), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n793), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n793), .A2(new_n855), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n859), .A2(G283), .B1(G87), .B2(new_n813), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n588), .B2(new_n803), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n289), .B(new_n792), .C1(G311), .C2(new_n788), .ZN(new_n862));
  INV_X1    g0662(.A(new_n774), .ZN(new_n863));
  INV_X1    g0663(.A(G303), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n862), .B1(new_n811), .B2(new_n863), .C1(new_n772), .C2(new_n864), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n861), .B(new_n865), .C1(G107), .C2(new_n783), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n761), .B1(new_n854), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n750), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n761), .A2(new_n758), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n334), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n867), .B(new_n870), .C1(new_n835), .C2(new_n759), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n841), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(G384));
  INV_X1    g0673(.A(new_n536), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n874), .A2(KEYINPUT35), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(KEYINPUT35), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n875), .A2(G116), .A3(new_n218), .A4(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(KEYINPUT99), .B(KEYINPUT36), .Z(new_n878));
  XNOR2_X1  g0678(.A(new_n877), .B(new_n878), .ZN(new_n879));
  OR3_X1    g0679(.A1(new_n215), .A2(new_n334), .A3(new_n386), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n252), .A2(G68), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n208), .B(G13), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n465), .A2(new_n729), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n744), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT101), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n744), .A2(new_n884), .A3(KEYINPUT101), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n650), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n635), .A2(new_n636), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n430), .B(new_n675), .C1(new_n891), .C2(new_n638), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n429), .A2(new_n676), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n461), .A2(new_n464), .A3(new_n894), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n892), .A2(new_n895), .B1(new_n838), .B2(new_n834), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n398), .A2(KEYINPUT16), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n385), .B1(new_n897), .B2(new_n399), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n415), .B1(new_n673), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n379), .A2(new_n898), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT37), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n408), .A2(new_n378), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n673), .B(KEYINPUT100), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n408), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n902), .A2(new_n904), .A3(new_n905), .A4(new_n415), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n898), .A2(new_n673), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n419), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n907), .A2(new_n909), .A3(KEYINPUT38), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n896), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n907), .A2(new_n909), .A3(KEYINPUT38), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n415), .B1(new_n379), .B2(new_n405), .ZN(new_n918));
  INV_X1    g0718(.A(new_n903), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n405), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT37), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n906), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n419), .A2(new_n920), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n916), .B1(new_n917), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n912), .A2(KEYINPUT39), .A3(new_n913), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n461), .A2(new_n675), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n641), .A2(new_n919), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n915), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n890), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n892), .A2(new_n895), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT87), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n652), .A2(new_n511), .A3(new_n676), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n934), .B1(new_n935), .B2(new_n625), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n721), .A2(new_n723), .A3(KEYINPUT87), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n836), .B1(new_n938), .B2(new_n719), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n933), .A2(new_n914), .A3(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n922), .A2(new_n923), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n911), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n941), .B1(new_n944), .B2(new_n913), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n933), .A3(new_n939), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n651), .A2(new_n726), .ZN(new_n948));
  OAI21_X1  g0748(.A(G330), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n947), .B2(new_n948), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n932), .A2(new_n950), .B1(new_n208), .B2(new_n747), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n932), .A2(new_n950), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n883), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT102), .ZN(G367));
  OAI221_X1 g0754(.A(new_n762), .B1(new_n507), .B2(new_n212), .C1(new_n236), .C2(new_n755), .ZN(new_n955));
  INV_X1    g0755(.A(new_n859), .ZN(new_n956));
  INV_X1    g0756(.A(G159), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n956), .A2(new_n957), .B1(new_n252), .B2(new_n803), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n796), .A2(new_n334), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n289), .B1(new_n787), .B2(new_n845), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n773), .A2(G143), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n791), .A2(new_n402), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n774), .B2(G150), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT109), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n783), .A2(G58), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n961), .A2(new_n962), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(G283), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n956), .A2(new_n811), .B1(new_n968), .B2(new_n803), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n796), .A2(new_n204), .ZN(new_n970));
  INV_X1    g0770(.A(G317), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n293), .B1(new_n787), .B2(new_n971), .C1(new_n205), .C2(new_n791), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n783), .A2(KEYINPUT46), .A3(G116), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n773), .A2(G311), .B1(G303), .B2(new_n776), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT46), .B1(new_n783), .B2(G116), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n967), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  INV_X1    g0779(.A(new_n761), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n750), .B(new_n955), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT110), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT110), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n478), .A2(new_n676), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n662), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n663), .B2(new_n984), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n982), .B(new_n983), .C1(new_n825), .C2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n694), .A2(new_n697), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n733), .A2(new_n675), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT104), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n542), .A2(new_n675), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n652), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT103), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT103), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n652), .A2(new_n994), .A3(new_n991), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n990), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT42), .B1(new_n988), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n988), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n993), .A2(new_n995), .ZN(new_n999));
  INV_X1    g0799(.A(new_n990), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT42), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n998), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n659), .B1(new_n1001), .B2(new_n583), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n997), .B(new_n1003), .C1(new_n1004), .C2(new_n675), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(KEYINPUT105), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT105), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1005), .A2(new_n1010), .A3(new_n1006), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1009), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1012), .A2(new_n1013), .B1(new_n695), .B2(new_n996), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1009), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n695), .A2(new_n996), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n701), .B(KEYINPUT41), .ZN(new_n1022));
  OAI211_X1 g0822(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n698), .C2(new_n1001), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n696), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n988), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n1026));
  OR2_X1    g0826(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1025), .A2(new_n996), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n698), .A2(new_n1001), .A3(KEYINPUT45), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT45), .B1(new_n698), .B2(new_n1001), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1023), .B(new_n1028), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n695), .A2(KEYINPUT107), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT45), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n1025), .B2(new_n996), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n698), .A2(new_n1001), .A3(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1032), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n1023), .A4(new_n1028), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n694), .A2(new_n697), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n998), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n686), .A2(KEYINPUT108), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n686), .B(KEYINPUT108), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1033), .A2(new_n1039), .A3(new_n1045), .A4(new_n745), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1022), .B1(new_n1046), .B2(new_n745), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n749), .A2(new_n208), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n987), .B1(new_n1021), .B2(new_n1050), .ZN(G387));
  AOI21_X1  g0851(.A(new_n701), .B1(new_n1045), .B2(new_n745), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n745), .B2(new_n1045), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n694), .A2(new_n825), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n751), .A2(new_n704), .B1(G107), .B2(new_n212), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n755), .B1(new_n233), .B2(G45), .ZN(new_n1056));
  XOR2_X1   g0856(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1057));
  OR3_X1    g0857(.A1(new_n1057), .A2(G50), .A3(new_n257), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n704), .A2(KEYINPUT111), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n479), .B1(new_n402), .B2(new_n334), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n704), .B2(KEYINPUT111), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1057), .B1(G50), .B2(new_n257), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1055), .B1(new_n1056), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n750), .B1(new_n1064), .B2(new_n763), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT113), .Z(new_n1066));
  AOI21_X1  g0866(.A(new_n289), .B1(new_n788), .B2(G326), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n782), .A2(new_n811), .B1(new_n968), .B2(new_n791), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G303), .A2(new_n804), .B1(new_n859), .B2(G311), .ZN(new_n1069));
  INV_X1    g0869(.A(G322), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1069), .B1(new_n772), .B2(new_n1070), .C1(new_n971), .C2(new_n775), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1068), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT49), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1067), .B1(new_n588), .B2(new_n796), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n783), .A2(G77), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n293), .B(new_n970), .C1(G150), .C2(new_n788), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT114), .Z(new_n1081));
  NAND2_X1  g0881(.A1(new_n804), .A2(G68), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G50), .A2(new_n774), .B1(new_n842), .B2(new_n380), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n957), .B2(new_n772), .C1(new_n507), .C2(new_n791), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1076), .A2(new_n1077), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1054), .B(new_n1066), .C1(new_n1086), .C2(new_n761), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1053), .A2(new_n1088), .ZN(G393));
  INV_X1    g0889(.A(new_n695), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1031), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1037), .A2(new_n695), .A3(new_n1023), .A4(new_n1028), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n1092), .A3(new_n1049), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n762), .B1(new_n204), .B2(new_n212), .C1(new_n243), .C2(new_n755), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n750), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n773), .A2(G317), .B1(G311), .B2(new_n774), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT52), .Z(new_n1097));
  NAND2_X1  g0897(.A1(new_n804), .A2(G294), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n859), .A2(G303), .B1(G116), .B2(new_n851), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n289), .B(new_n797), .C1(G322), .C2(new_n788), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n968), .B2(new_n782), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT115), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n772), .A2(new_n259), .B1(new_n957), .B2(new_n863), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT51), .Z(new_n1105));
  AOI22_X1  g0905(.A1(new_n380), .A2(new_n804), .B1(new_n859), .B2(G50), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n293), .B1(new_n788), .B2(G143), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n334), .B2(new_n791), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G87), .B2(new_n813), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1106), .B(new_n1109), .C1(new_n402), .C2(new_n782), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1100), .A2(new_n1103), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1095), .B1(new_n1111), .B2(new_n761), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1001), .B2(new_n825), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1093), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT116), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT116), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1093), .A2(new_n1116), .A3(new_n1113), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1045), .A2(new_n745), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(new_n702), .A3(new_n1046), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(KEYINPUT117), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT117), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1121), .A2(new_n1124), .A3(new_n702), .A4(new_n1046), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1118), .A2(new_n1123), .A3(new_n1125), .ZN(G390));
  NAND2_X1  g0926(.A1(new_n925), .A2(new_n926), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n896), .B2(new_n927), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n933), .A2(G330), .A3(new_n939), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n742), .A2(new_n676), .A3(new_n833), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n834), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n933), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n927), .B1(new_n913), .B2(new_n944), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1128), .A2(new_n1129), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1129), .B1(new_n1128), .B2(new_n1134), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n728), .A2(new_n651), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n889), .A2(new_n650), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n726), .A2(G330), .A3(new_n835), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(new_n895), .A3(new_n892), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1131), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1141), .A2(new_n1129), .A3(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n838), .A2(new_n834), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n1141), .B2(new_n1129), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1137), .A2(new_n1139), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n889), .A2(new_n650), .A3(new_n1138), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n1148), .A2(new_n1149), .B1(new_n1136), .B2(new_n1135), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n702), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1127), .A2(new_n758), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n869), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n750), .B1(new_n380), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n863), .A2(new_n588), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n293), .B1(new_n787), .B2(new_n811), .C1(new_n334), .C2(new_n791), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(new_n773), .C2(G283), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n859), .A2(G107), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n804), .A2(G97), .B1(G68), .B2(new_n813), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1157), .A2(new_n784), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n863), .A2(new_n848), .ZN(new_n1161));
  INV_X1    g0961(.A(G125), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n289), .B1(new_n787), .B2(new_n1162), .C1(new_n957), .C2(new_n791), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1161), .B(new_n1163), .C1(new_n773), .C2(G128), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n956), .A2(new_n845), .B1(new_n252), .B2(new_n796), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT54), .B(G143), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1165), .B1(new_n804), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT53), .B1(new_n782), .B2(new_n259), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n782), .A2(KEYINPUT53), .A3(new_n259), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1160), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1154), .B1(new_n1172), .B2(new_n761), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1137), .A2(new_n1049), .B1(new_n1152), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1151), .A2(new_n1174), .ZN(G378));
  NAND2_X1  g0975(.A1(new_n315), .A2(new_n365), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n673), .B1(new_n270), .B2(new_n265), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OR3_X1    g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n940), .A2(new_n941), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n946), .A2(G330), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n942), .A2(G330), .A3(new_n946), .A4(new_n1184), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1188), .A2(new_n931), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n931), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1049), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n750), .B1(G50), .B2(new_n1153), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n289), .A2(G41), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G50), .B(new_n1194), .C1(new_n284), .C2(new_n700), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n773), .A2(G116), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1194), .B1(new_n968), .B2(new_n787), .C1(new_n204), .C2(new_n793), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n963), .B(new_n1197), .C1(G107), .C2(new_n774), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n804), .A2(new_n340), .B1(G58), .B2(new_n813), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1196), .A2(new_n1078), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT58), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1195), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G128), .A2(new_n774), .B1(new_n842), .B2(G132), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n259), .B2(new_n791), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G137), .B2(new_n804), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n1162), .B2(new_n772), .C1(new_n782), .C2(new_n1166), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n813), .A2(G159), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G33), .B(G41), .C1(new_n788), .C2(G124), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1202), .B1(new_n1201), .B2(new_n1200), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1193), .B1(new_n1212), .B2(new_n761), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1184), .B2(new_n759), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1192), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(KEYINPUT57), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1148), .B1(new_n1137), .B2(new_n1146), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n702), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n930), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1188), .A2(new_n931), .A3(new_n1189), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1136), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1128), .A2(new_n1134), .A3(new_n1129), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1139), .B1(new_n1225), .B2(new_n1149), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT57), .B1(new_n1222), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1215), .B1(new_n1218), .B2(new_n1227), .ZN(G375));
  INV_X1    g1028(.A(KEYINPUT118), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1149), .B2(new_n1048), .ZN(new_n1230));
  OAI211_X1 g1030(.A(KEYINPUT118), .B(new_n1049), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n933), .A2(new_n759), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT119), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n868), .B1(new_n402), .B2(new_n869), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n293), .B1(new_n788), .B2(G128), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n252), .B2(new_n791), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G58), .B2(new_n813), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1237), .B1(new_n259), .B2(new_n803), .C1(new_n782), .C2(new_n957), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n773), .A2(G132), .B1(new_n859), .B2(new_n1167), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n845), .B2(new_n775), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1238), .B1(new_n1240), .B2(KEYINPUT120), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(KEYINPUT120), .B2(new_n1240), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n293), .B1(new_n787), .B2(new_n864), .C1(new_n863), .C2(new_n968), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n959), .B(new_n1243), .C1(new_n773), .C2(G294), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n783), .A2(G97), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n859), .A2(G116), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n804), .A2(G107), .B1(new_n340), .B2(new_n851), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1242), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1233), .B(new_n1234), .C1(new_n980), .C2(new_n1249), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1230), .A2(new_n1231), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1139), .A2(new_n1146), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1022), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(G381));
  NOR2_X1   g1056(.A1(G393), .A2(G396), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n872), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(G387), .A2(new_n1258), .A3(G390), .A4(G381), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT121), .ZN(new_n1260));
  OR2_X1    g1060(.A1(G375), .A2(G378), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1260), .A2(new_n1261), .ZN(G407));
  OAI211_X1 g1062(.A(G407), .B(G213), .C1(G343), .C2(new_n1261), .ZN(G409));
  INV_X1    g1063(.A(KEYINPUT124), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1118), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(G387), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n829), .B1(new_n1053), .B2(new_n1088), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1257), .A2(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(G387), .A2(new_n1265), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1014), .B(new_n1020), .C1(new_n1047), .C2(new_n1049), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G390), .B1(new_n1270), .B2(new_n987), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n1266), .A2(new_n1268), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(G387), .A2(new_n1265), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1268), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G390), .A2(new_n1270), .A3(new_n987), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1273), .A2(new_n1274), .A3(new_n1264), .A4(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G375), .A2(G378), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n674), .A2(G213), .ZN(new_n1280));
  AND4_X1   g1080(.A1(new_n1151), .A2(new_n1174), .A3(new_n1192), .A4(new_n1214), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1222), .A2(new_n1253), .A3(new_n1226), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1280), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1148), .A2(new_n1149), .A3(KEYINPUT60), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n702), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT60), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1230), .A2(new_n1231), .A3(new_n1250), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n872), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT60), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1254), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(new_n702), .A3(new_n1252), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G384), .B(new_n1251), .C1(new_n1292), .C2(new_n1284), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1289), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1279), .A2(new_n1283), .A3(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1297));
  OR3_X1    g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1295), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT123), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1289), .A2(new_n1293), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1301), .B1(new_n1289), .B2(new_n1293), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1280), .A2(G2897), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1302), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1279), .A2(new_n1283), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1289), .A2(new_n1293), .A3(new_n1301), .A4(new_n1304), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1278), .B1(new_n1300), .B2(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1279), .A2(new_n1283), .A3(new_n1294), .A4(KEYINPUT63), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1309), .A2(new_n1310), .A3(new_n1277), .A4(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT122), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1316), .B1(new_n1295), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1295), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(KEYINPUT125), .B1(new_n1315), .B2(new_n1321), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1295), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1323), .A2(new_n1318), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT125), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1324), .A2(new_n1314), .A3(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1312), .B1(new_n1322), .B2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(KEYINPUT127), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1329), .B(new_n1312), .C1(new_n1322), .C2(new_n1326), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(G405));
  NAND2_X1  g1131(.A1(new_n1261), .A2(new_n1279), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1332), .B(new_n1294), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1333), .B(new_n1277), .ZN(G402));
endmodule


