//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(G250), .B1(G257), .B2(G264), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n210), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n217), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT64), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G68), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  INV_X1    g0029(.A(G87), .ZN(new_n230));
  INV_X1    g0030(.A(G250), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n233));
  INV_X1    g0033(.A(G58), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  INV_X1    g0035(.A(G257), .ZN(new_n236));
  OAI221_X1 g0036(.A(new_n233), .B1(new_n234), .B2(new_n235), .C1(new_n205), .C2(new_n236), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n212), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT1), .Z(new_n239));
  NAND2_X1  g0039(.A1(new_n226), .A2(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n235), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT2), .B(G226), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT66), .ZN(new_n247));
  XOR2_X1   g0047(.A(G264), .B(G270), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n245), .B(new_n249), .Z(G358));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n251), .B(new_n252), .Z(new_n253));
  XOR2_X1   g0053(.A(G107), .B(G116), .Z(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT7), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n258), .A2(new_n259), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(KEYINPUT7), .B1(new_n265), .B2(new_n210), .ZN(new_n266));
  OAI21_X1  g0066(.A(G68), .B1(new_n260), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n234), .A2(new_n228), .ZN(new_n268));
  OAI21_X1  g0068(.A(G20), .B1(new_n268), .B2(new_n201), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G159), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n267), .A2(KEYINPUT16), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT16), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n259), .B1(new_n258), .B2(G20), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n228), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n278), .B2(new_n272), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n221), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n274), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  XOR2_X1   g0082(.A(KEYINPUT8), .B(G58), .Z(new_n283));
  NAND2_X1  g0083(.A1(new_n209), .A2(G20), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(new_n221), .A3(new_n280), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n286), .ZN(new_n289));
  INV_X1    g0089(.A(new_n283), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n285), .A2(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n282), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(G226), .A2(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n262), .A2(new_n264), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT75), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G87), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n262), .A2(new_n264), .A3(G223), .A4(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n262), .A2(new_n264), .A3(new_n293), .A4(KEYINPUT75), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n296), .A2(new_n297), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G41), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(G1), .A3(G13), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT67), .ZN(new_n306));
  AND2_X1   g0106(.A1(G33), .A2(G41), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n221), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n302), .A2(KEYINPUT67), .A3(G1), .A4(G13), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G232), .ZN(new_n312));
  INV_X1    g0112(.A(G274), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n311), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n305), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n310), .A2(KEYINPUT76), .A3(new_n314), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT76), .B1(new_n310), .B2(new_n314), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n305), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n318), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n292), .A2(KEYINPUT17), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT17), .ZN(new_n327));
  INV_X1    g0127(.A(new_n324), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(new_n321), .B1(new_n317), .B2(new_n316), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n282), .A2(new_n291), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n327), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT79), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT18), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT76), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n311), .A2(new_n313), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(G232), .B2(new_n311), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n308), .A2(new_n309), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G179), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n310), .A2(KEYINPUT76), .A3(new_n314), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n305), .A2(new_n339), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT77), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT75), .B1(new_n258), .B2(new_n293), .ZN(new_n346));
  AND4_X1   g0146(.A1(KEYINPUT75), .A2(new_n262), .A3(new_n264), .A4(new_n293), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n299), .A2(new_n297), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n303), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n315), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n345), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(G179), .B1(new_n301), .B2(new_n304), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n353), .A2(KEYINPUT77), .A3(new_n339), .A4(new_n341), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n344), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT78), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n292), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n344), .A2(KEYINPUT78), .A3(new_n352), .A4(new_n354), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n334), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n354), .A2(new_n352), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT77), .B1(new_n321), .B2(new_n353), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n356), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n362), .A2(new_n334), .A3(new_n330), .A4(new_n358), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n333), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n330), .A3(new_n358), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT18), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n367), .A2(KEYINPUT79), .A3(new_n363), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n332), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n258), .A2(G222), .A3(new_n298), .ZN(new_n370));
  INV_X1    g0170(.A(G77), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n258), .A2(G1698), .ZN(new_n372));
  INV_X1    g0172(.A(G223), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n370), .B1(new_n371), .B2(new_n258), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n304), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n310), .A2(new_n336), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n377));
  XOR2_X1   g0177(.A(KEYINPUT68), .B(G226), .Z(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n375), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT72), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n381), .A2(G190), .B1(new_n382), .B2(KEYINPUT10), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(G200), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n382), .A2(KEYINPUT10), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT9), .ZN(new_n388));
  INV_X1    g0188(.A(new_n281), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT69), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n261), .B2(G20), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n210), .A2(KEYINPUT69), .A3(G33), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n283), .A2(new_n393), .B1(G150), .B2(new_n270), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT70), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n394), .A2(new_n395), .B1(G20), .B2(new_n203), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n389), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n284), .A2(G50), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n287), .A2(new_n399), .B1(G50), .B2(new_n286), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n388), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n398), .A2(new_n400), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT9), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n385), .A2(new_n387), .A3(new_n401), .A4(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n383), .A2(new_n403), .A3(new_n401), .A4(new_n384), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n386), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n380), .A2(new_n345), .ZN(new_n407));
  OAI221_X1 g0207(.A(new_n407), .B1(G179), .B2(new_n380), .C1(new_n398), .C2(new_n400), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n258), .A2(G232), .A3(G1698), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n258), .A2(G226), .A3(new_n298), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G97), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n413), .A2(new_n304), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n308), .A2(G238), .A3(new_n309), .A4(new_n311), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n376), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT13), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n304), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT13), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n418), .A2(new_n419), .A3(new_n376), .A4(new_n415), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(G190), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n284), .A2(G68), .ZN(new_n422));
  OR3_X1    g0222(.A1(new_n287), .A2(KEYINPUT73), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT73), .B1(new_n287), .B2(new_n422), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n371), .B1(new_n391), .B2(new_n392), .ZN(new_n426));
  INV_X1    g0226(.A(new_n270), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n427), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n281), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT11), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n425), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n430), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n289), .A2(new_n228), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT12), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n421), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n317), .B1(new_n417), .B2(new_n420), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT74), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n417), .A2(new_n420), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G200), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT74), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n436), .A4(new_n421), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n436), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT14), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n440), .A2(new_n446), .A3(G169), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n417), .A2(G179), .A3(new_n420), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n440), .B2(G169), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n372), .A2(new_n229), .B1(new_n206), .B2(new_n258), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n265), .A2(new_n235), .A3(G1698), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n304), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n377), .A2(G244), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n376), .A3(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n456), .A2(new_n345), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n284), .A2(G77), .ZN(new_n458));
  OAI22_X1  g0258(.A1(new_n287), .A2(new_n458), .B1(G77), .B2(new_n286), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT71), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n283), .A2(new_n270), .B1(G20), .B2(G77), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT15), .B(G87), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n393), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n460), .B1(new_n465), .B2(new_n389), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n461), .A2(new_n464), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(KEYINPUT71), .A3(new_n281), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n459), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n456), .A2(G179), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n457), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n456), .A2(G200), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n469), .B(new_n473), .C1(new_n323), .C2(new_n456), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n444), .A2(new_n451), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n409), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n369), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n262), .A2(new_n264), .A3(G244), .A4(new_n298), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT4), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n258), .A2(KEYINPUT4), .A3(G244), .A4(new_n298), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n304), .ZN(new_n486));
  INV_X1    g0286(.A(G45), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n487), .A2(new_n313), .A3(G1), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT5), .B(G41), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n308), .A2(new_n488), .A3(new_n489), .A4(new_n309), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n487), .A2(G1), .ZN(new_n491));
  AND2_X1   g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  NOR2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n494), .A2(new_n308), .A3(G257), .A4(new_n309), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n486), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n345), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n490), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n485), .B2(new_n304), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n340), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n501));
  OR2_X1    g0301(.A1(KEYINPUT80), .A2(G97), .ZN(new_n502));
  NAND2_X1  g0302(.A1(KEYINPUT80), .A2(G97), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G97), .A2(G107), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT6), .B1(new_n207), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(G20), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n371), .B2(new_n427), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n206), .B1(new_n276), .B2(new_n277), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n281), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n286), .A2(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n209), .A2(G33), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n286), .A2(new_n512), .A3(new_n221), .A4(new_n280), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n511), .B1(new_n514), .B2(G97), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n497), .A2(new_n500), .A3(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n499), .A2(G190), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT81), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n496), .A2(G200), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n499), .A2(new_n519), .A3(G190), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(new_n510), .A3(new_n515), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n517), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n262), .A2(new_n264), .A3(new_n210), .A4(G87), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT22), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT22), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n258), .A2(new_n527), .A3(new_n210), .A4(G87), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT84), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n530), .B(KEYINPUT23), .C1(new_n210), .C2(G107), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n206), .A2(G20), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n530), .B1(new_n533), .B2(KEYINPUT23), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT23), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(new_n206), .A3(G20), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n532), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT24), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n529), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n529), .B2(new_n539), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n281), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT25), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n286), .B2(G107), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n286), .A2(new_n544), .A3(G107), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n546), .A2(new_n547), .B1(new_n206), .B2(new_n513), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n494), .A2(new_n308), .A3(G264), .A4(new_n309), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G250), .A2(G1698), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n236), .B2(G1698), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(new_n258), .B1(G33), .B2(G294), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n490), .B(new_n550), .C1(new_n553), .C2(new_n303), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G190), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(G200), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n543), .A2(new_n549), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n463), .A2(new_n286), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n513), .A2(new_n230), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n502), .A2(new_n230), .A3(new_n206), .A4(new_n503), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n210), .B1(new_n412), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n258), .A2(new_n210), .A3(G68), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n391), .A2(new_n392), .B1(new_n502), .B2(new_n503), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n564), .B(new_n565), .C1(KEYINPUT19), .C2(new_n566), .ZN(new_n567));
  AOI211_X1 g0367(.A(new_n559), .B(new_n560), .C1(new_n567), .C2(new_n281), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n262), .A2(new_n264), .A3(G244), .A4(G1698), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n262), .A2(new_n264), .A3(G238), .A4(new_n298), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G116), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT82), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT82), .A4(new_n571), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n304), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n488), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n491), .B2(new_n231), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n310), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(G190), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n303), .B1(new_n572), .B2(new_n573), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(new_n575), .B1(new_n310), .B2(new_n578), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n568), .B(new_n580), .C1(new_n317), .C2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n576), .A2(new_n340), .A3(new_n579), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n567), .A2(new_n281), .ZN(new_n585));
  INV_X1    g0385(.A(new_n559), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n514), .A2(new_n463), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n584), .B(new_n588), .C1(G169), .C2(new_n582), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n558), .A2(new_n583), .A3(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n524), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n529), .A2(new_n539), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT24), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n529), .A2(new_n539), .A3(new_n540), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n389), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT85), .B1(new_n595), .B2(new_n548), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT85), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n543), .A2(new_n597), .A3(new_n549), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n554), .A2(G169), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n340), .B2(new_n554), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(G116), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n289), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n513), .B2(new_n602), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT20), .ZN(new_n605));
  AOI21_X1  g0405(.A(G33), .B1(new_n502), .B2(new_n503), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n484), .A2(new_n210), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n280), .A2(new_n221), .B1(G20), .B2(new_n602), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n605), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(KEYINPUT20), .B(new_n609), .C1(new_n606), .C2(new_n607), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n604), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n262), .A2(new_n264), .A3(G257), .A4(new_n298), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT83), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT83), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n258), .A2(new_n616), .A3(G257), .A4(new_n298), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n262), .A2(new_n264), .A3(G1698), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n619), .A2(G264), .B1(G303), .B2(new_n265), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n303), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n494), .A2(new_n308), .A3(G270), .A4(new_n309), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n490), .ZN(new_n623));
  NOR4_X1   g0423(.A1(new_n613), .A2(new_n621), .A3(new_n340), .A4(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n604), .ZN(new_n625));
  INV_X1    g0425(.A(new_n503), .ZN(new_n626));
  NOR2_X1   g0426(.A1(KEYINPUT80), .A2(G97), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n261), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(new_n210), .A3(new_n484), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT20), .B1(new_n629), .B2(new_n609), .ZN(new_n630));
  INV_X1    g0430(.A(new_n612), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n625), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G169), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n621), .A2(new_n623), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT21), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n618), .A2(new_n620), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n304), .ZN(new_n637));
  INV_X1    g0437(.A(new_n623), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT21), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n639), .A2(new_n640), .A3(G169), .A4(new_n632), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n624), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n632), .B1(new_n639), .B2(G200), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n323), .B2(new_n639), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n478), .A2(new_n591), .A3(new_n601), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g0447(.A(new_n647), .B(KEYINPUT86), .Z(G372));
  OAI21_X1  g0448(.A(KEYINPUT18), .B1(new_n355), .B2(new_n292), .ZN(new_n649));
  INV_X1    g0449(.A(new_n360), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n650), .A2(new_n334), .A3(new_n330), .A4(new_n344), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n441), .A2(new_n436), .A3(new_n421), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n471), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n451), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n332), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n404), .A2(new_n406), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n408), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT87), .B1(new_n524), .B2(new_n590), .ZN(new_n661));
  INV_X1    g0461(.A(new_n523), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n499), .A2(new_n317), .ZN(new_n663));
  OAI22_X1  g0463(.A1(new_n663), .A2(KEYINPUT81), .B1(new_n323), .B2(new_n496), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n496), .A2(new_n345), .B1(new_n510), .B2(new_n515), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n662), .A2(new_n664), .B1(new_n500), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n590), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT87), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n642), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n543), .A2(new_n549), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(new_n600), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n661), .B(new_n669), .C1(new_n670), .C2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n589), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n583), .A2(new_n589), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n517), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n497), .A2(new_n500), .A3(new_n516), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n678), .A2(KEYINPUT26), .A3(new_n589), .A4(new_n583), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n674), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n660), .B1(new_n477), .B2(new_n682), .ZN(G369));
  NAND3_X1  g0483(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n613), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n670), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n645), .B2(new_n691), .ZN(new_n693));
  XNOR2_X1  g0493(.A(KEYINPUT88), .B(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT89), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n601), .A2(new_n690), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n596), .A2(new_n598), .A3(new_n689), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n601), .A2(new_n699), .A3(new_n558), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n670), .A2(new_n690), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n700), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n672), .B2(new_n690), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT90), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT90), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n704), .A2(new_n710), .ZN(G399));
  NOR2_X1   g0511(.A1(new_n214), .A2(G41), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n209), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n561), .A2(G116), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n713), .A2(new_n714), .B1(new_n220), .B2(new_n712), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  NAND2_X1  g0516(.A1(new_n601), .A2(new_n642), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n666), .A3(new_n667), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n689), .B1(new_n680), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n681), .A2(new_n690), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(KEYINPUT29), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n591), .A2(new_n646), .A3(new_n601), .A4(new_n690), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n622), .A2(G179), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n554), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n582), .A2(new_n727), .A3(new_n499), .A4(new_n637), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT30), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n621), .A2(new_n554), .A3(new_n726), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(new_n499), .A4(new_n582), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n634), .A2(new_n582), .A3(G179), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n496), .A2(KEYINPUT91), .A3(new_n554), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT91), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n499), .B2(new_n555), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n690), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n733), .A2(KEYINPUT92), .A3(new_n738), .ZN(new_n743));
  AOI21_X1  g0543(.A(KEYINPUT92), .B1(new_n733), .B2(new_n738), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n743), .A2(new_n744), .A3(new_n690), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n725), .B(new_n742), .C1(new_n745), .C2(KEYINPUT31), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n746), .A2(new_n695), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n724), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n716), .B1(new_n750), .B2(G1), .ZN(G364));
  NAND2_X1  g0551(.A1(new_n210), .A2(G13), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT93), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G45), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n713), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n697), .B(new_n755), .C1(new_n695), .C2(new_n693), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n756), .A2(KEYINPUT94), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(KEYINPUT94), .ZN(new_n758));
  INV_X1    g0558(.A(new_n755), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n213), .A2(new_n258), .ZN(new_n760));
  INV_X1    g0560(.A(G355), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n761), .B1(G116), .B2(new_n213), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n214), .A2(new_n258), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n487), .B2(new_n220), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n253), .A2(new_n487), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT95), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n221), .B1(G20), .B2(new_n345), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n759), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G283), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n210), .A2(G179), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(new_n323), .A3(G200), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n776), .A2(G190), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(G303), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n775), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n210), .A2(new_n340), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G190), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n317), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G326), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n782), .A2(G200), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n780), .B(new_n786), .C1(G322), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G190), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n781), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n781), .A2(new_n323), .A3(G200), .ZN(new_n792));
  XOR2_X1   g0592(.A(KEYINPUT33), .B(G317), .Z(new_n793));
  OAI221_X1 g0593(.A(new_n265), .B1(new_n790), .B2(new_n791), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G179), .A2(G200), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT96), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n796), .A2(G20), .A3(new_n323), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n794), .B1(G329), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G294), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n210), .B1(new_n796), .B2(G190), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT98), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(KEYINPUT98), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n788), .B(new_n799), .C1(new_n800), .C2(new_n804), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT99), .ZN(new_n806));
  INV_X1    g0606(.A(new_n787), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n807), .A2(new_n234), .B1(new_n784), .B2(new_n202), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n258), .B1(new_n790), .B2(new_n371), .C1(new_n228), .C2(new_n792), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n777), .A2(new_n206), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n778), .A2(new_n230), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G159), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n797), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(KEYINPUT97), .B(KEYINPUT32), .Z(new_n815));
  XNOR2_X1  g0615(.A(new_n814), .B(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n812), .B(new_n816), .C1(new_n205), .C2(new_n804), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n805), .A2(KEYINPUT99), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n806), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n774), .B1(new_n819), .B2(new_n771), .ZN(new_n820));
  INV_X1    g0620(.A(new_n770), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n693), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT100), .ZN(new_n823));
  AND3_X1   g0623(.A1(new_n757), .A2(new_n758), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NOR2_X1   g0625(.A1(new_n472), .A2(new_n689), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n474), .B1(new_n469), .B2(new_n690), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n472), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n722), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n826), .B1(new_n472), .B2(new_n828), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n681), .A2(new_n690), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n759), .B1(new_n834), .B2(new_n748), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n748), .B2(new_n834), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n771), .A2(new_n768), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n755), .B1(new_n371), .B2(new_n837), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n265), .B1(new_n790), .B2(new_n602), .C1(new_n775), .C2(new_n792), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n787), .A2(G294), .B1(new_n783), .B2(G303), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n840), .B1(new_n230), .B2(new_n777), .C1(new_n206), .C2(new_n778), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n839), .B(new_n841), .C1(G311), .C2(new_n798), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n205), .B2(new_n804), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n798), .A2(G132), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n258), .B1(new_n778), .B2(new_n202), .C1(new_n228), .C2(new_n777), .ZN(new_n845));
  INV_X1    g0645(.A(new_n792), .ZN(new_n846));
  INV_X1    g0646(.A(new_n790), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n846), .A2(G150), .B1(new_n847), .B2(G159), .ZN(new_n848));
  INV_X1    g0648(.A(G143), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n848), .B1(new_n807), .B2(new_n849), .C1(new_n850), .C2(new_n784), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n844), .B(new_n845), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n853), .B1(new_n852), .B2(new_n851), .C1(new_n234), .C2(new_n804), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n843), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n771), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n838), .B1(new_n855), .B2(new_n856), .C1(new_n832), .C2(new_n769), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n836), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(G384));
  INV_X1    g0659(.A(KEYINPUT105), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT92), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n739), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n733), .A2(KEYINPUT92), .A3(new_n738), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n862), .A2(new_n741), .A3(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n725), .B(new_n864), .C1(new_n745), .C2(KEYINPUT31), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n445), .A2(new_n689), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n451), .A2(new_n653), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n449), .A2(new_n450), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n444), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n867), .B1(new_n869), .B2(new_n866), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n865), .A2(new_n832), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n366), .A2(KEYINPUT102), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT102), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n357), .A2(new_n873), .A3(new_n358), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n292), .A2(new_n325), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  INV_X1    g0676(.A(new_n687), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n330), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n872), .A2(new_n874), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n878), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n355), .A2(new_n292), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n369), .B2(new_n878), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT38), .B(new_n884), .C1(new_n369), .C2(new_n878), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n871), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n860), .B1(new_n889), .B2(KEYINPUT40), .ZN(new_n890));
  INV_X1    g0690(.A(new_n871), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n367), .A2(KEYINPUT79), .A3(new_n363), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT79), .B1(new_n367), .B2(new_n363), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n656), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n878), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n896), .B2(new_n884), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n875), .A2(new_n878), .ZN(new_n898));
  INV_X1    g0698(.A(new_n882), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n876), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(KEYINPUT102), .B2(new_n366), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n900), .B1(new_n874), .B2(new_n902), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n886), .B(new_n903), .C1(new_n894), .C2(new_n895), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n891), .B1(new_n897), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(KEYINPUT105), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n880), .A2(KEYINPUT103), .A3(new_n883), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n649), .A2(new_n651), .A3(new_n331), .A4(new_n326), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n895), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT104), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n909), .A2(KEYINPUT104), .A3(new_n895), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n908), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT103), .B1(new_n880), .B2(new_n883), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n886), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n888), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n871), .A2(new_n906), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n890), .A2(new_n907), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n862), .A2(new_n689), .A3(new_n863), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n743), .A2(new_n744), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n740), .A2(new_n920), .B1(new_n921), .B2(new_n741), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n477), .B1(new_n725), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n695), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n919), .B2(new_n923), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n917), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n451), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n690), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n887), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n927), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n887), .A2(new_n888), .ZN(new_n933));
  INV_X1    g0733(.A(new_n870), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n833), .B2(new_n827), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n933), .A2(new_n935), .B1(new_n652), .B2(new_n687), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n659), .B1(new_n723), .B2(new_n478), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n937), .B(new_n938), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n925), .A2(new_n939), .B1(new_n209), .B2(new_n753), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n939), .B2(new_n925), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n219), .A2(new_n371), .A3(new_n268), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n202), .A2(G68), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n209), .B(G13), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n504), .A2(new_n506), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT35), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT35), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n946), .A2(G116), .A3(new_n222), .A4(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(KEYINPUT101), .B(KEYINPUT36), .Z(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  OR3_X1    g0750(.A1(new_n941), .A2(new_n944), .A3(new_n950), .ZN(G367));
  NAND2_X1  g0751(.A1(new_n516), .A2(new_n689), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n666), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n678), .A2(new_n689), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT107), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n954), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT107), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n703), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(KEYINPUT109), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n601), .B1(new_n956), .B2(new_n959), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n690), .B1(new_n963), .B2(new_n678), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n706), .ZN(new_n966));
  OR3_X1    g0766(.A1(new_n966), .A2(new_n955), .A3(KEYINPUT42), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT42), .B1(new_n966), .B2(new_n955), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT108), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT108), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n964), .A2(new_n971), .A3(new_n968), .A4(new_n967), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n568), .A2(new_n690), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n674), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT106), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(new_n676), .C2(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n975), .B2(new_n974), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT43), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n970), .A2(new_n972), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n970), .A2(new_n972), .B1(new_n978), .B2(new_n977), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n962), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n961), .A2(KEYINPUT109), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n970), .A2(new_n972), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n977), .A2(new_n978), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n980), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n990), .A2(new_n962), .A3(new_n984), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n712), .B(KEYINPUT41), .Z(new_n992));
  AOI21_X1  g0792(.A(new_n955), .B1(new_n708), .B2(new_n709), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT45), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n708), .A2(new_n709), .A3(new_n955), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT44), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n703), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n706), .B1(new_n702), .B2(new_n705), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n697), .B(new_n1000), .Z(new_n1001));
  NOR2_X1   g0801(.A1(new_n1001), .A2(new_n749), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n994), .A2(new_n997), .A3(new_n704), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n999), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n992), .B1(new_n1004), .B2(new_n750), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n754), .A2(G1), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n986), .B(new_n991), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n258), .B1(new_n790), .B2(new_n202), .C1(new_n813), .C2(new_n792), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n777), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n787), .A2(G150), .B1(new_n1009), .B2(G77), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n234), .B2(new_n778), .C1(new_n849), .C2(new_n784), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1008), .B(new_n1011), .C1(G137), .C2(new_n798), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n804), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(G68), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n804), .A2(new_n206), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT46), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n778), .A2(new_n1017), .A3(new_n602), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n265), .B1(new_n790), .B2(new_n775), .C1(new_n800), .C2(new_n792), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(G317), .C2(new_n798), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n807), .A2(new_n779), .B1(new_n784), .B2(new_n791), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n502), .A2(new_n503), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1021), .B1(new_n1022), .B2(new_n1009), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1017), .B1(new_n778), .B2(new_n602), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT110), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1020), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1015), .B1(new_n1016), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT47), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n771), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n977), .A2(new_n770), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n773), .B1(new_n214), .B2(new_n463), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n249), .A2(new_n763), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n755), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n1029), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1007), .A2(new_n1035), .ZN(G387));
  INV_X1    g0836(.A(new_n1002), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1001), .A2(new_n749), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n712), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n763), .B1(new_n245), .B2(new_n487), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n714), .B2(new_n760), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n283), .A2(new_n202), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT111), .Z(new_n1043));
  OR2_X1    g0843(.A1(new_n1043), .A2(KEYINPUT50), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g0845(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1044), .A2(new_n714), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1041), .A2(new_n1047), .B1(new_n206), .B2(new_n214), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n759), .B1(new_n1048), .B2(new_n773), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n258), .B1(new_n790), .B2(new_n228), .C1(new_n290), .C2(new_n792), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n787), .A2(G50), .B1(new_n1009), .B2(G97), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n371), .B2(new_n778), .C1(new_n813), .C2(new_n784), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(G150), .C2(new_n798), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1013), .A2(new_n463), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n846), .A2(G311), .B1(new_n847), .B2(G303), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n787), .A2(G317), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n783), .A2(G322), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT48), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n775), .B2(new_n804), .C1(new_n800), .C2(new_n778), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT49), .Z(new_n1062));
  OAI221_X1 g0862(.A(new_n265), .B1(new_n602), .B2(new_n777), .C1(new_n797), .C2(new_n785), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1055), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1049), .B1(new_n1064), .B2(new_n771), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n701), .B2(new_n821), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1006), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1039), .B(new_n1066), .C1(new_n1067), .C2(new_n1001), .ZN(G393));
  AND3_X1   g0868(.A1(new_n994), .A2(new_n997), .A3(new_n704), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n704), .B1(new_n994), .B2(new_n997), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1037), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n1004), .A3(new_n712), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1067), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1022), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n772), .B1(new_n213), .B2(new_n1074), .C1(new_n764), .C2(new_n256), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT112), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n755), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n1076), .B2(new_n1075), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n787), .A2(G311), .B1(new_n783), .B2(G317), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT52), .Z(new_n1080));
  OAI22_X1  g0880(.A1(new_n206), .A2(new_n777), .B1(new_n778), .B2(new_n775), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n265), .B1(new_n790), .B2(new_n800), .C1(new_n779), .C2(new_n792), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(G322), .C2(new_n798), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1080), .B(new_n1083), .C1(new_n602), .C2(new_n804), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1013), .A2(G77), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n202), .B2(new_n792), .C1(new_n290), .C2(new_n790), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT113), .Z(new_n1087));
  AOI22_X1  g0887(.A1(new_n787), .A2(G159), .B1(new_n783), .B2(G150), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT51), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n265), .B1(new_n1009), .B2(G87), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n228), .B2(new_n778), .C1(new_n797), .C2(new_n849), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1084), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1078), .B1(new_n1093), .B2(new_n771), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n960), .B2(new_n821), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1073), .A2(KEYINPUT114), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT114), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n999), .A2(new_n1006), .A3(new_n1003), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n1095), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1072), .B1(new_n1097), .B2(new_n1100), .ZN(G390));
  INV_X1    g0901(.A(KEYINPUT116), .ZN(new_n1102));
  INV_X1    g0902(.A(G330), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n830), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n865), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1102), .B1(new_n1105), .B2(new_n934), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n865), .A2(new_n1104), .A3(KEYINPUT116), .A4(new_n870), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n935), .A2(new_n930), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n927), .B2(new_n931), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n680), .A2(new_n718), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(new_n690), .A3(new_n829), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n827), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(KEYINPUT115), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT115), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(new_n1115), .A3(new_n827), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1114), .A2(new_n870), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n917), .A2(new_n1117), .A3(new_n929), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1108), .B1(new_n1110), .B2(new_n1119), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n935), .A2(new_n930), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n887), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n1122));
  AOI21_X1  g0922(.A(KEYINPUT39), .B1(new_n916), .B2(new_n888), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n746), .A2(new_n695), .A3(new_n832), .A4(new_n870), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n1118), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1120), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n865), .A2(new_n369), .A3(new_n476), .A4(G330), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT117), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n938), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n832), .A2(G330), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n922), .B2(new_n725), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1125), .B1(new_n1133), .B2(new_n870), .ZN(new_n1134));
  AOI211_X1 g0934(.A(KEYINPUT115), .B(new_n826), .C1(new_n719), .C2(new_n829), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1115), .B1(new_n1112), .B2(new_n827), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT118), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT118), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1105), .A2(new_n934), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1125), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n746), .A2(new_n695), .A3(new_n832), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n934), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1106), .A2(new_n1145), .A3(new_n1107), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n833), .A2(new_n827), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1131), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1127), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1120), .A2(new_n1126), .A3(new_n1149), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n712), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1120), .A2(new_n1126), .A3(new_n1006), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n258), .B1(new_n790), .B2(new_n1155), .C1(new_n850), .C2(new_n792), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n787), .A2(G132), .B1(new_n783), .B2(G128), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n202), .B2(new_n777), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1156), .B(new_n1158), .C1(G125), .C2(new_n798), .ZN(new_n1159));
  INV_X1    g0959(.A(G150), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n778), .A2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT53), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1159), .B(new_n1162), .C1(new_n813), .C2(new_n804), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n811), .B1(G68), .B2(new_n1009), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n787), .A2(G116), .B1(new_n783), .B2(G283), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n265), .B1(new_n792), .B2(new_n206), .C1(new_n1074), .C2(new_n790), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G294), .B2(new_n798), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1085), .A2(new_n1164), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n856), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n755), .B(new_n1169), .C1(new_n290), .C2(new_n837), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(new_n769), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1153), .A2(new_n1154), .A3(new_n1172), .ZN(G378));
  NOR2_X1   g0973(.A1(new_n402), .A2(new_n687), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT120), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n409), .B(new_n1175), .ZN(new_n1176));
  XOR2_X1   g0976(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1177));
  XNOR2_X1  g0977(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n890), .A2(new_n907), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1103), .B1(new_n917), .B2(new_n918), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1180), .A2(new_n937), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n937), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1179), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(KEYINPUT105), .B1(new_n905), .B2(new_n906), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n889), .A2(new_n860), .A3(KEYINPUT40), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1181), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n937), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1180), .A2(new_n937), .A3(new_n1181), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(new_n1178), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1184), .A2(new_n1006), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n837), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n759), .B1(G50), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n258), .A2(G41), .ZN(new_n1195));
  INV_X1    g0995(.A(G41), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G50), .B(new_n1195), .C1(new_n261), .C2(new_n1196), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n784), .A2(new_n602), .B1(new_n778), .B2(new_n371), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n807), .A2(new_n206), .B1(new_n777), .B2(new_n234), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1195), .B1(new_n790), .B2(new_n462), .C1(new_n205), .C2(new_n792), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G283), .B2(new_n798), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1014), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  XOR2_X1   g1003(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1204));
  AOI21_X1  g1004(.A(new_n1197), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1013), .A2(G150), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n778), .A2(new_n1155), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n846), .A2(G132), .B1(new_n847), .B2(G137), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n787), .A2(G128), .B1(new_n783), .B2(G125), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n261), .B(new_n1196), .C1(new_n777), .C2(new_n813), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n798), .B2(G124), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1205), .B1(new_n1204), .B2(new_n1203), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1194), .B1(new_n1216), .B2(new_n771), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1178), .B2(new_n769), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1192), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1131), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1152), .A2(new_n1220), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1184), .A2(new_n1191), .A3(KEYINPUT57), .A4(new_n1221), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1222), .A2(new_n712), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1184), .A2(new_n1221), .A3(new_n1191), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT57), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1219), .B1(new_n1223), .B2(new_n1226), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT121), .Z(G375));
  INV_X1    g1028(.A(new_n992), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1143), .A2(new_n1131), .A3(new_n1148), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1150), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n265), .B1(new_n790), .B2(new_n206), .C1(new_n602), .C2(new_n792), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n787), .A2(G283), .B1(new_n783), .B2(G294), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n371), .B2(new_n777), .C1(new_n205), .C2(new_n778), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1232), .B(new_n1234), .C1(G303), .C2(new_n798), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n258), .B1(new_n790), .B2(new_n1160), .C1(new_n792), .C2(new_n1155), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n787), .A2(G137), .B1(new_n783), .B2(G132), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1237), .B1(new_n234), .B2(new_n777), .C1(new_n813), .C2(new_n778), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1236), .B(new_n1238), .C1(G128), .C2(new_n798), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1013), .A2(G50), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1054), .A2(new_n1235), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n759), .B1(G68), .B2(new_n1193), .C1(new_n1241), .C2(new_n856), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n934), .B2(new_n768), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1143), .A2(new_n1148), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(new_n1006), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1231), .A2(new_n1245), .ZN(G381));
  OR3_X1    g1046(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1247));
  OR4_X1    g1047(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1247), .ZN(new_n1248));
  OR3_X1    g1048(.A1(G375), .A2(new_n1248), .A3(G378), .ZN(G407));
  INV_X1    g1049(.A(G378), .ZN(new_n1250));
  INV_X1    g1050(.A(G213), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1251), .A2(G343), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G407), .B(G213), .C1(G375), .C2(new_n1253), .ZN(G409));
  AND2_X1   g1054(.A1(new_n1192), .A2(new_n1218), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1222), .A2(new_n712), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G378), .B(new_n1255), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1184), .A2(new_n1191), .A3(new_n1229), .A4(new_n1221), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(new_n1192), .A3(new_n1218), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1250), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1252), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT122), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1138), .A2(new_n1142), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n712), .B1(new_n1265), .B2(new_n1131), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT60), .B1(new_n1265), .B2(new_n1131), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1265), .A2(KEYINPUT60), .A3(new_n1131), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1264), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n712), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1244), .B2(new_n1220), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1230), .A2(new_n1273), .ZN(new_n1274));
  AND4_X1   g1074(.A1(new_n1264), .A2(new_n1272), .A3(new_n1269), .A4(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1245), .B1(new_n1270), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n858), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G384), .B(new_n1245), .C1(new_n1270), .C2(new_n1275), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1262), .A2(new_n1263), .A3(new_n1279), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(KEYINPUT62), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT124), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1277), .A2(new_n1282), .A3(new_n1278), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1252), .A2(G2897), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1283), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1279), .A2(new_n1282), .A3(new_n1285), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1260), .A2(new_n1250), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1227), .B2(G378), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1287), .B(new_n1288), .C1(new_n1290), .C2(new_n1252), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT61), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT114), .B1(new_n1073), .B2(new_n1096), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1099), .A2(new_n1098), .A3(new_n1095), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1069), .A2(new_n1070), .A3(new_n1037), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1296), .A2(new_n1271), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n1294), .A2(new_n1295), .B1(new_n1297), .B2(new_n1071), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n986), .A2(new_n991), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1229), .B1(new_n1296), .B2(new_n749), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(new_n1067), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1298), .B1(new_n1301), .B2(new_n1034), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(G393), .B(new_n824), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(G390), .A2(new_n1007), .A3(new_n1035), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1302), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1303), .B1(new_n1302), .B2(new_n1304), .ZN(new_n1306));
  OAI22_X1  g1106(.A1(new_n1281), .A2(new_n1293), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT125), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1262), .A2(KEYINPUT63), .A3(new_n1263), .A4(new_n1279), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1291), .A2(new_n1292), .A3(new_n1309), .A4(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT123), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1280), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1313), .B1(new_n1280), .B2(new_n1314), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1308), .B1(new_n1312), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1319));
  AOI211_X1 g1119(.A(new_n1252), .B(new_n1319), .C1(new_n1258), .C2(new_n1261), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT123), .B1(new_n1320), .B2(KEYINPUT63), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1280), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(new_n1323), .A2(new_n1311), .A3(KEYINPUT125), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1307), .B1(new_n1318), .B2(new_n1324), .ZN(G405));
  OAI21_X1  g1125(.A(new_n1319), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1303), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1302), .A2(new_n1304), .A3(new_n1303), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1329), .A2(new_n1279), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1326), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1332), .B(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT126), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(G375), .A2(new_n1335), .A3(new_n1250), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(G375), .A2(new_n1250), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1258), .A2(new_n1335), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1334), .A2(new_n1336), .A3(new_n1339), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1332), .B(KEYINPUT127), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1339), .A2(new_n1336), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1340), .A2(new_n1343), .ZN(G402));
endmodule


