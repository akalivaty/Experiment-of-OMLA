//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n558, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(KEYINPUT65), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(G125), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n458), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n458), .A2(G101), .A3(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n459), .A2(G137), .A3(new_n458), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G112), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G2105), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n459), .A2(KEYINPUT67), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n459), .A2(KEYINPUT67), .ZN(new_n478));
  OAI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n476), .B1(new_n480), .B2(G124), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n458), .B1(new_n477), .B2(new_n478), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT68), .B(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(new_n458), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n491), .A2(KEYINPUT68), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(KEYINPUT68), .ZN(new_n493));
  OAI211_X1 g068(.A(KEYINPUT69), .B(G2105), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n487), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n459), .A2(KEYINPUT4), .A3(G138), .A4(new_n458), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n459), .A2(G126), .A3(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n461), .A2(G138), .A3(new_n458), .A4(new_n464), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT70), .B1(new_n506), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n509), .B2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(new_n506), .A3(G543), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n507), .A2(new_n510), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n505), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n507), .A2(new_n510), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n511), .A2(new_n513), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n517), .A2(new_n518), .A3(new_n505), .A4(new_n515), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n517), .A2(new_n518), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n515), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(G651), .B1(G50), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n522), .A2(new_n529), .ZN(G166));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n534), .B1(new_n514), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n517), .A2(new_n518), .A3(new_n515), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n538), .A2(G89), .A3(new_n519), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  NAND3_X1  g116(.A1(new_n517), .A2(new_n518), .A3(G64), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n544), .A2(G651), .B1(G52), .B2(new_n528), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n538), .A2(G90), .A3(new_n519), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND3_X1  g123(.A1(new_n517), .A2(new_n518), .A3(G56), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G651), .B1(G43), .B2(new_n528), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n538), .A2(G81), .A3(new_n519), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  XOR2_X1   g132(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n558));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n524), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n515), .A2(G53), .A3(G543), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n569), .B1(new_n516), .B2(new_n520), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n538), .A2(KEYINPUT74), .A3(new_n519), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n568), .B1(new_n572), .B2(G91), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G299));
  NAND2_X1  g149(.A1(new_n522), .A2(new_n529), .ZN(G303));
  NAND2_X1  g150(.A1(new_n572), .A2(G87), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  INV_X1    g152(.A(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n527), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n528), .A2(KEYINPUT75), .A3(G49), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n514), .A2(G74), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n579), .A2(new_n580), .B1(new_n581), .B2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n576), .A2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n524), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  INV_X1    g162(.A(G48), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT76), .B1(new_n527), .B2(new_n588), .ZN(new_n589));
  OR3_X1    g164(.A1(new_n527), .A2(KEYINPUT76), .A3(new_n588), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  AND3_X1   g167(.A1(new_n538), .A2(KEYINPUT74), .A3(new_n519), .ZN(new_n593));
  AOI21_X1  g168(.A(KEYINPUT74), .B1(new_n538), .B2(new_n519), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G60), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n524), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(G47), .B2(new_n528), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n538), .A2(G85), .A3(new_n519), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT77), .Z(new_n605));
  NAND2_X1  g180(.A1(new_n528), .A2(G54), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n517), .A2(new_n518), .A3(G66), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT78), .Z(new_n609));
  NOR2_X1   g184(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G651), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n606), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(new_n570), .B2(new_n571), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(G92), .B1(new_n593), .B2(new_n594), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(KEYINPUT10), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n605), .B1(G868), .B2(new_n620), .ZN(G284));
  OAI21_X1  g196(.A(new_n605), .B1(G868), .B2(new_n620), .ZN(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n573), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n623), .B1(new_n573), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n620), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n552), .A2(new_n553), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n618), .A2(KEYINPUT10), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n572), .A2(new_n616), .A3(G92), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n629), .A2(new_n626), .A3(new_n630), .A4(new_n613), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT79), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n612), .B1(new_n618), .B2(KEYINPUT10), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT79), .ZN(new_n634));
  NAND4_X1  g209(.A1(new_n633), .A2(new_n634), .A3(new_n626), .A4(new_n630), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  MUX2_X1   g211(.A(new_n628), .B(new_n636), .S(G868), .Z(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g213(.A1(new_n461), .A2(new_n464), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n639), .A2(G2104), .A3(new_n458), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT12), .Z(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT13), .Z(new_n642));
  INV_X1    g217(.A(G2100), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n483), .A2(G135), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n480), .A2(G123), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n458), .A2(G111), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n646), .B(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2096), .Z(new_n651));
  NAND3_X1  g226(.A1(new_n644), .A2(new_n645), .A3(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT80), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2430), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n661), .B(new_n662), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n659), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(G14), .B1(new_n664), .B2(new_n666), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  AOI21_X1  g249(.A(KEYINPUT18), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n675), .B(new_n677), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2096), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT81), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(KEYINPUT82), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  OR3_X1    g263(.A1(new_n682), .A2(new_n683), .A3(KEYINPUT82), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n682), .A2(new_n683), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n684), .A2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(new_n694), .B(new_n693), .S(new_n688), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(G229));
  NAND2_X1  g279(.A1(new_n620), .A2(G16), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G4), .B2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G1348), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n639), .A2(G127), .ZN(new_n709));
  NAND2_X1  g284(.A1(G115), .A2(G2104), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n458), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT25), .Z(new_n713));
  INV_X1    g288(.A(G139), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n482), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G29), .ZN(new_n717));
  NOR2_X1   g292(.A1(G29), .A2(G33), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT94), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT95), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(G2072), .Z(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G35), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G162), .B2(new_n723), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT29), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(G2090), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n722), .B1(KEYINPUT99), .B2(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(KEYINPUT99), .ZN(new_n729));
  OR2_X1    g304(.A1(G104), .A2(G2105), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n730), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT92), .Z(new_n732));
  INV_X1    g307(.A(G140), .ZN(new_n733));
  INV_X1    g308(.A(G128), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n732), .B1(new_n482), .B2(new_n733), .C1(new_n734), .C2(new_n479), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G29), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT93), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n723), .A2(G26), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G2067), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  AND4_X1   g317(.A1(new_n708), .A2(new_n728), .A3(new_n729), .A4(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G20), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT23), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n573), .B2(new_n744), .ZN(new_n747));
  INV_X1    g322(.A(G1956), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G2078), .ZN(new_n750));
  NAND2_X1  g325(.A1(G164), .A2(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G27), .B2(G29), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT26), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n458), .A2(G2104), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n755), .A2(new_n756), .B1(G105), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G141), .ZN(new_n759));
  INV_X1    g334(.A(G129), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n758), .B1(new_n482), .B2(new_n759), .C1(new_n760), .C2(new_n479), .ZN(new_n761));
  MUX2_X1   g336(.A(G32), .B(new_n761), .S(G29), .Z(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT27), .B(G1996), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n750), .A2(new_n752), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  NAND2_X1  g341(.A1(G160), .A2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n723), .B1(new_n768), .B2(G34), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n769), .A2(KEYINPUT97), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(G34), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n769), .B2(KEYINPUT97), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n767), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n765), .B1(new_n750), .B2(new_n752), .C1(new_n766), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G2090), .B2(new_n726), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n762), .A2(new_n764), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT98), .Z(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  NOR2_X1   g353(.A1(G171), .A2(new_n744), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G5), .B2(new_n744), .ZN(new_n780));
  NOR2_X1   g355(.A1(G168), .A2(new_n744), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n744), .B2(G21), .ZN(new_n782));
  INV_X1    g357(.A(G1966), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n778), .A2(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n778), .B2(new_n780), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT30), .B(G28), .ZN(new_n786));
  OR2_X1    g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  NAND2_X1  g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n786), .A2(new_n723), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n650), .B2(new_n723), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n766), .B2(new_n773), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n783), .B2(new_n782), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n744), .A2(G19), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n554), .B2(new_n744), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1341), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n785), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  AND4_X1   g371(.A1(new_n749), .A2(new_n775), .A3(new_n777), .A4(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n706), .A2(new_n707), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n743), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n744), .A2(G22), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G166), .B2(new_n744), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1971), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT33), .B(G1976), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT89), .ZN(new_n804));
  NOR2_X1   g379(.A1(G16), .A2(G23), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT88), .Z(new_n806));
  AND2_X1   g381(.A1(new_n576), .A2(new_n582), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G16), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n802), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n744), .A2(G6), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n591), .B1(new_n572), .B2(G86), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n744), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT32), .B(G1981), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n808), .A2(new_n804), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n809), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT90), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT34), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n723), .A2(G25), .ZN(new_n823));
  OR2_X1    g398(.A1(G95), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n825));
  INV_X1    g400(.A(G119), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n479), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G131), .B2(new_n483), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT84), .Z(new_n829));
  OAI21_X1  g404(.A(new_n823), .B1(new_n829), .B2(new_n723), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT85), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(KEYINPUT85), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G1991), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n744), .A2(G24), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT86), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(G290), .B2(G16), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT87), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G1986), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n834), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n831), .A2(new_n842), .A3(new_n832), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n835), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n818), .A2(KEYINPUT34), .A3(new_n819), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n822), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT91), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT36), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n844), .B1(new_n820), .B2(new_n821), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n852), .A2(new_n849), .A3(new_n846), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n799), .B1(new_n851), .B2(new_n853), .ZN(G311));
  INV_X1    g429(.A(new_n799), .ZN(new_n855));
  INV_X1    g430(.A(new_n853), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n849), .B1(new_n852), .B2(new_n846), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(G150));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n538), .A2(G93), .A3(new_n519), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n515), .A2(G55), .A3(G543), .ZN(new_n861));
  NAND2_X1  g436(.A1(G80), .A2(G543), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n514), .B2(G67), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n861), .B1(new_n864), .B2(new_n611), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n859), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n861), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n517), .A2(new_n518), .A3(G67), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n862), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n867), .B1(new_n869), .B2(G651), .ZN(new_n870));
  INV_X1    g445(.A(G93), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n538), .A2(new_n519), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n870), .B(KEYINPUT100), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n866), .A2(new_n628), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n860), .A2(new_n865), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n554), .A2(new_n875), .A3(KEYINPUT100), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n620), .A2(G559), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n881));
  AOI21_X1  g456(.A(G860), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n881), .B2(new_n880), .ZN(new_n883));
  INV_X1    g458(.A(new_n875), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G860), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT37), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT101), .ZN(G145));
  XNOR2_X1  g463(.A(G162), .B(new_n650), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(G160), .ZN(new_n890));
  OR2_X1    g465(.A1(G106), .A2(G2105), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n891), .B(G2104), .C1(G118), .C2(new_n458), .ZN(new_n892));
  INV_X1    g467(.A(G142), .ZN(new_n893));
  INV_X1    g468(.A(G130), .ZN(new_n894));
  OAI221_X1 g469(.A(new_n892), .B1(new_n482), .B2(new_n893), .C1(new_n894), .C2(new_n479), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT102), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n641), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n829), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n898), .A2(KEYINPUT103), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n735), .B(new_n503), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n761), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n716), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(KEYINPUT103), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n899), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n899), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n890), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n899), .A2(new_n902), .A3(new_n903), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n902), .A2(new_n898), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(new_n890), .ZN(new_n909));
  AOI21_X1  g484(.A(G37), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n906), .A2(new_n910), .A3(KEYINPUT40), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT40), .B1(new_n906), .B2(new_n910), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(G395));
  NAND2_X1  g488(.A1(G305), .A2(G166), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n915));
  NAND2_X1  g490(.A1(G290), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n601), .A2(KEYINPUT107), .A3(new_n602), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n807), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n811), .A2(G303), .ZN(new_n920));
  NAND3_X1  g495(.A1(G288), .A2(new_n916), .A3(new_n917), .ZN(new_n921));
  AND4_X1   g496(.A1(new_n914), .A2(new_n919), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n919), .A2(new_n921), .B1(new_n914), .B2(new_n920), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n925));
  AND4_X1   g500(.A1(new_n573), .A2(new_n629), .A3(new_n630), .A4(new_n613), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n573), .B1(new_n633), .B2(new_n630), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(G299), .B1(new_n617), .B2(new_n619), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n633), .A2(new_n573), .A3(new_n630), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT104), .ZN(new_n931));
  INV_X1    g506(.A(new_n877), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n632), .A2(new_n635), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n632), .B2(new_n635), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n928), .B(new_n931), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  XOR2_X1   g510(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(new_n926), .B2(new_n927), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n929), .A2(new_n930), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n632), .A2(new_n635), .A3(new_n932), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n636), .A2(new_n877), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n935), .A2(new_n944), .A3(KEYINPUT105), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n942), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n928), .A4(new_n931), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n946), .B1(new_n945), .B2(new_n949), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n924), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n945), .A2(new_n949), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n922), .A2(new_n923), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n952), .A2(new_n957), .A3(G868), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n959));
  INV_X1    g534(.A(G868), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n884), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n952), .A2(new_n957), .A3(new_n959), .A4(G868), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(G295));
  AND2_X1   g539(.A1(new_n962), .A2(new_n963), .ZN(G331));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n966));
  NAND2_X1  g541(.A1(G171), .A2(G168), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n546), .A2(new_n545), .B1(new_n536), .B2(new_n539), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n877), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n874), .A2(new_n876), .A3(new_n967), .A4(new_n969), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(KEYINPUT110), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n974));
  AND4_X1   g549(.A1(new_n539), .A2(new_n545), .A3(new_n536), .A4(new_n546), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(new_n968), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n932), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n929), .A2(new_n930), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n972), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n976), .A2(KEYINPUT109), .A3(new_n876), .A4(new_n874), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n984), .A3(new_n971), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n929), .A2(new_n930), .A3(new_n939), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n936), .B1(new_n929), .B2(new_n930), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n981), .A2(new_n988), .A3(new_n955), .ZN(new_n989));
  INV_X1    g564(.A(G37), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n971), .A2(new_n984), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n992), .A2(new_n928), .A3(new_n931), .A4(new_n983), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n939), .B1(new_n926), .B2(new_n927), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n929), .A2(new_n930), .A3(new_n937), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n994), .A2(new_n973), .A3(new_n977), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n955), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT111), .B(KEYINPUT43), .C1(new_n991), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n993), .A2(new_n996), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n924), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(new_n990), .A3(new_n989), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT111), .B1(new_n1002), .B2(KEYINPUT43), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n983), .A2(new_n992), .B1(new_n938), .B2(new_n940), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n979), .B1(new_n973), .B2(new_n977), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n924), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n990), .A4(new_n989), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT44), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n999), .A2(new_n1003), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1006), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT43), .B1(new_n1011), .B2(new_n991), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1001), .A2(new_n1007), .A3(new_n990), .A4(new_n989), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT44), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n966), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(KEYINPUT44), .A3(new_n998), .A4(new_n1008), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1014), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(KEYINPUT112), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1015), .A2(new_n1021), .ZN(G397));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT116), .B(G1981), .Z(new_n1024));
  NOR2_X1   g599(.A1(G305), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1981), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n521), .A2(G86), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n592), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1023), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT49), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1023), .B(new_n1031), .C1(new_n1025), .C2(new_n1028), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1384), .B1(new_n499), .B2(new_n502), .ZN(new_n1033));
  INV_X1    g608(.A(G40), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n467), .A2(new_n1034), .A3(new_n472), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1030), .A2(new_n1032), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n576), .A2(G1976), .A3(new_n582), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1043), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1040), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G303), .A2(G8), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(KEYINPUT55), .ZN(new_n1050));
  INV_X1    g625(.A(G1971), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G160), .A2(G40), .ZN(new_n1052));
  INV_X1    g627(.A(G1384), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n503), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT45), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT113), .B(G1384), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1033), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1035), .B1(new_n1033), .B2(new_n1060), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G2090), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1051), .A2(new_n1059), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1050), .B1(new_n1066), .B2(new_n1038), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT119), .B1(new_n1048), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1040), .A2(new_n1067), .A3(new_n1070), .A4(new_n1047), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1050), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1971), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1054), .A2(KEYINPUT50), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(new_n1035), .A3(new_n1061), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(G2090), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1072), .B(G8), .C1(new_n1073), .C2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1035), .B1(new_n1033), .B2(KEYINPUT45), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n783), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1074), .A2(new_n766), .A3(new_n1035), .A4(new_n1061), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(G8), .A3(G168), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT63), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1069), .A2(new_n1071), .A3(new_n1077), .A4(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1040), .A2(new_n1077), .A3(new_n1067), .A4(new_n1047), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT118), .B1(new_n1087), .B2(new_n1083), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n1084), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1087), .A2(KEYINPUT118), .A3(new_n1083), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1086), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1048), .A2(new_n1077), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1040), .A2(new_n1045), .A3(new_n807), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(G305), .B2(new_n1024), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1092), .B1(new_n1094), .B2(new_n1039), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1080), .A2(new_n1081), .A3(G168), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G8), .ZN(new_n1097));
  AOI21_X1  g672(.A(G168), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT51), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1096), .A2(new_n1101), .A3(G8), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1059), .B2(G2078), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1056), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n1108));
  OAI221_X1 g683(.A(new_n1106), .B1(G1961), .B2(new_n1064), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G171), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1103), .A2(new_n1104), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1052), .B1(new_n1054), .B2(KEYINPUT50), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1348), .B1(new_n1112), .B2(new_n1061), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1036), .A2(G2067), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT121), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n707), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1114), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n620), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1075), .A2(new_n748), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(G2072), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1056), .A2(new_n1058), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n573), .B(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1120), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n573), .B(KEYINPUT57), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT122), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1129), .A2(new_n1134), .A3(new_n1131), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT123), .B(G1996), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1056), .A2(new_n1058), .A3(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT58), .B(G1341), .Z(new_n1140));
  NAND2_X1  g715(.A1(new_n1036), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n628), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1136), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1143), .B2(new_n1142), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1130), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OR3_X1    g724(.A1(new_n1142), .A2(new_n1143), .A3(KEYINPUT59), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1128), .A2(new_n1131), .A3(KEYINPUT61), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1145), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1117), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT60), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1115), .A2(new_n1156), .A3(new_n1119), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n620), .A3(new_n1157), .ZN(new_n1158));
  OAI221_X1 g733(.A(KEYINPUT60), .B1(new_n619), .B2(new_n617), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1133), .B(new_n1135), .C1(new_n1152), .C2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(G301), .B(KEYINPUT54), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1109), .A2(new_n1162), .ZN(new_n1163));
  AND4_X1   g738(.A1(KEYINPUT53), .A2(new_n1058), .A3(new_n750), .A4(new_n1035), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT45), .B1(new_n503), .B2(new_n1057), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1162), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1106), .B(new_n1167), .C1(G1961), .C2(new_n1064), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1169), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1111), .B1(new_n1161), .B2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1091), .B(new_n1095), .C1(new_n1171), .C2(new_n1087), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1165), .A2(new_n1035), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n735), .B(new_n741), .ZN(new_n1174));
  INV_X1    g749(.A(G1996), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n761), .B(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1173), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT114), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1173), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n829), .A2(new_n834), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n829), .A2(new_n834), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1179), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  XOR2_X1   g758(.A(G290), .B(G1986), .Z(new_n1184));
  OAI21_X1  g759(.A(new_n1183), .B1(new_n1173), .B2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT115), .Z(new_n1186));
  NAND2_X1  g761(.A1(new_n1172), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n735), .A2(G2067), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1189), .A2(KEYINPUT125), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1179), .ZN(new_n1192));
  AOI21_X1  g767(.A(KEYINPUT125), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1188), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1174), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1179), .B1(new_n1195), .B2(new_n761), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1179), .A2(KEYINPUT46), .A3(new_n1175), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT46), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1198), .B1(new_n1173), .B2(G1996), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1200));
  XOR2_X1   g775(.A(new_n1200), .B(KEYINPUT47), .Z(new_n1201));
  NOR3_X1   g776(.A1(new_n1173), .A2(G1986), .A3(G290), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT48), .Z(new_n1203));
  AOI21_X1  g778(.A(new_n1201), .B1(new_n1183), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1194), .A2(new_n1204), .ZN(new_n1205));
  NOR3_X1   g780(.A1(new_n1192), .A2(new_n1188), .A3(new_n1193), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1187), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g783(.A(G319), .B1(new_n667), .B2(new_n668), .ZN(new_n1210));
  NOR2_X1   g784(.A1(G227), .A2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g785(.A(new_n1211), .B1(new_n702), .B2(new_n703), .ZN(new_n1212));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n1213));
  XNOR2_X1  g787(.A(new_n1212), .B(new_n1213), .ZN(new_n1214));
  AOI21_X1  g788(.A(new_n1214), .B1(new_n906), .B2(new_n910), .ZN(new_n1215));
  NAND2_X1  g789(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1216));
  AND2_X1   g790(.A1(new_n1215), .A2(new_n1216), .ZN(G308));
  NAND2_X1  g791(.A1(new_n1215), .A2(new_n1216), .ZN(G225));
endmodule


