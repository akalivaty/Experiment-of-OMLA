//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n188));
  INV_X1    g002(.A(G113), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(KEYINPUT69), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT69), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n191), .B1(KEYINPUT2), .B2(G113), .ZN(new_n192));
  AOI22_X1  g006(.A1(new_n190), .A2(new_n192), .B1(KEYINPUT2), .B2(G113), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G116), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT70), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n195), .A2(new_n197), .A3(KEYINPUT70), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n200), .B1(new_n204), .B2(new_n193), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G137), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  OAI211_X1 g026(.A(KEYINPUT66), .B(new_n212), .C1(new_n209), .C2(G137), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(G134), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT66), .B1(new_n215), .B2(new_n212), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n211), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n211), .B(new_n219), .C1(new_n214), .C2(new_n216), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(KEYINPUT67), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n217), .A2(new_n222), .A3(G131), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G143), .ZN(new_n225));
  INV_X1    g039(.A(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT0), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT64), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT64), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n228), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G143), .B(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n236), .A2(KEYINPUT65), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n237), .B1(new_n228), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n235), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n221), .A2(new_n223), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT68), .B(G128), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(G143), .B2(new_n224), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n228), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n225), .A2(new_n227), .A3(new_n245), .A4(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n215), .A2(new_n210), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n249), .B(new_n220), .C1(new_n219), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n243), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT30), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT30), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n243), .A2(new_n254), .A3(new_n251), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n206), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n243), .A2(new_n206), .A3(new_n251), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT31), .B1(new_n256), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n252), .A2(new_n205), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(new_n257), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n243), .A2(new_n206), .A3(new_n251), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(KEYINPUT28), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n263), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n243), .A2(new_n254), .A3(new_n251), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n254), .B1(new_n243), .B2(new_n251), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n205), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n276));
  NAND4_X1  g090(.A1(new_n275), .A2(new_n257), .A3(new_n264), .A4(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n266), .A2(new_n272), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n279));
  NOR2_X1   g093(.A1(G472), .A2(G902), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n278), .B2(new_n280), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G472), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n206), .B1(new_n243), .B2(new_n251), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT28), .B1(new_n270), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n263), .B1(new_n257), .B2(new_n267), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(KEYINPUT29), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n263), .B1(new_n256), .B2(new_n270), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT29), .B1(new_n286), .B2(new_n287), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n290), .B1(new_n293), .B2(KEYINPUT73), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n291), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n284), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n187), .B1(new_n283), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n278), .A2(new_n280), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT32), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n293), .A2(KEYINPUT73), .ZN(new_n303));
  INV_X1    g117(.A(new_n290), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n296), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G472), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n302), .A2(new_n306), .A3(KEYINPUT74), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT22), .B(G137), .ZN(new_n308));
  INV_X1    g122(.A(G953), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(G221), .A3(G234), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n308), .B(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT77), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n316), .A3(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT78), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n313), .B2(G140), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT76), .A3(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n314), .A2(new_n316), .A3(new_n324), .A4(G140), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n318), .A2(KEYINPUT16), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT77), .B(G125), .ZN(new_n327));
  OR3_X1    g141(.A1(new_n327), .A2(KEYINPUT16), .A3(G140), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n326), .A2(G146), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(G146), .B1(new_n326), .B2(new_n328), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n244), .A2(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n194), .A2(G128), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT24), .B(G110), .Z(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n194), .B2(G128), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n333), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT75), .B1(new_n332), .B2(new_n336), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n244), .A2(new_n340), .A3(KEYINPUT23), .A4(G119), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n338), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G110), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n335), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n331), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n334), .B1(new_n332), .B2(new_n333), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n342), .B2(new_n343), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n326), .A2(G146), .A3(new_n328), .ZN(new_n348));
  XNOR2_X1  g162(.A(G125), .B(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n224), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n312), .B1(new_n345), .B2(new_n352), .ZN(new_n353));
  AOI211_X1 g167(.A(G110), .B(new_n338), .C1(new_n339), .C2(new_n341), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n350), .B(new_n348), .C1(new_n354), .C2(new_n346), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n355), .B(new_n311), .C1(new_n331), .C2(new_n344), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G234), .ZN(new_n358));
  AOI21_X1  g172(.A(G902), .B1(new_n358), .B2(G217), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  OR2_X1    g174(.A1(new_n360), .A2(KEYINPUT79), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n357), .A2(new_n362), .A3(new_n289), .ZN(new_n363));
  OAI21_X1  g177(.A(G217), .B1(new_n358), .B2(G902), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n353), .A2(new_n289), .A3(new_n356), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n360), .A2(KEYINPUT79), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n361), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n298), .A2(new_n307), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT80), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n298), .A2(new_n307), .A3(new_n373), .A4(new_n370), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G113), .B(G122), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT92), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT91), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n380), .A2(KEYINPUT19), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(KEYINPUT19), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n349), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n318), .A2(new_n323), .A3(new_n325), .ZN(new_n385));
  AOI211_X1 g199(.A(G146), .B(new_n384), .C1(new_n385), .C2(KEYINPUT19), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n379), .B1(new_n386), .B2(new_n329), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n259), .A2(G214), .ZN(new_n388));
  OR2_X1    g202(.A1(KEYINPUT89), .A2(G143), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT89), .A2(G143), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n388), .A2(new_n390), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n219), .ZN(new_n394));
  OAI21_X1  g208(.A(G131), .B1(new_n391), .B2(new_n392), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n325), .A2(new_n323), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n324), .B1(new_n327), .B2(G140), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT19), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n224), .A3(new_n383), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT92), .A3(new_n348), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n387), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n395), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT18), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n385), .A2(G146), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n350), .ZN(new_n406));
  NAND2_X1  g220(.A1(KEYINPUT18), .A2(G131), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n393), .A2(KEYINPUT90), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT90), .B1(new_n393), .B2(new_n407), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n404), .B(new_n406), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n378), .B1(new_n402), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n403), .A2(KEYINPUT17), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n394), .A2(new_n413), .A3(new_n395), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n331), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n415), .A2(new_n378), .A3(new_n410), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT93), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(G475), .A2(G902), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n401), .A2(new_n396), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT92), .B1(new_n400), .B2(new_n348), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n410), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n378), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n415), .A2(new_n378), .A3(new_n410), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n417), .A2(new_n418), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n423), .A2(new_n425), .ZN(new_n428));
  NOR3_X1   g242(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n427), .A2(KEYINPUT20), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n378), .B1(new_n415), .B2(new_n410), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n416), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n289), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n433), .A2(G475), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n196), .A2(G122), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n435), .B(KEYINPUT94), .Z(new_n436));
  NAND2_X1  g250(.A1(new_n196), .A2(G122), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G107), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n436), .A2(G107), .A3(new_n437), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n436), .A2(KEYINPUT14), .A3(G107), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT95), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n244), .A2(G143), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n226), .A2(G128), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G134), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n447), .A2(G134), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n444), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n450), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT95), .A3(new_n448), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n436), .A2(KEYINPUT14), .A3(G107), .A4(new_n437), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n443), .A2(new_n451), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n447), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT13), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n209), .B1(new_n445), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n456), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n440), .A3(new_n441), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT9), .B(G234), .ZN(new_n461));
  INV_X1    g275(.A(G217), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n461), .A2(new_n462), .A3(G953), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n455), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n463), .B1(new_n455), .B2(new_n460), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n289), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G478), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(KEYINPUT15), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI221_X1 g283(.A(new_n289), .B1(KEYINPUT15), .B2(new_n467), .C1(new_n464), .C2(new_n465), .ZN(new_n470));
  NAND2_X1  g284(.A1(G234), .A2(G237), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n471), .A2(G952), .A3(new_n309), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(G902), .A3(G953), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT96), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(G898), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n469), .A2(new_n470), .A3(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n430), .A2(new_n434), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G214), .B1(G237), .B2(G902), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n309), .A2(G224), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT7), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n247), .A2(new_n327), .A3(new_n248), .ZN(new_n485));
  INV_X1    g299(.A(new_n327), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n486), .B(new_n235), .C1(new_n239), .C2(new_n241), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n485), .B1(new_n487), .B2(KEYINPUT87), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n238), .B1(new_n236), .B2(KEYINPUT65), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n228), .A2(new_n240), .A3(new_n237), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n225), .A2(new_n227), .B1(new_n231), .B2(new_n232), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n490), .A2(new_n491), .B1(new_n492), .B2(new_n234), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n489), .B1(new_n493), .B2(new_n486), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n484), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n195), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT5), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n189), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n203), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT70), .B1(new_n195), .B2(new_n197), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n498), .B1(new_n501), .B2(new_n497), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n377), .A2(G107), .ZN(new_n503));
  AND2_X1   g317(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n504));
  NOR2_X1   g318(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G101), .ZN(new_n507));
  OR2_X1    g321(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n439), .A2(G104), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n377), .A2(G107), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n506), .A2(new_n507), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n511), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G101), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n502), .A2(new_n515), .A3(new_n200), .ZN(new_n516));
  NAND2_X1  g330(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n509), .B1(new_n508), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n511), .B1(new_n503), .B2(new_n505), .ZN(new_n519));
  OAI21_X1  g333(.A(G101), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT4), .A3(new_n512), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT4), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n522), .B(G101), .C1(new_n518), .C2(new_n519), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n205), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(G110), .B(G122), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n516), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n512), .A2(new_n514), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n502), .A2(new_n527), .A3(new_n200), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n498), .B1(new_n497), .B2(new_n198), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n200), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n515), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n525), .B(KEYINPUT8), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n487), .A2(KEYINPUT87), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n493), .A2(new_n489), .A3(new_n486), .ZN(new_n535));
  INV_X1    g349(.A(new_n484), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n485), .A4(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n495), .A2(new_n526), .A3(new_n533), .A4(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n538), .A2(new_n289), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n516), .A2(new_n524), .ZN(new_n540));
  INV_X1    g354(.A(new_n525), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(KEYINPUT6), .A3(new_n526), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT6), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n540), .A2(new_n544), .A3(new_n541), .ZN(new_n545));
  OAI211_X1 g359(.A(G224), .B(new_n309), .C1(new_n488), .C2(new_n494), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n534), .A2(new_n535), .A3(new_n483), .A4(new_n485), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n543), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n539), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G210), .B1(G237), .B2(G902), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n552), .B(KEYINPUT88), .Z(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n539), .A2(new_n549), .A3(new_n552), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n482), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT86), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT12), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n248), .A2(KEYINPUT84), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT84), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n236), .A2(new_n560), .A3(new_n245), .A4(G128), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n228), .B1(new_n246), .B2(new_n230), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n512), .A3(new_n514), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n247), .A2(new_n248), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n527), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n221), .A2(new_n223), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n558), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(new_n566), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n570), .A2(KEYINPUT12), .A3(new_n223), .A4(new_n221), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT85), .ZN(new_n573));
  XNOR2_X1  g387(.A(G110), .B(G140), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n309), .A2(G227), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n521), .A2(new_n242), .A3(new_n523), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n578), .B1(new_n579), .B2(new_n527), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n515), .A2(KEYINPUT10), .A3(new_n249), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n577), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n576), .B1(new_n582), .B2(new_n568), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT85), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n569), .A2(new_n584), .A3(new_n571), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n573), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n577), .A2(new_n580), .A3(new_n581), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n223), .A3(new_n221), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n568), .A2(new_n577), .A3(new_n580), .A4(new_n581), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n576), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G469), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n289), .ZN(new_n594));
  INV_X1    g408(.A(new_n576), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n588), .A2(new_n589), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n569), .A2(new_n571), .B1(new_n582), .B2(new_n568), .ZN(new_n597));
  OAI211_X1 g411(.A(G469), .B(new_n596), .C1(new_n597), .C2(new_n595), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n593), .A2(new_n289), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(G221), .B1(new_n461), .B2(G902), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n604), .B(KEYINPUT81), .Z(new_n605));
  XOR2_X1   g419(.A(new_n605), .B(KEYINPUT82), .Z(new_n606));
  AOI21_X1  g420(.A(new_n557), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(G902), .B1(new_n586), .B2(new_n591), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n601), .B1(new_n608), .B2(new_n593), .ZN(new_n609));
  INV_X1    g423(.A(new_n606), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n609), .A2(KEYINPUT86), .A3(new_n610), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n480), .B(new_n556), .C1(new_n607), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT97), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n603), .A2(new_n557), .A3(new_n606), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT86), .B1(new_n609), .B2(new_n610), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n480), .A4(new_n556), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n375), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT98), .B(G101), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G3));
  INV_X1    g436(.A(new_n299), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n284), .B1(new_n278), .B2(new_n289), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n369), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n626), .A2(new_n616), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n427), .A2(KEYINPUT20), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n428), .A2(new_n429), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n433), .A2(G475), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n466), .A2(new_n467), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n464), .A2(new_n465), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT100), .B(KEYINPUT33), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(KEYINPUT100), .A2(KEYINPUT33), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n636), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n289), .A2(G478), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n633), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n539), .A2(new_n549), .A3(new_n552), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n552), .B1(new_n539), .B2(new_n549), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n481), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT99), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n648), .B(new_n481), .C1(new_n644), .C2(new_n645), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n647), .A2(new_n478), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n627), .A2(new_n643), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT34), .B(G104), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  NAND2_X1  g467(.A1(new_n469), .A2(new_n470), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT20), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n417), .A2(new_n426), .A3(new_n655), .A4(new_n418), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n434), .B1(new_n628), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n650), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n627), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  OAI22_X1  g476(.A1(new_n345), .A2(new_n352), .B1(KEYINPUT36), .B2(new_n312), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n312), .A2(KEYINPUT36), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n355), .B(new_n664), .C1(new_n331), .C2(new_n344), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n663), .A2(new_n359), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n363), .B2(new_n366), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n625), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n613), .A2(new_n618), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT37), .B(G110), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G12));
  NOR3_X1   g485(.A1(new_n283), .A2(new_n297), .A3(new_n187), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT74), .B1(new_n302), .B2(new_n306), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n628), .A2(new_n656), .ZN(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n472), .B1(new_n475), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n675), .A2(new_n631), .A3(new_n654), .A4(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n667), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n647), .A2(new_n649), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n674), .A2(new_n681), .A3(new_n616), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XOR2_X1   g500(.A(new_n677), .B(KEYINPUT39), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n616), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n554), .A2(new_n555), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT38), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT38), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n554), .A2(new_n693), .A3(new_n555), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n481), .A3(new_n667), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n256), .A2(new_n265), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n264), .B1(new_n268), .B2(new_n257), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n289), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G472), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n302), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n632), .A2(new_n654), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n689), .A2(new_n690), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  OAI211_X1 g520(.A(new_n641), .B(new_n678), .C1(new_n430), .C2(new_n434), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n674), .A2(new_n616), .A3(new_n684), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  NAND2_X1  g524(.A1(KEYINPUT102), .A2(G469), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n608), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n608), .A2(new_n711), .ZN(new_n713));
  INV_X1    g527(.A(new_n605), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n298), .A2(new_n307), .A3(new_n370), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n643), .A2(new_n650), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT41), .B(G113), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  AND3_X1   g535(.A1(new_n298), .A2(new_n307), .A3(new_n370), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(KEYINPUT103), .A3(new_n659), .A4(new_n716), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n724), .B1(new_n717), .B2(new_n658), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NOR2_X1   g541(.A1(new_n683), .A2(new_n715), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n298), .A2(new_n728), .A3(new_n307), .A4(new_n480), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  NOR2_X1   g544(.A1(new_n715), .A2(new_n477), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n647), .A2(new_n649), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n280), .B(KEYINPUT104), .Z(new_n733));
  AND2_X1   g547(.A1(new_n278), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n369), .A2(new_n734), .A3(new_n624), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n704), .A2(new_n731), .A3(new_n732), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  NOR3_X1   g551(.A1(new_n734), .A2(new_n624), .A3(new_n667), .ZN(new_n738));
  AND4_X1   g552(.A1(new_n732), .A2(new_n708), .A3(new_n716), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n313), .ZN(G27));
  OAI21_X1  g554(.A(KEYINPUT105), .B1(new_n609), .B2(new_n605), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  AOI211_X1 g556(.A(G469), .B(G902), .C1(new_n586), .C2(new_n591), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n742), .B(new_n714), .C1(new_n743), .C2(new_n601), .ZN(new_n744));
  INV_X1    g558(.A(new_n553), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n481), .B(new_n555), .C1(new_n550), .C2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n741), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n298), .A3(new_n307), .A4(new_n370), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n707), .A2(KEYINPUT42), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n369), .B1(new_n302), .B2(new_n306), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n748), .A2(new_n708), .A3(new_n752), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n750), .A2(new_n751), .B1(KEYINPUT42), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  XNOR2_X1  g569(.A(new_n679), .B(KEYINPUT101), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n749), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n209), .ZN(G36));
  NOR2_X1   g572(.A1(new_n430), .A2(new_n434), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n641), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n762), .B1(new_n632), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n761), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n625), .A2(new_n682), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT107), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n765), .A2(new_n767), .A3(KEYINPUT44), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n747), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n596), .B1(new_n597), .B2(new_n595), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n593), .B1(new_n775), .B2(new_n776), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n600), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(KEYINPUT46), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n594), .B1(new_n781), .B2(KEYINPUT46), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n605), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n770), .A2(KEYINPUT108), .A3(new_n747), .A4(new_n771), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n774), .A2(new_n687), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(KEYINPUT47), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(KEYINPUT47), .ZN(new_n791));
  OAI221_X1 g605(.A(new_n714), .B1(new_n790), .B2(new_n791), .C1(new_n783), .C2(new_n782), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n785), .B2(new_n791), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n369), .A2(new_n747), .ZN(new_n794));
  OR4_X1    g608(.A1(new_n674), .A2(new_n793), .A3(new_n707), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n626), .A2(new_n478), .A3(new_n616), .A4(new_n556), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n759), .A2(new_n654), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n669), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n642), .B(KEYINPUT111), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n798), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n620), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n801), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n739), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n682), .A2(new_n609), .A3(new_n605), .A4(new_n677), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n704), .A2(new_n809), .A3(new_n732), .A4(new_n701), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n685), .A2(new_n709), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n616), .A2(new_n298), .A3(new_n307), .A4(new_n684), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n739), .B1(new_n814), .B2(new_n681), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT52), .A3(new_n709), .A4(new_n810), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n803), .B1(new_n375), .B2(new_n619), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT112), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n469), .A2(new_n470), .A3(new_n678), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n746), .A2(new_n667), .A3(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(new_n657), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n298), .A3(new_n616), .A4(new_n307), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n748), .A2(new_n708), .A3(new_n738), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n757), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n729), .A2(new_n736), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n719), .A2(new_n827), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n726), .A2(new_n826), .A3(new_n754), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n807), .A2(new_n817), .A3(new_n819), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n797), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n815), .A2(new_n812), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n831), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n801), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n818), .B2(KEYINPUT112), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n620), .A2(KEYINPUT112), .A3(new_n804), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n726), .A2(new_n826), .A3(new_n754), .A4(new_n828), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(KEYINPUT113), .A3(KEYINPUT53), .A4(new_n817), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n832), .A2(new_n834), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT54), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT53), .B1(new_n830), .B2(new_n833), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n839), .A2(new_n831), .A3(new_n817), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n712), .A2(new_n713), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n793), .B1(new_n606), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n765), .A2(new_n472), .A3(new_n735), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n747), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n764), .B(new_n760), .ZN(new_n852));
  INV_X1    g666(.A(new_n472), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n715), .A2(new_n746), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n738), .A3(new_n855), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n472), .A2(new_n702), .A3(new_n370), .A4(new_n855), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n632), .A2(new_n641), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n692), .A2(new_n482), .A3(new_n694), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n715), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT114), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n854), .A2(new_n863), .A3(new_n735), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT50), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n850), .A2(KEYINPUT50), .A3(new_n863), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n860), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(KEYINPUT51), .B(new_n851), .C1(new_n868), .C2(KEYINPUT115), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n868), .A2(KEYINPUT115), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n867), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n856), .A3(new_n851), .A4(new_n859), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n850), .A2(new_n732), .A3(new_n716), .ZN(new_n876));
  INV_X1    g690(.A(G952), .ZN(new_n877));
  AOI211_X1 g691(.A(new_n877), .B(G953), .C1(new_n857), .C2(new_n643), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n854), .A2(new_n752), .A3(new_n855), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n880), .A2(KEYINPUT48), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(KEYINPUT48), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n875), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n871), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n842), .A2(new_n847), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT116), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n842), .A2(new_n885), .A3(new_n888), .A4(new_n847), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n877), .A2(new_n309), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n370), .A2(new_n606), .A3(new_n481), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n695), .B(new_n892), .C1(KEYINPUT49), .C2(new_n848), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n848), .A2(KEYINPUT49), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT110), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n893), .A2(new_n702), .A3(new_n761), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n891), .A2(KEYINPUT117), .A3(new_n896), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(G75));
  NOR2_X1   g715(.A1(new_n309), .A2(G952), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n543), .A2(new_n545), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n548), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n845), .A2(new_n289), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(G210), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n906), .A2(new_n553), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n905), .A2(new_n908), .ZN(new_n911));
  AOI211_X1 g725(.A(new_n902), .B(new_n909), .C1(new_n910), .C2(new_n911), .ZN(G51));
  XNOR2_X1  g726(.A(new_n845), .B(KEYINPUT54), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n599), .B(KEYINPUT57), .Z(new_n914));
  OAI21_X1  g728(.A(new_n592), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n906), .A2(new_n777), .A3(new_n778), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n902), .B1(new_n915), .B2(new_n916), .ZN(G54));
  NAND3_X1  g731(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n417), .A2(new_n426), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT118), .ZN(new_n921));
  INV_X1    g735(.A(new_n902), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n918), .A2(new_n923), .A3(new_n919), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n918), .B2(new_n919), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n921), .A2(new_n926), .ZN(G60));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  NOR3_X1   g743(.A1(new_n913), .A2(new_n639), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n842), .A2(new_n847), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n931), .A2(new_n929), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n902), .B(new_n930), .C1(new_n932), .C2(new_n639), .ZN(G63));
  XNOR2_X1  g747(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n462), .A2(new_n289), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n843), .A2(new_n844), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n665), .A3(new_n663), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n938), .B(new_n922), .C1(new_n357), .C2(new_n937), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT61), .Z(G66));
  INV_X1    g754(.A(G224), .ZN(new_n941));
  OAI21_X1  g755(.A(G953), .B1(new_n476), .B2(new_n941), .ZN(new_n942));
  AND4_X1   g756(.A1(new_n726), .A2(new_n807), .A3(new_n819), .A4(new_n828), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(G953), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n903), .B1(G898), .B2(new_n309), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT121), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n944), .B(new_n946), .ZN(G69));
  INV_X1    g761(.A(new_n757), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n704), .A2(new_n732), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n785), .A2(new_n687), .A3(new_n950), .A4(new_n752), .ZN(new_n951));
  AND4_X1   g765(.A1(new_n754), .A2(new_n795), .A3(new_n948), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n815), .A2(new_n709), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT123), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n952), .A2(new_n787), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n309), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n253), .A2(new_n255), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n399), .A2(new_n383), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT122), .Z(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n956), .B(new_n960), .C1(new_n676), .C2(new_n309), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n954), .A2(new_n705), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n963), .A2(KEYINPUT124), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(KEYINPUT124), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI211_X1 g780(.A(new_n688), .B(new_n746), .C1(new_n802), .C2(new_n799), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n375), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n787), .A2(new_n795), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(KEYINPUT62), .B2(new_n962), .ZN(new_n970));
  AOI21_X1  g784(.A(G953), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n961), .B1(new_n971), .B2(new_n960), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n309), .B1(G227), .B2(G900), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(G72));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n955), .B2(new_n943), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n275), .A2(new_n257), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT125), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n263), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n922), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n291), .B1(new_n256), .B2(new_n265), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n976), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT127), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n983), .B1(new_n841), .B2(new_n986), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n970), .B(new_n943), .C1(new_n964), .C2(new_n965), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n976), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT126), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n981), .A2(new_n263), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n990), .B1(new_n989), .B2(new_n991), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(G57));
endmodule


