//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT65), .Z(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n463), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  NAND4_X1  g057(.A1(new_n471), .A2(new_n473), .A3(G126), .A4(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n471), .A2(new_n473), .A3(G138), .A4(new_n463), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n462), .A2(new_n490), .A3(G138), .A4(new_n463), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n487), .B1(new_n489), .B2(new_n491), .ZN(G164));
  INV_X1    g067(.A(G543), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT5), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G543), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT6), .B(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G88), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G50), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n497), .A2(G62), .ZN(new_n505));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  XOR2_X1   g081(.A(new_n506), .B(KEYINPUT66), .Z(new_n507));
  AOI21_X1  g082(.A(new_n504), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n503), .A2(new_n508), .ZN(G303));
  INV_X1    g084(.A(G303), .ZN(G166));
  NAND3_X1  g085(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT7), .ZN(new_n512));
  INV_X1    g087(.A(G51), .ZN(new_n513));
  INV_X1    g088(.A(G89), .ZN(new_n514));
  OAI221_X1 g089(.A(new_n512), .B1(new_n501), .B2(new_n513), .C1(new_n499), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n494), .A2(new_n496), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT67), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n494), .A2(new_n496), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n515), .A2(new_n521), .ZN(G168));
  AND2_X1   g097(.A1(new_n497), .A2(new_n498), .ZN(new_n523));
  INV_X1    g098(.A(new_n501), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT69), .B(G52), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n523), .A2(G90), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n494), .A2(new_n496), .A3(new_n518), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n518), .B1(new_n494), .B2(new_n496), .ZN(new_n528));
  OAI21_X1  g103(.A(G64), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n530), .B1(new_n529), .B2(new_n531), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n526), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n529), .A2(new_n531), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT68), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n539), .A2(G651), .A3(new_n532), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT70), .B1(new_n540), .B2(new_n526), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n523), .A2(G81), .B1(new_n524), .B2(G43), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n545), .B2(new_n504), .ZN(new_n546));
  INV_X1    g121(.A(G860), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n546), .A2(new_n547), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  NAND3_X1  g128(.A1(new_n498), .A2(G53), .A3(G543), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT9), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n497), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n504), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n499), .B(KEYINPUT71), .ZN(new_n558));
  INV_X1    g133(.A(G91), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n555), .B(new_n557), .C1(new_n558), .C2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G168), .ZN(G286));
  OR2_X1    g136(.A1(new_n520), .A2(G74), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(G49), .B2(new_n524), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n499), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G288));
  AOI22_X1  g142(.A1(new_n565), .A2(G86), .B1(G48), .B2(new_n524), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n497), .A2(G61), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n569), .A2(new_n570), .B1(G73), .B2(G543), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n497), .A2(KEYINPUT72), .A3(G61), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n504), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n568), .A2(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n523), .A2(G85), .B1(new_n524), .B2(G47), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n520), .A2(G60), .ZN(new_n577));
  INV_X1    g152(.A(G72), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n493), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT73), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n579), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n576), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT74), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT74), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n585), .B(new_n576), .C1(new_n581), .C2(new_n582), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n524), .A2(KEYINPUT75), .ZN(new_n589));
  INV_X1    g164(.A(G54), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n590), .B1(new_n501), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT76), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n516), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n589), .A2(new_n592), .B1(new_n596), .B2(G651), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n565), .A2(KEYINPUT10), .A3(G92), .ZN(new_n598));
  AOI21_X1  g173(.A(KEYINPUT10), .B1(new_n565), .B2(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT77), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n588), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n588), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(G168), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(new_n605), .B2(G168), .ZN(G280));
  NOR2_X1   g183(.A1(new_n601), .A2(G559), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(G860), .B2(new_n602), .ZN(G148));
  NAND2_X1  g185(.A1(new_n546), .A2(new_n605), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n609), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n462), .A2(new_n460), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT12), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(G2100), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n475), .A2(G123), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n477), .A2(G135), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n463), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2096), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n616), .A2(G2100), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n617), .A2(new_n623), .A3(new_n624), .ZN(G156));
  INV_X1    g200(.A(G14), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2435), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(KEYINPUT14), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n626), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(KEYINPUT17), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n644), .A2(new_n645), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n649), .B(new_n651), .C1(new_n652), .C2(new_n648), .ZN(new_n653));
  OR3_X1    g228(.A1(new_n651), .A2(KEYINPUT18), .A3(new_n647), .ZN(new_n654));
  OAI21_X1  g229(.A(KEYINPUT18), .B1(new_n651), .B2(new_n647), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2096), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT20), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n662), .B2(new_n663), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n666), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT80), .Z(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n673), .B(new_n679), .ZN(G229));
  MUX2_X1   g255(.A(G6), .B(G305), .S(G16), .Z(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT32), .B(G1981), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n684), .A2(G23), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(G288), .B2(G16), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT33), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n681), .A2(new_n682), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n684), .A2(G22), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G166), .B2(new_n684), .ZN(new_n692));
  INV_X1    g267(.A(G1971), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n686), .A2(new_n689), .ZN(new_n695));
  NAND4_X1  g270(.A1(new_n683), .A2(new_n690), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT34), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G25), .A2(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n475), .A2(G119), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n477), .A2(G131), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n463), .A2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT81), .Z(new_n705));
  AOI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(G29), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XOR2_X1   g282(.A(new_n706), .B(new_n707), .Z(new_n708));
  INV_X1    g283(.A(G1986), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n684), .A2(G24), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G290), .B2(G16), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n708), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n698), .B(new_n712), .C1(new_n709), .C2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(G168), .A2(G16), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT88), .Z(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G16), .B2(G21), .ZN(new_n718));
  INV_X1    g293(.A(G1966), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT31), .B(G11), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT89), .B(KEYINPUT30), .Z(new_n722));
  AOI21_X1  g297(.A(G29), .B1(new_n722), .B2(G28), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G28), .B2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n721), .B(new_n724), .C1(new_n622), .C2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G1961), .ZN(new_n728));
  NOR2_X1   g303(.A1(G171), .A2(new_n684), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G5), .B2(new_n684), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n727), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n725), .A2(G35), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G162), .B2(new_n725), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT29), .Z(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(G2090), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT91), .ZN(new_n740));
  INV_X1    g315(.A(G299), .ZN(new_n741));
  OAI21_X1  g316(.A(KEYINPUT23), .B1(new_n741), .B2(new_n684), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n684), .A2(G20), .ZN(new_n743));
  MUX2_X1   g318(.A(KEYINPUT23), .B(new_n742), .S(new_n743), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G1956), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(G1956), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n740), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT28), .ZN(new_n748));
  INV_X1    g323(.A(G26), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G29), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(G29), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n475), .A2(KEYINPUT84), .A3(G128), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT84), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n462), .A2(G2105), .ZN(new_n754));
  INV_X1    g329(.A(G128), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n477), .A2(G140), .ZN(new_n757));
  OR2_X1    g332(.A1(G104), .A2(G2105), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n758), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n752), .A2(new_n756), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n751), .B1(new_n760), .B2(G29), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n750), .B1(new_n761), .B2(new_n748), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(G2067), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(G2067), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n725), .A2(G32), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n477), .A2(G141), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT85), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n460), .A2(G105), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT26), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n769), .B(new_n771), .C1(G129), .C2(new_n475), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT86), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n765), .B1(new_n774), .B2(new_n725), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT87), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n763), .B(new_n764), .C1(new_n775), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G29), .A2(G33), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n460), .A2(G103), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT25), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G139), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n782), .B1(new_n464), .B2(new_n783), .C1(new_n784), .C2(new_n463), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(G29), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(G2072), .Z(new_n788));
  INV_X1    g363(.A(KEYINPUT24), .ZN(new_n789));
  INV_X1    g364(.A(G34), .ZN(new_n790));
  AOI21_X1  g365(.A(G29), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G160), .B2(new_n725), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G2084), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n725), .A2(G27), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G164), .B2(new_n725), .ZN(new_n796));
  INV_X1    g371(.A(G2078), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n788), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n775), .B2(new_n777), .ZN(new_n800));
  MUX2_X1   g375(.A(G19), .B(new_n546), .S(G16), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1341), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G2090), .B2(new_n738), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n747), .A2(new_n778), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G4), .A2(G16), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n602), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1348), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n728), .B2(new_n730), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n733), .A2(new_n734), .A3(new_n805), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n715), .A2(new_n810), .ZN(G311));
  XNOR2_X1  g386(.A(new_n713), .B(KEYINPUT36), .ZN(new_n812));
  AND3_X1   g387(.A1(new_n734), .A2(new_n805), .A3(new_n809), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n812), .A2(new_n733), .A3(new_n813), .ZN(G150));
  NAND2_X1  g389(.A1(new_n602), .A2(G559), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT92), .B(KEYINPUT38), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT39), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT94), .B(G55), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n523), .A2(G93), .B1(new_n524), .B2(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT93), .B1(new_n821), .B2(new_n504), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n821), .A2(KEYINPUT93), .A3(new_n504), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n825), .A2(KEYINPUT95), .A3(new_n546), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n546), .A2(KEYINPUT95), .ZN(new_n827));
  OR3_X1    g402(.A1(new_n821), .A2(KEYINPUT93), .A3(new_n504), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(new_n822), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n546), .A2(KEYINPUT95), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n827), .A2(new_n829), .A3(new_n830), .A4(new_n820), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n818), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n818), .A2(new_n832), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n833), .A2(new_n547), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n825), .A2(G860), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT97), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT96), .B(KEYINPUT37), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n835), .A2(new_n839), .ZN(G145));
  XOR2_X1   g415(.A(new_n622), .B(G160), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n481), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n475), .A2(new_n843), .A3(G130), .ZN(new_n844));
  INV_X1    g419(.A(G130), .ZN(new_n845));
  OAI21_X1  g420(.A(KEYINPUT98), .B1(new_n754), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n477), .A2(G142), .ZN(new_n847));
  OR2_X1    g422(.A1(G106), .A2(G2105), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n844), .A2(new_n846), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n704), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT99), .ZN(new_n852));
  INV_X1    g427(.A(new_n615), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n774), .A2(new_n786), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n773), .A2(new_n785), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n760), .B(G164), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n860), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n857), .A2(new_n862), .A3(new_n858), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n856), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n854), .A2(new_n861), .A3(new_n855), .A4(new_n863), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n842), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n870), .A2(new_n866), .A3(new_n865), .ZN(new_n871));
  AOI21_X1  g446(.A(G37), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(KEYINPUT101), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n865), .A2(KEYINPUT100), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n856), .A2(new_n864), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n868), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n873), .A2(new_n874), .A3(new_n876), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n842), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT40), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n872), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(G395));
  XNOR2_X1  g460(.A(new_n609), .B(new_n832), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n600), .A2(new_n741), .ZN(new_n887));
  OAI211_X1 g462(.A(G299), .B(new_n597), .C1(new_n598), .C2(new_n599), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(KEYINPUT103), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n600), .A2(new_n741), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n888), .ZN(new_n894));
  XNOR2_X1  g469(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n893), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n886), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n826), .A2(new_n831), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n609), .B(new_n899), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n898), .A2(KEYINPUT105), .B1(new_n900), .B2(new_n894), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n886), .A2(new_n902), .A3(new_n897), .ZN(new_n903));
  NAND2_X1  g478(.A1(G290), .A2(G166), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n584), .A2(G303), .A3(new_n586), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(G305), .B(G288), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT42), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n901), .A2(new_n903), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n901), .B2(new_n903), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n825), .A2(new_n605), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(G295));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n916), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n537), .B2(new_n541), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n535), .A2(new_n536), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n540), .A2(KEYINPUT70), .A3(new_n526), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(KEYINPUT106), .A3(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n921), .A2(G286), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G286), .B1(new_n921), .B2(new_n924), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n925), .A2(new_n926), .A3(new_n832), .ZN(new_n927));
  INV_X1    g502(.A(new_n924), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT106), .B1(new_n922), .B2(new_n923), .ZN(new_n929));
  OAI21_X1  g504(.A(G168), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n921), .A2(G286), .A3(new_n924), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n899), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n894), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n832), .B1(new_n925), .B2(new_n926), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(new_n899), .A3(new_n931), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n897), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n911), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G37), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n911), .B1(new_n933), .B2(new_n936), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n919), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n890), .B1(new_n889), .B2(new_n892), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n934), .A2(new_n935), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n894), .A2(new_n896), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n933), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n911), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n947), .A2(KEYINPUT43), .A3(new_n938), .A4(new_n937), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT44), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n939), .B2(new_n940), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n947), .A2(new_n919), .A3(new_n938), .A4(new_n937), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n950), .A2(new_n955), .ZN(G397));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G164), .B2(G1384), .ZN(new_n958));
  INV_X1    g533(.A(G125), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n468), .B1(new_n474), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(G2105), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n477), .A2(G137), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n961), .A2(new_n962), .A3(G40), .A4(new_n461), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(G1996), .A3(new_n773), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(KEYINPUT108), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(KEYINPUT108), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n760), .A2(G2067), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n760), .A2(G2067), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1996), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n964), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT107), .Z(new_n974));
  AOI211_X1 g549(.A(new_n966), .B(new_n971), .C1(new_n974), .C2(new_n774), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n975), .A2(new_n707), .A3(new_n705), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n964), .B1(new_n976), .B2(new_n969), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n974), .A2(KEYINPUT46), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n964), .A2(new_n773), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n970), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n980), .B(KEYINPUT125), .Z(new_n981));
  NAND2_X1  g556(.A1(new_n974), .A2(KEYINPUT46), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n978), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT47), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n977), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n964), .ZN(new_n986));
  NOR3_X1   g561(.A1(G290), .A2(G1986), .A3(new_n986), .ZN(new_n987));
  XOR2_X1   g562(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n988));
  XNOR2_X1  g563(.A(new_n987), .B(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n704), .B(new_n707), .Z(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n964), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n975), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n989), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n985), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(G288), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT52), .B1(G288), .B2(new_n998), .ZN(new_n1000));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n466), .A2(new_n469), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n489), .A2(new_n491), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n483), .A2(new_n486), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n563), .A2(new_n566), .A3(KEYINPUT112), .A4(G1976), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n999), .A2(new_n1000), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n999), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1981), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n568), .A2(new_n1015), .A3(new_n574), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n523), .A2(G86), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n524), .A2(G48), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1020), .A2(new_n573), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1016), .B1(new_n1022), .B2(new_n1015), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1016), .B(KEYINPUT49), .C1(new_n1022), .C2(new_n1015), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n1009), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1025), .A2(KEYINPUT114), .A3(new_n1026), .A4(new_n1009), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1014), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G303), .A2(G8), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT55), .ZN(new_n1033));
  AOI211_X1 g608(.A(new_n957), .B(G1384), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n958), .B1(new_n1034), .B2(KEYINPUT110), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1036));
  INV_X1    g611(.A(G1384), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT110), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n957), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1035), .A2(new_n1040), .A3(new_n1002), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1041), .A2(new_n693), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1043));
  NOR3_X1   g618(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1002), .B(new_n1043), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT111), .B(G2090), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1005), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(KEYINPUT116), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1042), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1033), .B1(new_n1052), .B2(new_n1008), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1043), .A2(new_n1002), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(new_n1044), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(new_n1047), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n1042), .B2(new_n1057), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1058), .A2(new_n1033), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1005), .A2(KEYINPUT45), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1005), .A2(KEYINPUT117), .A3(KEYINPUT45), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1062), .A2(new_n958), .A3(new_n1002), .A4(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT118), .B(G2084), .Z(new_n1065));
  AOI22_X1  g640(.A1(new_n1064), .A2(new_n719), .B1(new_n1055), .B2(new_n1065), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1066), .A2(new_n1008), .A3(G286), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1031), .A2(new_n1053), .A3(new_n1059), .A4(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1058), .A2(new_n1033), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1067), .A2(KEYINPUT63), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1031), .A2(new_n1059), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1016), .B(KEYINPUT115), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n563), .A2(new_n998), .A3(new_n566), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1059), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1078), .A2(new_n1009), .B1(new_n1079), .B2(new_n1031), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1064), .A2(new_n719), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1055), .A2(new_n1065), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1082), .B(G8), .C1(new_n1085), .C2(G286), .ZN(new_n1086));
  NOR2_X1   g661(.A1(G168), .A2(new_n1008), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT51), .B(new_n1088), .C1(new_n1066), .C2(new_n1008), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT124), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n958), .A2(KEYINPUT53), .A3(new_n797), .A4(new_n1002), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NOR4_X1   g671(.A1(G164), .A2(new_n1061), .A3(new_n957), .A4(G1384), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT117), .B1(new_n1005), .B2(KEYINPUT45), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(G1961), .B2(new_n1055), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1035), .A2(new_n797), .A3(new_n1040), .A4(new_n1002), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(KEYINPUT123), .A3(new_n1103), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1101), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1094), .B1(new_n1108), .B2(G301), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1102), .A2(KEYINPUT123), .A3(new_n1103), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT123), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(KEYINPUT124), .B(G171), .C1(new_n1112), .C2(new_n1101), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1093), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n963), .B1(new_n1038), .B2(KEYINPUT50), .ZN(new_n1117));
  AOI21_X1  g692(.A(G1348), .B1(new_n1117), .B2(new_n1049), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1006), .A2(G2067), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1116), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1348), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1054), .B2(new_n1044), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1006), .A2(G2067), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(KEYINPUT120), .A3(new_n1123), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n600), .ZN(new_n1126));
  INV_X1    g701(.A(G1956), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n1129));
  NAND2_X1  g704(.A1(G299), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n565), .A2(G91), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1131), .A2(new_n555), .A3(KEYINPUT57), .A4(new_n557), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT56), .B(G2072), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1035), .A2(new_n1040), .A3(new_n1002), .A4(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1128), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1125), .A2(new_n1126), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1128), .A2(new_n1135), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1133), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1035), .A2(new_n972), .A3(new_n1040), .A4(new_n1002), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT58), .B(G1341), .Z(new_n1143));
  NAND2_X1  g718(.A1(new_n1006), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n546), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1146), .ZN(new_n1148));
  AOI211_X1 g723(.A(new_n546), .B(new_n1148), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1128), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1133), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1140), .A2(KEYINPUT61), .A3(new_n1136), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1150), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1120), .A2(new_n1157), .A3(new_n1124), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1158), .A2(new_n1159), .A3(new_n1126), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n1158), .B2(new_n1126), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1125), .A2(new_n1157), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1156), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1160), .A2(new_n1161), .B1(new_n1157), .B2(new_n1125), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1141), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1056), .A2(new_n728), .B1(new_n1060), .B2(new_n1096), .ZN(new_n1167));
  OAI211_X1 g742(.A(G301), .B(new_n1167), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1109), .A2(new_n1113), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT54), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1086), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1167), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(G171), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1170), .B1(new_n1108), .B2(G301), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1172), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1115), .B1(new_n1166), .B2(new_n1177), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1031), .A2(new_n1053), .A3(new_n1059), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1081), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(G290), .B(new_n709), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n975), .B(new_n991), .C1(new_n1181), .C2(new_n986), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT109), .Z(new_n1183));
  OAI21_X1  g758(.A(new_n996), .B1(new_n1180), .B2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g759(.A1(new_n658), .A2(G319), .ZN(new_n1186));
  OR3_X1    g760(.A1(G401), .A2(G229), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g761(.A(new_n1187), .B1(new_n872), .B2(new_n880), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1188), .A2(new_n953), .ZN(G225));
  INV_X1    g763(.A(G225), .ZN(G308));
endmodule


