//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT66), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g0026(.A1(new_n224), .A2(new_n225), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n202), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n207), .ZN(new_n233));
  AND2_X1   g0033(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NOR4_X1   g0034(.A1(new_n213), .A2(new_n226), .A3(new_n227), .A4(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G226), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT67), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n202), .ZN(new_n248));
  INV_X1    g0048(.A(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT68), .ZN(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n250), .B(new_n254), .Z(G351));
  INV_X1    g0055(.A(G13), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G1), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G50), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n260), .A2(new_n232), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n258), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n262), .B1(new_n206), .B2(G20), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n259), .B1(new_n263), .B2(G50), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n249), .A2(KEYINPUT70), .A3(KEYINPUT8), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT8), .B(G58), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT70), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(new_n207), .A3(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n264), .B1(new_n272), .B2(new_n261), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G169), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n277), .B1(new_n282), .B2(G226), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT69), .B(G223), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G1698), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G222), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n288), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(G77), .B2(new_n288), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n283), .B1(new_n294), .B2(new_n279), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n274), .B1(new_n275), .B2(new_n295), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n295), .A2(G179), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n273), .B(KEYINPUT9), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n295), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(G190), .B2(new_n295), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n301), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n302), .A2(KEYINPUT74), .A3(KEYINPUT10), .A4(new_n305), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n261), .A2(new_n258), .A3(KEYINPUT73), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT73), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n256), .A2(new_n207), .A3(G1), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n260), .A2(new_n232), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n206), .A2(G20), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  MUX2_X1   g0117(.A(new_n258), .B(new_n317), .S(G77), .Z(new_n318));
  INV_X1    g0118(.A(new_n266), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(new_n270), .B1(G20), .B2(G77), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT72), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n207), .A2(G33), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n320), .A2(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n313), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n318), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT3), .B(G33), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(G232), .A3(new_n291), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(G238), .A3(G1698), .ZN(new_n331));
  INV_X1    g0131(.A(G107), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n330), .B(new_n331), .C1(new_n332), .C2(new_n329), .ZN(new_n333));
  INV_X1    g0133(.A(new_n279), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n277), .B1(new_n282), .B2(G244), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G169), .ZN(new_n338));
  INV_X1    g0138(.A(G179), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n337), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n328), .A2(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n335), .A2(new_n336), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(G200), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n337), .A2(G190), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n327), .B(new_n318), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  AND4_X1   g0146(.A1(new_n300), .A2(new_n308), .A3(new_n309), .A4(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n277), .B1(new_n282), .B2(G238), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n329), .A2(G232), .A3(G1698), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G97), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT75), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n291), .A2(G226), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n288), .B2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n329), .A2(KEYINPUT75), .A3(G226), .A4(new_n291), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n348), .B1(new_n356), .B2(new_n279), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT13), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(KEYINPUT76), .A3(KEYINPUT13), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT76), .B1(new_n357), .B2(KEYINPUT13), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G169), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT14), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT14), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(new_n367), .A3(G169), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n357), .A2(KEYINPUT13), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n360), .A2(G179), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n366), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G68), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n317), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT78), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n270), .A2(G50), .B1(G20), .B2(new_n372), .ZN(new_n376));
  INV_X1    g0176(.A(G77), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n324), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n313), .ZN(new_n379));
  XOR2_X1   g0179(.A(KEYINPUT77), .B(KEYINPUT11), .Z(new_n380));
  OR2_X1    g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n380), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n257), .A2(G20), .A3(new_n372), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT12), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n375), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n371), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n386), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n364), .A2(G200), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n360), .A2(G190), .A3(new_n369), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n347), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n329), .B2(G20), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n284), .A2(G33), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT7), .B(new_n207), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n372), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n249), .A2(new_n372), .ZN(new_n400));
  OAI21_X1  g0200(.A(G20), .B1(new_n400), .B2(new_n201), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n270), .A2(G159), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n393), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT81), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT79), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n286), .B2(KEYINPUT3), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n284), .A2(KEYINPUT79), .A3(G33), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n287), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n207), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT7), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n394), .A3(new_n207), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(G68), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n403), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(KEYINPUT16), .A3(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(KEYINPUT81), .B(new_n393), .C1(new_n399), .C2(new_n403), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n406), .A2(new_n416), .A3(new_n313), .A4(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n268), .A2(new_n258), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n263), .B2(new_n268), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n276), .B1(new_n281), .B2(new_n239), .ZN(new_n421));
  AND2_X1   g0221(.A1(G226), .A2(G1698), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(G223), .B2(new_n291), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n410), .A2(new_n423), .B1(new_n286), .B2(new_n215), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n421), .B1(new_n424), .B2(new_n334), .ZN(new_n425));
  INV_X1    g0225(.A(G190), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(G200), .B2(new_n425), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n418), .A2(KEYINPUT84), .A3(new_n420), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT83), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT83), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n418), .A2(new_n431), .A3(new_n420), .A4(new_n428), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(KEYINPUT17), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(KEYINPUT83), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT82), .B1(new_n425), .B2(G169), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n425), .A2(new_n339), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n425), .A2(KEYINPUT82), .A3(new_n339), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n418), .A2(new_n420), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT18), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n438), .A2(new_n439), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n420), .B2(new_n418), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n433), .A2(new_n435), .A3(new_n443), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n206), .A2(G33), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n310), .A2(new_n314), .A3(G116), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G116), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n312), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(G20), .B1(new_n286), .B2(G97), .ZN(new_n454));
  INV_X1    g0254(.A(G283), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n286), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT89), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n451), .A2(G20), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n313), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n457), .B1(new_n313), .B2(new_n458), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(KEYINPUT20), .B(new_n456), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n453), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT5), .B(G41), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(G274), .A3(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n279), .ZN(new_n473));
  INV_X1    g0273(.A(G270), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G264), .A2(G1698), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n218), .B2(G1698), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n477), .A2(new_n408), .A3(new_n409), .A4(new_n287), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n288), .A2(G303), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n279), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n475), .A2(new_n480), .A3(new_n339), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT90), .B1(new_n465), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n463), .A2(new_n464), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n450), .A2(new_n452), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT90), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(new_n481), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n475), .A2(new_n480), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(new_n275), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n486), .A2(KEYINPUT21), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n486), .A2(new_n491), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT21), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n489), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT91), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n465), .B(new_n497), .C1(new_n303), .C2(new_n490), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n490), .A2(new_n303), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT91), .B1(new_n486), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n490), .A2(G190), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n469), .B1(new_n473), .B2(new_n218), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT85), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(KEYINPUT85), .B(new_n469), .C1(new_n473), .C2(new_n218), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n291), .A2(KEYINPUT4), .A3(G244), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n216), .B2(new_n291), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(new_n329), .B1(G33), .B2(G283), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n408), .A2(new_n409), .A3(G244), .A4(new_n287), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(G1698), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n512), .B2(KEYINPUT4), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n506), .A2(new_n507), .B1(new_n513), .B2(new_n334), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n339), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n334), .ZN(new_n516));
  INV_X1    g0316(.A(new_n504), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n275), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n332), .A2(KEYINPUT6), .A3(G97), .ZN(new_n520));
  XOR2_X1   g0320(.A(G97), .B(G107), .Z(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(KEYINPUT6), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(G20), .B1(G77), .B2(new_n270), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n395), .A2(new_n398), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G107), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n313), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n258), .A2(G97), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n261), .A2(new_n258), .A3(new_n449), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n530), .B2(G97), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n515), .A2(new_n519), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n531), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n526), .B2(new_n313), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n516), .A2(G190), .A3(new_n517), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n536), .C1(new_n514), .C2(new_n303), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n207), .A2(G107), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n257), .A2(new_n539), .A3(KEYINPUT25), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n540), .A2(KEYINPUT92), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT25), .B1(new_n257), .B2(new_n539), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n542), .B2(KEYINPUT92), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n541), .A2(new_n543), .B1(new_n530), .B2(G107), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n207), .A2(G87), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n288), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n207), .B2(G107), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n332), .A2(KEYINPUT23), .A3(G20), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n286), .A2(new_n451), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n549), .A2(new_n550), .B1(new_n551), .B2(new_n207), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n408), .A2(new_n409), .A3(new_n207), .A4(new_n287), .ZN(new_n553));
  NAND2_X1  g0353(.A1(KEYINPUT22), .A2(G87), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n547), .B(new_n552), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n313), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n547), .A2(new_n552), .ZN(new_n558));
  OR2_X1    g0358(.A1(new_n553), .A2(new_n554), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT24), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n544), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G257), .A2(G1698), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n216), .B2(G1698), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(new_n408), .A3(new_n409), .A4(new_n287), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G294), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n279), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n472), .A2(G264), .A3(new_n279), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n567), .A2(G179), .A3(new_n569), .A4(new_n469), .ZN(new_n570));
  INV_X1    g0370(.A(new_n469), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n566), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n572), .B2(new_n275), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n561), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n555), .A2(new_n556), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n559), .A2(KEYINPUT24), .A3(new_n547), .A4(new_n552), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n313), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n572), .A2(G200), .ZN(new_n578));
  NOR4_X1   g0378(.A1(new_n566), .A2(new_n568), .A3(new_n571), .A4(G190), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n577), .B(new_n544), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT93), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n574), .A2(new_n580), .A3(KEYINPUT93), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n538), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT87), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n408), .A2(new_n409), .A3(new_n287), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT86), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n207), .A4(G68), .ZN(new_n589));
  OAI21_X1  g0389(.A(KEYINPUT86), .B1(new_n553), .B2(new_n372), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OR2_X1    g0391(.A1(KEYINPUT19), .A2(G20), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(new_n350), .ZN(new_n593));
  NOR2_X1   g0393(.A1(G87), .A2(G97), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n332), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n350), .A2(new_n207), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n593), .B1(new_n597), .B2(KEYINPUT19), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n586), .B1(new_n591), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n598), .B1(new_n589), .B2(new_n590), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n261), .B1(new_n600), .B2(KEYINPUT87), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n325), .A2(new_n312), .ZN(new_n603));
  INV_X1    g0403(.A(new_n325), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n530), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(G250), .B1(new_n467), .B2(G1), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n468), .A2(G274), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n334), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(G238), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n610), .A2(G1698), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n408), .A2(new_n409), .A3(new_n611), .A4(new_n287), .ZN(new_n612));
  OAI221_X1 g0412(.A(new_n612), .B1(new_n286), .B2(new_n451), .C1(new_n511), .C2(new_n291), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n609), .B1(new_n613), .B2(new_n334), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n339), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(G169), .B2(new_n614), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n606), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT88), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n599), .A2(new_n601), .B1(new_n312), .B2(new_n325), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n530), .A2(G87), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n614), .A2(new_n426), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(G200), .B2(new_n614), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n618), .B2(new_n624), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n503), .B(new_n585), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n392), .A2(new_n448), .A3(new_n627), .ZN(G372));
  NOR2_X1   g0428(.A1(new_n392), .A2(new_n448), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n616), .B1(new_n620), .B2(new_n605), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  INV_X1    g0431(.A(new_n533), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n631), .A2(new_n618), .A3(new_n624), .A4(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n495), .A2(new_n492), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(KEYINPUT94), .A3(new_n489), .A4(new_n574), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n489), .A2(new_n492), .A3(new_n495), .A4(new_n574), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT94), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n618), .A2(new_n624), .ZN(new_n640));
  INV_X1    g0440(.A(new_n580), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n640), .A2(new_n641), .A3(new_n538), .ZN(new_n642));
  AOI211_X1 g0442(.A(new_n630), .B(new_n633), .C1(new_n639), .C2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT88), .B1(new_n644), .B2(new_n630), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n631), .B1(new_n647), .B2(new_n632), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n629), .A2(KEYINPUT95), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n300), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n447), .A2(new_n443), .ZN(new_n653));
  INV_X1    g0453(.A(new_n341), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n371), .A2(new_n386), .B1(new_n391), .B2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n429), .A2(KEYINPUT83), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n432), .A2(KEYINPUT17), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n435), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n653), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n308), .A2(new_n309), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n652), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n651), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT95), .B1(new_n629), .B2(new_n650), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n662), .A2(new_n663), .ZN(G369));
  INV_X1    g0464(.A(new_n257), .ZN(new_n665));
  OR3_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .A3(G20), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT27), .B1(new_n665), .B2(G20), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n496), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n583), .A2(new_n584), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n561), .A2(new_n670), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT96), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(KEYINPUT96), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n672), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n574), .A2(new_n670), .ZN(new_n681));
  OR3_X1    g0481(.A1(new_n680), .A2(KEYINPUT97), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT97), .B1(new_n680), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n678), .A2(new_n679), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n561), .A2(new_n573), .A3(new_n670), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n465), .A2(new_n671), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n634), .A2(new_n489), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n503), .B2(new_n688), .ZN(new_n690));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n684), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n210), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n594), .A2(new_n332), .A3(new_n451), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n697), .A2(G1), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n231), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n697), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT31), .B1(new_n627), .B2(new_n670), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT98), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n481), .A2(new_n614), .A3(new_n569), .A4(new_n567), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n518), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT30), .ZN(new_n708));
  NOR4_X1   g0508(.A1(new_n614), .A2(new_n572), .A3(new_n490), .A4(G179), .ZN(new_n709));
  INV_X1    g0509(.A(new_n514), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n707), .A2(KEYINPUT30), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n705), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n713), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(KEYINPUT98), .A3(new_n708), .A4(new_n711), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n671), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n704), .A2(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(KEYINPUT31), .B(new_n670), .C1(new_n712), .C2(new_n713), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n691), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n644), .A2(new_n630), .ZN(new_n723));
  INV_X1    g0523(.A(new_n538), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n723), .A2(new_n580), .A3(new_n724), .A4(new_n636), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT26), .B1(new_n640), .B2(new_n533), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(new_n618), .A3(new_n726), .ZN(new_n727));
  AOI211_X1 g0527(.A(KEYINPUT26), .B(new_n533), .C1(new_n645), .C2(new_n646), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT29), .B(new_n671), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n670), .B1(new_n643), .B2(new_n649), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n722), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n703), .B1(new_n733), .B2(G1), .ZN(G364));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n232), .B1(G20), .B2(new_n275), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n695), .A2(new_n587), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n250), .A2(G45), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n701), .A2(new_n467), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n210), .A2(new_n329), .ZN(new_n745));
  INV_X1    g0545(.A(G355), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n746), .B1(G116), .B2(new_n210), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n739), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n256), .A2(G20), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G45), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n697), .A2(G1), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n207), .A2(G190), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n303), .A2(G179), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n332), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n207), .A2(new_n426), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n339), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n329), .B1(new_n758), .B2(new_n249), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n756), .A2(new_n753), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n755), .B(new_n759), .C1(G87), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G179), .A2(G200), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n207), .B1(new_n763), .B2(G190), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n217), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n752), .A2(new_n763), .ZN(new_n767));
  INV_X1    g0567(.A(G159), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT32), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n339), .A2(new_n303), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n756), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n752), .A2(new_n757), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n772), .A2(new_n202), .B1(new_n773), .B2(new_n377), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n771), .A2(new_n752), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n774), .B1(G68), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n762), .A2(new_n766), .A3(new_n770), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G326), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n772), .A2(new_n779), .B1(new_n773), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n764), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(G294), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT99), .Z(new_n784));
  INV_X1    g0584(.A(new_n754), .ZN(new_n785));
  INV_X1    g0585(.A(new_n767), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G283), .A2(new_n785), .B1(new_n786), .B2(G329), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT100), .ZN(new_n788));
  INV_X1    g0588(.A(G303), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n288), .B1(new_n760), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n758), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(G322), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT33), .B(G317), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n775), .B1(new_n794), .B2(KEYINPUT101), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(KEYINPUT101), .B2(new_n794), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n788), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n778), .B1(new_n784), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n751), .B1(new_n798), .B2(new_n738), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n748), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n690), .B2(new_n737), .ZN(new_n801));
  INV_X1    g0601(.A(new_n751), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n692), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n690), .A2(new_n691), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  OAI22_X1  g0606(.A1(new_n775), .A2(new_n455), .B1(new_n773), .B2(new_n451), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT102), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G294), .A2(new_n791), .B1(new_n786), .B2(G311), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n754), .A2(new_n215), .ZN(new_n810));
  INV_X1    g0610(.A(new_n772), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n810), .B1(G303), .B2(new_n811), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n329), .B(new_n765), .C1(G107), .C2(new_n761), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n808), .A2(new_n809), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G132), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n754), .A2(new_n372), .B1(new_n767), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G50), .B2(new_n761), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n410), .B1(new_n782), .B2(G58), .ZN(new_n818));
  INV_X1    g0618(.A(new_n773), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n811), .A2(G137), .B1(new_n819), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G150), .ZN(new_n821));
  XOR2_X1   g0621(.A(KEYINPUT103), .B(G143), .Z(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n821), .B2(new_n775), .C1(new_n758), .C2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT34), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n817), .B(new_n818), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n814), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n738), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n738), .A2(new_n735), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n751), .B1(new_n377), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n341), .A2(new_n670), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n671), .B1(new_n318), .B2(new_n327), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n832), .A2(KEYINPUT104), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(KEYINPUT104), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(new_n345), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n831), .B1(new_n835), .B2(new_n341), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n828), .B(new_n830), .C1(new_n836), .C2(new_n736), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n730), .A2(new_n836), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT105), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n639), .A2(new_n642), .ZN(new_n840));
  INV_X1    g0640(.A(new_n633), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n840), .A2(new_n618), .A3(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n671), .B(new_n836), .C1(new_n842), .C2(new_n648), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n838), .A2(new_n839), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n839), .B2(new_n838), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n802), .B1(new_n845), .B2(new_n721), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n721), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n837), .B1(new_n847), .B2(new_n848), .ZN(G384));
  NAND2_X1  g0649(.A1(new_n522), .A2(KEYINPUT35), .ZN(new_n850));
  OAI211_X1 g0650(.A(G116), .B(new_n233), .C1(new_n522), .C2(KEYINPUT35), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(KEYINPUT106), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(KEYINPUT106), .B2(new_n851), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT36), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(KEYINPUT36), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n701), .A2(new_n377), .A3(new_n400), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n372), .A2(G50), .ZN(new_n857));
  OAI211_X1 g0657(.A(G1), .B(new_n256), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n854), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT107), .Z(new_n860));
  INV_X1    g0660(.A(new_n836), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n717), .A2(KEYINPUT31), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(new_n719), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n414), .A2(new_n415), .ZN(new_n865));
  INV_X1    g0665(.A(new_n393), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n416), .B(new_n313), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n420), .ZN(new_n868));
  INV_X1    g0668(.A(new_n668), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n429), .A2(KEYINPUT83), .A3(new_n434), .ZN(new_n871));
  INV_X1    g0671(.A(new_n657), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n430), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n870), .B1(new_n873), .B2(new_n653), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n444), .A2(new_n668), .B1(new_n867), .B2(new_n420), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n418), .A2(new_n420), .A3(new_n428), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n441), .A2(new_n869), .ZN(new_n879));
  XNOR2_X1  g0679(.A(KEYINPUT108), .B(KEYINPUT37), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n442), .A2(new_n879), .A3(new_n876), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n864), .B1(new_n874), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n870), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n448), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n882), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n386), .A2(new_n670), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n387), .A2(new_n391), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n391), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n386), .B(new_n670), .C1(new_n891), .C2(new_n371), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n863), .A2(new_n888), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n445), .A2(new_n877), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT110), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(new_n898), .A3(new_n879), .A4(new_n880), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n881), .A2(KEYINPUT110), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n442), .A2(new_n879), .A3(new_n876), .ZN(new_n901));
  INV_X1    g0701(.A(new_n880), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n899), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n879), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n447), .A2(new_n443), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n905), .B1(new_n658), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n864), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n887), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n863), .A2(KEYINPUT40), .A3(new_n910), .A4(new_n893), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n896), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT112), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n719), .A2(new_n862), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n914), .A2(new_n629), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n691), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n915), .B2(new_n913), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n629), .B(new_n729), .C1(new_n730), .C2(KEYINPUT29), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n661), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT111), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n371), .A2(new_n386), .A3(new_n671), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n909), .A2(new_n923), .A3(new_n887), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT109), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n924), .A2(new_n925), .B1(new_n888), .B2(KEYINPUT39), .ZN(new_n926));
  AOI221_X4 g0726(.A(new_n864), .B1(new_n881), .B2(new_n878), .C1(new_n448), .C2(new_n885), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT38), .B1(new_n886), .B2(new_n882), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n925), .B(KEYINPUT39), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n922), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n653), .A2(new_n869), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n890), .A2(new_n892), .ZN(new_n933));
  INV_X1    g0733(.A(new_n831), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n933), .B1(new_n843), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n932), .B1(new_n935), .B2(new_n888), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n920), .B(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n917), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT113), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n940), .B1(new_n206), .B2(new_n749), .C1(new_n938), .C2(new_n917), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n939), .A2(KEYINPUT113), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n860), .B1(new_n941), .B2(new_n942), .ZN(G367));
  OAI21_X1  g0743(.A(new_n724), .B1(new_n535), .B2(new_n671), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n632), .A2(new_n670), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n687), .A2(new_n496), .A3(new_n671), .A4(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT42), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(KEYINPUT42), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n533), .B1(new_n944), .B2(new_n574), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n671), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT43), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n671), .B1(new_n620), .B2(new_n621), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT114), .Z(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(new_n723), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n618), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n952), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n953), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT115), .ZN(new_n961));
  INV_X1    g0761(.A(new_n946), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n693), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n961), .B(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n959), .B(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n696), .B(KEYINPUT41), .Z(new_n966));
  AND3_X1   g0766(.A1(new_n684), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT45), .B1(new_n684), .B2(new_n946), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n682), .A2(new_n683), .A3(new_n962), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT44), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n693), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n692), .B(new_n687), .C1(new_n969), .C2(new_n971), .ZN(new_n974));
  MUX2_X1   g0774(.A(new_n685), .B(new_n687), .S(new_n672), .Z(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(new_n692), .Z(new_n976));
  NAND4_X1  g0776(.A1(new_n973), .A2(new_n974), .A3(new_n733), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n966), .B1(new_n977), .B2(new_n733), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n750), .A2(G1), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT116), .Z(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n965), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n739), .B1(new_n210), .B2(new_n325), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n244), .B2(new_n740), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT117), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n751), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n985), .B2(new_n984), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G50), .A2(new_n819), .B1(new_n785), .B2(G77), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n821), .B2(new_n758), .C1(new_n768), .C2(new_n775), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n764), .A2(new_n372), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n329), .B1(new_n772), .B2(new_n822), .ZN(new_n991));
  INV_X1    g0791(.A(G137), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n760), .A2(new_n249), .B1(new_n767), .B2(new_n992), .ZN(new_n993));
  NOR4_X1   g0793(.A1(new_n989), .A2(new_n990), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT119), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n761), .A2(KEYINPUT46), .A3(G116), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT46), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n760), .B2(new_n451), .ZN(new_n998));
  INV_X1    g0798(.A(G294), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n996), .B(new_n998), .C1(new_n999), .C2(new_n775), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(KEYINPUT118), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(KEYINPUT118), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n410), .B1(new_n754), .B2(new_n217), .C1(new_n789), .C2(new_n758), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G107), .B2(new_n782), .ZN(new_n1004));
  INV_X1    g0804(.A(G317), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n772), .A2(new_n780), .B1(new_n767), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G283), .B2(new_n819), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1002), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n995), .B1(new_n1001), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1010), .A2(KEYINPUT47), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n738), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n1010), .B2(KEYINPUT47), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n987), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n958), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n737), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n982), .A2(new_n1017), .ZN(G387));
  OAI22_X1  g0818(.A1(new_n745), .A2(new_n699), .B1(G107), .B2(new_n210), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n240), .A2(G45), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n266), .A2(G50), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  AOI211_X1 g0822(.A(G45), .B(new_n698), .C1(G68), .C2(G77), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n741), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1019), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n739), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n802), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n687), .A2(new_n1016), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n772), .A2(new_n768), .B1(new_n760), .B2(new_n377), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n758), .A2(new_n202), .B1(new_n773), .B2(new_n372), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n782), .A2(new_n604), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n754), .A2(new_n217), .B1(new_n767), .B2(new_n821), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1033), .A2(new_n410), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n268), .A2(new_n776), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n760), .A2(new_n999), .B1(new_n764), .B2(new_n455), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n773), .A2(new_n789), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n780), .A2(new_n775), .B1(new_n758), .B2(new_n1005), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G322), .C2(new_n811), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1037), .B1(new_n1040), .B2(KEYINPUT48), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(KEYINPUT48), .B2(new_n1040), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT49), .Z(new_n1043));
  OAI221_X1 g0843(.A(new_n410), .B1(new_n767), .B2(new_n779), .C1(new_n451), .C2(new_n754), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1036), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1027), .B(new_n1028), .C1(new_n738), .C2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n976), .B2(new_n981), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n976), .A2(new_n733), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n696), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n976), .A2(new_n733), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1047), .B1(new_n1049), .B2(new_n1050), .ZN(G393));
  NAND2_X1  g0851(.A1(new_n962), .A2(new_n737), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n254), .A2(new_n740), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n739), .B1(new_n217), .B2(new_n210), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n802), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n772), .A2(new_n1005), .B1(new_n758), .B2(new_n780), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT52), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G303), .A2(new_n776), .B1(new_n786), .B2(G322), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G283), .A2(new_n761), .B1(new_n819), .B2(G294), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n329), .B(new_n755), .C1(G116), .C2(new_n782), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n410), .B(new_n810), .C1(new_n319), .C2(new_n819), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n782), .A2(G77), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G50), .A2(new_n776), .B1(new_n761), .B2(G68), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n767), .C2(new_n822), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n772), .A2(new_n821), .B1(new_n758), .B2(new_n768), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT51), .Z(new_n1068));
  OAI21_X1  g0868(.A(new_n1061), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1055), .B1(new_n1069), .B2(new_n738), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1052), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n973), .A2(new_n974), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1071), .B1(new_n1072), .B2(new_n980), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n977), .A2(new_n696), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1048), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(G390));
  NAND3_X1  g0877(.A1(new_n914), .A2(new_n629), .A3(G330), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n918), .A2(new_n1078), .A3(new_n661), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT122), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n863), .A2(G330), .A3(new_n893), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n647), .A2(new_n503), .A3(new_n585), .A4(new_n671), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n717), .B1(new_n1082), .B2(KEYINPUT31), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n720), .ZN(new_n1084));
  OAI211_X1 g0884(.A(G330), .B(new_n836), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1081), .B1(new_n893), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n843), .A2(new_n934), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n721), .A2(KEYINPUT121), .A3(new_n836), .A4(new_n893), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT121), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n1085), .B2(new_n933), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n835), .A2(new_n341), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n671), .B(new_n1094), .C1(new_n727), .C2(new_n728), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n934), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n863), .A2(G330), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n933), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1093), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1080), .B1(new_n1089), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT120), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n921), .B(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n910), .A2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1095), .A2(new_n934), .B1(new_n890), .B2(new_n892), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT38), .B1(new_n904), .B2(new_n907), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n927), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT109), .B1(new_n1107), .B2(new_n923), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n923), .B1(new_n884), .B2(new_n887), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n929), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n922), .B1(new_n1088), .B2(new_n893), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1093), .B(new_n1105), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n924), .A2(new_n925), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1109), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n930), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1088), .A2(new_n893), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n921), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1113), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1112), .B1(new_n1119), .B2(new_n1081), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n697), .B1(new_n1100), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n1120), .B2(new_n1100), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1120), .A2(new_n980), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n829), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n802), .B1(new_n268), .B2(new_n1124), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n772), .A2(new_n455), .B1(new_n754), .B2(new_n372), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n329), .B(new_n1126), .C1(G87), .C2(new_n761), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G107), .A2(new_n776), .B1(new_n791), .B2(G116), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G97), .A2(new_n819), .B1(new_n786), .B2(G294), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1127), .A2(new_n1063), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n775), .A2(new_n992), .B1(new_n773), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G159), .B2(new_n782), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT123), .Z(new_n1134));
  NOR2_X1   g0934(.A1(new_n760), .A2(new_n821), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT53), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n329), .B1(new_n815), .B2(new_n758), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n1136), .B2(new_n1135), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n786), .A2(G125), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G128), .A2(new_n811), .B1(new_n785), .B2(G50), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1130), .B1(new_n1134), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1125), .B1(new_n1142), .B2(new_n738), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n1110), .B2(new_n736), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1122), .A2(new_n1123), .A3(new_n1144), .ZN(G378));
  NAND3_X1  g0945(.A1(new_n896), .A2(G330), .A3(new_n911), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n660), .A2(new_n300), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n274), .A2(new_n668), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n931), .A2(new_n936), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n931), .B2(new_n936), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1147), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1156), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n921), .B1(new_n1161), .B2(new_n929), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1088), .A2(new_n888), .A3(new_n893), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n653), .B2(new_n869), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1160), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n931), .A2(new_n936), .A3(new_n1156), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n1146), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1159), .A2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1093), .A2(new_n1098), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1080), .B1(new_n1120), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n696), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1168), .A2(new_n981), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n751), .B1(new_n202), .B2(new_n829), .ZN(new_n1176));
  INV_X1    g0976(.A(G125), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n772), .A2(new_n1177), .B1(new_n775), .B2(new_n815), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1131), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1179), .A2(new_n761), .B1(new_n791), .B2(G128), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n992), .B2(new_n773), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1178), .B(new_n1181), .C1(G150), .C2(new_n782), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n786), .A2(G124), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G33), .B(G41), .C1(new_n785), .C2(G159), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n773), .A2(new_n325), .B1(new_n767), .B2(new_n455), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n587), .A2(G41), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n217), .C2(new_n775), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n760), .A2(new_n377), .B1(new_n754), .B2(new_n249), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n772), .A2(new_n451), .B1(new_n758), .B2(new_n332), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1192), .A2(new_n990), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT58), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1195), .A2(KEYINPUT58), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1191), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1198), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1199));
  AND4_X1   g0999(.A1(new_n1188), .A2(new_n1196), .A3(new_n1197), .A4(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1176), .B1(new_n1012), .B2(new_n1200), .C1(new_n1160), .C2(new_n736), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1175), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1174), .A2(new_n1203), .ZN(G375));
  OAI22_X1  g1004(.A1(new_n451), .A2(new_n775), .B1(new_n758), .B2(new_n455), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n329), .B(new_n1205), .C1(G77), .C2(new_n785), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G97), .A2(new_n761), .B1(new_n786), .B2(G303), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n811), .A2(G294), .B1(new_n819), .B2(G107), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1206), .A2(new_n1032), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n772), .A2(new_n815), .B1(new_n758), .B2(new_n992), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G159), .B2(new_n761), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G58), .A2(new_n785), .B1(new_n819), .B2(G150), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n776), .A2(new_n1179), .B1(new_n786), .B2(G128), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n410), .B1(new_n782), .B2(G50), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1012), .B1(new_n1209), .B2(new_n1215), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n751), .B(new_n1216), .C1(new_n372), .C2(new_n829), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n893), .B2(new_n736), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1169), .B2(new_n980), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1100), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(new_n966), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1079), .B(KEYINPUT122), .Z(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1169), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1220), .B1(new_n1222), .B2(new_n1225), .ZN(G381));
  AND3_X1   g1026(.A1(new_n1076), .A2(new_n982), .A3(new_n1017), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(G375), .A2(G378), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(G407));
  INV_X1    g1030(.A(G213), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(G343), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1228), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(G407), .A2(G213), .A3(new_n1233), .ZN(G409));
  XNOR2_X1  g1034(.A(G393), .B(new_n805), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1076), .B1(new_n982), .B2(new_n1017), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1235), .B1(new_n1227), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G387), .A2(G390), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1076), .A2(new_n982), .A3(new_n1017), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1235), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(new_n966), .ZN(new_n1244));
  AOI21_X1  g1044(.A(G378), .B1(new_n1203), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1243), .A2(KEYINPUT57), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1202), .B1(new_n1249), .B2(new_n696), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT124), .B1(new_n1250), .B2(G378), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1174), .A2(G378), .A3(KEYINPUT124), .A4(new_n1203), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1246), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT62), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1232), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1224), .A2(KEYINPUT60), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1224), .A2(KEYINPUT60), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1100), .A2(new_n696), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(G384), .A3(new_n1220), .ZN(new_n1263));
  INV_X1    g1063(.A(G384), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1260), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1264), .B1(new_n1265), .B2(new_n1219), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1232), .A2(G2897), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1263), .A2(new_n1266), .A3(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1271), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1174), .A2(G378), .A3(new_n1203), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT124), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1245), .B1(new_n1277), .B2(new_n1252), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1274), .B1(new_n1278), .B2(new_n1232), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1269), .A2(new_n1270), .A3(new_n1279), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1278), .A2(new_n1232), .A3(new_n1267), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(new_n1255), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1242), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1279), .A2(KEYINPUT63), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1254), .A2(new_n1256), .A3(new_n1268), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1237), .A2(new_n1241), .A3(new_n1270), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1281), .B2(KEYINPUT63), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1283), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT125), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT125), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1283), .A2(new_n1289), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(G405));
  INV_X1    g1094(.A(G378), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G375), .A2(new_n1295), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1296), .B(KEYINPUT126), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1277), .A2(new_n1252), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  XOR2_X1   g1099(.A(new_n1299), .B(KEYINPUT127), .Z(new_n1300));
  XNOR2_X1  g1100(.A(new_n1242), .B(new_n1267), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1300), .B(new_n1301), .ZN(G402));
endmodule


