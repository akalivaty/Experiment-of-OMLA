

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U553 ( .A(KEYINPUT92), .ZN(n682) );
  XNOR2_X1 U554 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U555 ( .A1(n692), .A2(n970), .ZN(n685) );
  NOR2_X1 U556 ( .A1(n719), .A2(n718), .ZN(n720) );
  INV_X1 U557 ( .A(KEYINPUT97), .ZN(n721) );
  XNOR2_X1 U558 ( .A(n722), .B(n721), .ZN(n728) );
  NOR2_X2 U559 ( .A1(n534), .A2(G2105), .ZN(n892) );
  INV_X1 U560 ( .A(G651), .ZN(n525) );
  NOR2_X1 U561 ( .A1(G543), .A2(n525), .ZN(n521) );
  XNOR2_X1 U562 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n520) );
  XNOR2_X1 U563 ( .A(n521), .B(n520), .ZN(n638) );
  NAND2_X1 U564 ( .A1(G64), .A2(n638), .ZN(n524) );
  XOR2_X1 U565 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  NOR2_X1 U566 ( .A1(n634), .A2(G651), .ZN(n522) );
  XOR2_X1 U567 ( .A(KEYINPUT65), .B(n522), .Z(n645) );
  NAND2_X1 U568 ( .A1(G52), .A2(n645), .ZN(n523) );
  NAND2_X1 U569 ( .A1(n524), .A2(n523), .ZN(n530) );
  NOR2_X1 U570 ( .A1(G543), .A2(G651), .ZN(n637) );
  NAND2_X1 U571 ( .A1(G90), .A2(n637), .ZN(n527) );
  NOR2_X1 U572 ( .A1(n634), .A2(n525), .ZN(n641) );
  NAND2_X1 U573 ( .A1(G77), .A2(n641), .ZN(n526) );
  NAND2_X1 U574 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U575 ( .A(KEYINPUT9), .B(n528), .Z(n529) );
  NOR2_X1 U576 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U577 ( .A(KEYINPUT69), .B(n531), .Z(G171) );
  INV_X1 U578 ( .A(G171), .ZN(G301) );
  AND2_X1 U579 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U580 ( .A(G2104), .B(KEYINPUT66), .Z(n534) );
  AND2_X1 U581 ( .A1(G2105), .A2(n534), .ZN(n895) );
  NAND2_X1 U582 ( .A1(n895), .A2(G123), .ZN(n533) );
  XNOR2_X1 U583 ( .A(KEYINPUT18), .B(KEYINPUT76), .ZN(n532) );
  XNOR2_X1 U584 ( .A(n533), .B(n532), .ZN(n542) );
  AND2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n897) );
  NAND2_X1 U586 ( .A1(G111), .A2(n897), .ZN(n536) );
  NAND2_X1 U587 ( .A1(G99), .A2(n892), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n540) );
  NOR2_X1 U589 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  XOR2_X2 U590 ( .A(KEYINPUT17), .B(n537), .Z(n891) );
  NAND2_X1 U591 ( .A1(G135), .A2(n891), .ZN(n538) );
  XNOR2_X1 U592 ( .A(KEYINPUT77), .B(n538), .ZN(n539) );
  NOR2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n542), .A2(n541), .ZN(n923) );
  XNOR2_X1 U595 ( .A(G2096), .B(n923), .ZN(n543) );
  OR2_X1 U596 ( .A1(G2100), .A2(n543), .ZN(G156) );
  INV_X1 U597 ( .A(G132), .ZN(G219) );
  INV_X1 U598 ( .A(G82), .ZN(G220) );
  INV_X1 U599 ( .A(G120), .ZN(G236) );
  INV_X1 U600 ( .A(G69), .ZN(G235) );
  INV_X1 U601 ( .A(G108), .ZN(G238) );
  NAND2_X1 U602 ( .A1(n891), .A2(G138), .ZN(n546) );
  NAND2_X1 U603 ( .A1(G114), .A2(n897), .ZN(n544) );
  XOR2_X1 U604 ( .A(KEYINPUT83), .B(n544), .Z(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G126), .A2(n895), .ZN(n548) );
  NAND2_X1 U607 ( .A1(G102), .A2(n892), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U609 ( .A1(n550), .A2(n549), .ZN(G164) );
  NAND2_X1 U610 ( .A1(G101), .A2(n892), .ZN(n551) );
  XOR2_X1 U611 ( .A(KEYINPUT23), .B(n551), .Z(n553) );
  NAND2_X1 U612 ( .A1(n897), .A2(G113), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n790) );
  NAND2_X1 U614 ( .A1(G125), .A2(n895), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G137), .A2(n891), .ZN(n554) );
  NAND2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n673) );
  NOR2_X1 U617 ( .A1(n790), .A2(n673), .ZN(G160) );
  XOR2_X1 U618 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n557) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n557), .B(n556), .ZN(G223) );
  INV_X1 U621 ( .A(G223), .ZN(n836) );
  NAND2_X1 U622 ( .A1(n836), .A2(G567), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT11), .B(n558), .Z(G234) );
  NAND2_X1 U624 ( .A1(n638), .A2(G56), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT14), .ZN(n561) );
  NAND2_X1 U626 ( .A1(G43), .A2(n645), .ZN(n560) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n637), .A2(G81), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U630 ( .A1(G68), .A2(n641), .ZN(n563) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT72), .B(n565), .Z(n566) );
  XNOR2_X1 U633 ( .A(KEYINPUT13), .B(n566), .ZN(n567) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n978) );
  NAND2_X1 U635 ( .A1(n978), .A2(G860), .ZN(G153) );
  NAND2_X1 U636 ( .A1(G868), .A2(G301), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G79), .A2(n641), .ZN(n570) );
  NAND2_X1 U638 ( .A1(G54), .A2(n645), .ZN(n569) );
  NAND2_X1 U639 ( .A1(n570), .A2(n569), .ZN(n575) );
  NAND2_X1 U640 ( .A1(G92), .A2(n637), .ZN(n572) );
  NAND2_X1 U641 ( .A1(G66), .A2(n638), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U643 ( .A(KEYINPUT73), .B(n573), .Z(n574) );
  NOR2_X1 U644 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U645 ( .A(KEYINPUT15), .B(n576), .ZN(n970) );
  INV_X1 U646 ( .A(G868), .ZN(n604) );
  NAND2_X1 U647 ( .A1(n970), .A2(n604), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n578), .A2(n577), .ZN(G284) );
  NAND2_X1 U649 ( .A1(n638), .A2(G63), .ZN(n579) );
  XNOR2_X1 U650 ( .A(n579), .B(KEYINPUT74), .ZN(n581) );
  NAND2_X1 U651 ( .A1(G51), .A2(n645), .ZN(n580) );
  NAND2_X1 U652 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U653 ( .A(KEYINPUT6), .B(n582), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n637), .A2(G89), .ZN(n583) );
  XNOR2_X1 U655 ( .A(n583), .B(KEYINPUT4), .ZN(n585) );
  NAND2_X1 U656 ( .A1(G76), .A2(n641), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U658 ( .A(n586), .B(KEYINPUT5), .Z(n587) );
  NOR2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U660 ( .A(KEYINPUT7), .B(n589), .Z(n590) );
  XOR2_X1 U661 ( .A(KEYINPUT75), .B(n590), .Z(G168) );
  XOR2_X1 U662 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U663 ( .A1(G78), .A2(n641), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G65), .A2(n638), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n637), .A2(G91), .ZN(n593) );
  XOR2_X1 U667 ( .A(KEYINPUT70), .B(n593), .Z(n594) );
  NOR2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n645), .A2(G53), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(G299) );
  NOR2_X1 U671 ( .A1(G286), .A2(n604), .ZN(n599) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n599), .A2(n598), .ZN(G297) );
  INV_X1 U674 ( .A(G860), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n600), .A2(G559), .ZN(n601) );
  INV_X1 U676 ( .A(n970), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n601), .A2(n607), .ZN(n602) );
  XNOR2_X1 U678 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U679 ( .A1(n607), .A2(G868), .ZN(n603) );
  NOR2_X1 U680 ( .A1(G559), .A2(n603), .ZN(n606) );
  AND2_X1 U681 ( .A1(n604), .A2(n978), .ZN(n605) );
  NOR2_X1 U682 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G559), .A2(n607), .ZN(n608) );
  XOR2_X1 U684 ( .A(n978), .B(n608), .Z(n655) );
  NOR2_X1 U685 ( .A1(n655), .A2(G860), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G67), .A2(n638), .ZN(n610) );
  NAND2_X1 U687 ( .A1(G55), .A2(n645), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G93), .A2(n637), .ZN(n612) );
  NAND2_X1 U690 ( .A1(G80), .A2(n641), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n657) );
  XNOR2_X1 U693 ( .A(n615), .B(n657), .ZN(G145) );
  NAND2_X1 U694 ( .A1(G85), .A2(n637), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G72), .A2(n641), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G60), .A2(n638), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G47), .A2(n645), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U701 ( .A(KEYINPUT68), .B(n622), .Z(G290) );
  NAND2_X1 U702 ( .A1(n638), .A2(G62), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n623), .B(KEYINPUT78), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G50), .A2(n645), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U706 ( .A(KEYINPUT79), .B(n626), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G88), .A2(n637), .ZN(n628) );
  NAND2_X1 U708 ( .A1(G75), .A2(n641), .ZN(n627) );
  AND2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(G303) );
  INV_X1 U711 ( .A(G303), .ZN(G166) );
  NAND2_X1 U712 ( .A1(G49), .A2(n645), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U715 ( .A1(n638), .A2(n633), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n634), .A2(G87), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U718 ( .A1(G86), .A2(n637), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G61), .A2(n638), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n641), .A2(G73), .ZN(n642) );
  XOR2_X1 U722 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n645), .A2(G48), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(G305) );
  XNOR2_X1 U726 ( .A(G290), .B(G166), .ZN(n654) );
  INV_X1 U727 ( .A(G299), .ZN(n974) );
  XNOR2_X1 U728 ( .A(n974), .B(n657), .ZN(n652) );
  XNOR2_X1 U729 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n649) );
  XNOR2_X1 U730 ( .A(G288), .B(KEYINPUT80), .ZN(n648) );
  XNOR2_X1 U731 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U732 ( .A(n650), .B(G305), .Z(n651) );
  XNOR2_X1 U733 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n654), .B(n653), .ZN(n906) );
  XNOR2_X1 U735 ( .A(n655), .B(n906), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n656), .A2(G868), .ZN(n659) );
  OR2_X1 U737 ( .A1(n657), .A2(G868), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2078), .A2(G2084), .ZN(n660) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n661), .ZN(n662) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U745 ( .A1(G235), .A2(G236), .ZN(n664) );
  XOR2_X1 U746 ( .A(KEYINPUT82), .B(n664), .Z(n665) );
  NOR2_X1 U747 ( .A1(G238), .A2(n665), .ZN(n666) );
  NAND2_X1 U748 ( .A1(G57), .A2(n666), .ZN(n840) );
  NAND2_X1 U749 ( .A1(n840), .A2(G567), .ZN(n671) );
  NOR2_X1 U750 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U751 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U752 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U753 ( .A1(G96), .A2(n669), .ZN(n841) );
  NAND2_X1 U754 ( .A1(n841), .A2(G2106), .ZN(n670) );
  NAND2_X1 U755 ( .A1(n671), .A2(n670), .ZN(n842) );
  NAND2_X1 U756 ( .A1(G483), .A2(G661), .ZN(n672) );
  NOR2_X1 U757 ( .A1(n842), .A2(n672), .ZN(n839) );
  NAND2_X1 U758 ( .A1(n839), .A2(G36), .ZN(G176) );
  INV_X1 U759 ( .A(G40), .ZN(n674) );
  OR2_X1 U760 ( .A1(n674), .A2(n673), .ZN(n789) );
  NOR2_X1 U761 ( .A1(n790), .A2(n789), .ZN(n676) );
  NOR2_X1 U762 ( .A1(G164), .A2(G1384), .ZN(n792) );
  AND2_X1 U763 ( .A1(n676), .A2(n792), .ZN(n677) );
  XNOR2_X1 U764 ( .A(n677), .B(KEYINPUT64), .ZN(n679) );
  NAND2_X1 U765 ( .A1(G1996), .A2(n679), .ZN(n678) );
  XNOR2_X1 U766 ( .A(n678), .B(KEYINPUT26), .ZN(n681) );
  INV_X1 U767 ( .A(n679), .ZN(n686) );
  NAND2_X1 U768 ( .A1(G1341), .A2(n686), .ZN(n680) );
  NAND2_X1 U769 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U770 ( .A1(n978), .A2(n684), .ZN(n692) );
  XNOR2_X1 U771 ( .A(n685), .B(KEYINPUT93), .ZN(n691) );
  INV_X1 U772 ( .A(n686), .ZN(n706) );
  NAND2_X1 U773 ( .A1(G2067), .A2(n706), .ZN(n688) );
  NAND2_X1 U774 ( .A1(n686), .A2(G1348), .ZN(n687) );
  NAND2_X1 U775 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U776 ( .A(KEYINPUT94), .B(n689), .ZN(n690) );
  NAND2_X1 U777 ( .A1(n691), .A2(n690), .ZN(n695) );
  NAND2_X1 U778 ( .A1(n970), .A2(n692), .ZN(n693) );
  XOR2_X1 U779 ( .A(KEYINPUT95), .B(n693), .Z(n694) );
  NAND2_X1 U780 ( .A1(n695), .A2(n694), .ZN(n700) );
  NAND2_X1 U781 ( .A1(G2072), .A2(n706), .ZN(n696) );
  XNOR2_X1 U782 ( .A(n696), .B(KEYINPUT27), .ZN(n698) );
  INV_X1 U783 ( .A(G1956), .ZN(n1010) );
  NOR2_X1 U784 ( .A1(n706), .A2(n1010), .ZN(n697) );
  NOR2_X1 U785 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U786 ( .A1(n974), .A2(n701), .ZN(n699) );
  NAND2_X1 U787 ( .A1(n700), .A2(n699), .ZN(n704) );
  NOR2_X1 U788 ( .A1(n974), .A2(n701), .ZN(n702) );
  XOR2_X1 U789 ( .A(n702), .B(KEYINPUT28), .Z(n703) );
  NAND2_X1 U790 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U791 ( .A(n705), .B(KEYINPUT29), .ZN(n710) );
  XOR2_X1 U792 ( .A(KEYINPUT25), .B(G2078), .Z(n954) );
  NOR2_X1 U793 ( .A1(n686), .A2(n954), .ZN(n708) );
  NOR2_X1 U794 ( .A1(G1961), .A2(n706), .ZN(n707) );
  NOR2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n714) );
  NOR2_X1 U796 ( .A1(G301), .A2(n714), .ZN(n709) );
  NOR2_X1 U797 ( .A1(n710), .A2(n709), .ZN(n719) );
  NAND2_X1 U798 ( .A1(n686), .A2(G8), .ZN(n765) );
  NOR2_X1 U799 ( .A1(G1966), .A2(n765), .ZN(n734) );
  NOR2_X1 U800 ( .A1(n686), .A2(G2084), .ZN(n731) );
  NOR2_X1 U801 ( .A1(n734), .A2(n731), .ZN(n711) );
  NAND2_X1 U802 ( .A1(G8), .A2(n711), .ZN(n712) );
  XNOR2_X1 U803 ( .A(KEYINPUT30), .B(n712), .ZN(n713) );
  NOR2_X1 U804 ( .A1(G168), .A2(n713), .ZN(n716) );
  AND2_X1 U805 ( .A1(G301), .A2(n714), .ZN(n715) );
  NOR2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U807 ( .A(n717), .B(KEYINPUT31), .ZN(n718) );
  XOR2_X1 U808 ( .A(KEYINPUT96), .B(n720), .Z(n733) );
  NAND2_X1 U809 ( .A1(n733), .A2(G286), .ZN(n722) );
  NOR2_X1 U810 ( .A1(G1971), .A2(n765), .ZN(n723) );
  XNOR2_X1 U811 ( .A(n723), .B(KEYINPUT98), .ZN(n725) );
  NOR2_X1 U812 ( .A1(n686), .A2(G2090), .ZN(n724) );
  NOR2_X1 U813 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U814 ( .A1(G303), .A2(n726), .ZN(n727) );
  NAND2_X1 U815 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U816 ( .A1(n729), .A2(G8), .ZN(n730) );
  XNOR2_X1 U817 ( .A(n730), .B(KEYINPUT32), .ZN(n764) );
  NAND2_X1 U818 ( .A1(G8), .A2(n731), .ZN(n732) );
  XOR2_X1 U819 ( .A(KEYINPUT91), .B(n732), .Z(n737) );
  INV_X1 U820 ( .A(n733), .ZN(n735) );
  NOR2_X1 U821 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U822 ( .A1(n737), .A2(n736), .ZN(n762) );
  NAND2_X1 U823 ( .A1(G288), .A2(G1976), .ZN(n738) );
  XOR2_X1 U824 ( .A(KEYINPUT100), .B(n738), .Z(n980) );
  INV_X1 U825 ( .A(n980), .ZN(n739) );
  AND2_X1 U826 ( .A1(n762), .A2(n739), .ZN(n745) );
  XNOR2_X1 U827 ( .A(G1981), .B(KEYINPUT101), .ZN(n740) );
  XNOR2_X1 U828 ( .A(n740), .B(G305), .ZN(n991) );
  NOR2_X1 U829 ( .A1(G288), .A2(G1976), .ZN(n741) );
  XNOR2_X1 U830 ( .A(n741), .B(KEYINPUT99), .ZN(n747) );
  NOR2_X1 U831 ( .A1(n765), .A2(n747), .ZN(n742) );
  NAND2_X1 U832 ( .A1(KEYINPUT33), .A2(n742), .ZN(n743) );
  NAND2_X1 U833 ( .A1(n991), .A2(n743), .ZN(n753) );
  INV_X1 U834 ( .A(n753), .ZN(n744) );
  AND2_X1 U835 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U836 ( .A1(n764), .A2(n746), .ZN(n761) );
  INV_X1 U837 ( .A(n747), .ZN(n749) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U839 ( .A1(n749), .A2(n748), .ZN(n987) );
  OR2_X1 U840 ( .A1(n987), .A2(n765), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n980), .A2(n750), .ZN(n751) );
  NOR2_X1 U842 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n759) );
  NOR2_X1 U844 ( .A1(G1981), .A2(G305), .ZN(n756) );
  XNOR2_X1 U845 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n754) );
  XNOR2_X1 U846 ( .A(n754), .B(KEYINPUT89), .ZN(n755) );
  XNOR2_X1 U847 ( .A(n756), .B(n755), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n757), .A2(n765), .ZN(n758) );
  NOR2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n760) );
  AND2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n772) );
  AND2_X1 U851 ( .A1(n762), .A2(n765), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n770) );
  INV_X1 U853 ( .A(n765), .ZN(n768) );
  NOR2_X1 U854 ( .A1(G2090), .A2(G303), .ZN(n766) );
  NAND2_X1 U855 ( .A1(G8), .A2(n766), .ZN(n767) );
  OR2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n769) );
  AND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n810) );
  NAND2_X1 U859 ( .A1(G107), .A2(n897), .ZN(n774) );
  NAND2_X1 U860 ( .A1(G119), .A2(n895), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G131), .A2(n891), .ZN(n776) );
  NAND2_X1 U863 ( .A1(G95), .A2(n892), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U865 ( .A1(n778), .A2(n777), .ZN(n872) );
  INV_X1 U866 ( .A(G1991), .ZN(n947) );
  NOR2_X1 U867 ( .A1(n872), .A2(n947), .ZN(n788) );
  NAND2_X1 U868 ( .A1(G105), .A2(n892), .ZN(n779) );
  XNOR2_X1 U869 ( .A(n779), .B(KEYINPUT38), .ZN(n786) );
  NAND2_X1 U870 ( .A1(G117), .A2(n897), .ZN(n781) );
  NAND2_X1 U871 ( .A1(G141), .A2(n891), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U873 ( .A1(G129), .A2(n895), .ZN(n782) );
  XNOR2_X1 U874 ( .A(KEYINPUT87), .B(n782), .ZN(n783) );
  NOR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n884) );
  AND2_X1 U877 ( .A1(n884), .A2(G1996), .ZN(n787) );
  NOR2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n929) );
  OR2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n822) );
  INV_X1 U881 ( .A(n822), .ZN(n793) );
  NOR2_X1 U882 ( .A1(n929), .A2(n793), .ZN(n814) );
  XOR2_X1 U883 ( .A(n814), .B(KEYINPUT88), .Z(n808) );
  XNOR2_X1 U884 ( .A(G1986), .B(G290), .ZN(n794) );
  XNOR2_X1 U885 ( .A(n794), .B(KEYINPUT84), .ZN(n989) );
  NAND2_X1 U886 ( .A1(n989), .A2(n822), .ZN(n795) );
  XOR2_X1 U887 ( .A(KEYINPUT85), .B(n795), .Z(n806) );
  NAND2_X1 U888 ( .A1(G116), .A2(n897), .ZN(n797) );
  NAND2_X1 U889 ( .A1(G128), .A2(n895), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U891 ( .A(n798), .B(KEYINPUT35), .ZN(n803) );
  NAND2_X1 U892 ( .A1(G140), .A2(n891), .ZN(n800) );
  NAND2_X1 U893 ( .A1(G104), .A2(n892), .ZN(n799) );
  NAND2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U895 ( .A(KEYINPUT34), .B(n801), .Z(n802) );
  NAND2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U897 ( .A(n804), .B(KEYINPUT36), .ZN(n888) );
  XOR2_X1 U898 ( .A(G2067), .B(KEYINPUT37), .Z(n819) );
  NAND2_X1 U899 ( .A1(n888), .A2(n819), .ZN(n805) );
  XOR2_X1 U900 ( .A(KEYINPUT86), .B(n805), .Z(n939) );
  NAND2_X1 U901 ( .A1(n822), .A2(n939), .ZN(n817) );
  AND2_X1 U902 ( .A1(n806), .A2(n817), .ZN(n807) );
  AND2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n825) );
  NOR2_X1 U905 ( .A1(n884), .A2(G1996), .ZN(n811) );
  XNOR2_X1 U906 ( .A(n811), .B(KEYINPUT102), .ZN(n931) );
  AND2_X1 U907 ( .A1(n947), .A2(n872), .ZN(n926) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n926), .A2(n812), .ZN(n813) );
  NOR2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U911 ( .A1(n931), .A2(n815), .ZN(n816) );
  XNOR2_X1 U912 ( .A(KEYINPUT39), .B(n816), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n888), .A2(n819), .ZN(n820) );
  XNOR2_X1 U915 ( .A(n820), .B(KEYINPUT103), .ZN(n936) );
  NAND2_X1 U916 ( .A1(n821), .A2(n936), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U920 ( .A(G1348), .B(G2454), .ZN(n827) );
  XNOR2_X1 U921 ( .A(n827), .B(G2430), .ZN(n828) );
  XNOR2_X1 U922 ( .A(n828), .B(G1341), .ZN(n834) );
  XOR2_X1 U923 ( .A(G2443), .B(G2427), .Z(n830) );
  XNOR2_X1 U924 ( .A(G2438), .B(G2446), .ZN(n829) );
  XNOR2_X1 U925 ( .A(n830), .B(n829), .ZN(n832) );
  XOR2_X1 U926 ( .A(G2451), .B(G2435), .Z(n831) );
  XNOR2_X1 U927 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U928 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n835), .A2(G14), .ZN(n911) );
  XOR2_X1 U930 ( .A(KEYINPUT104), .B(n911), .Z(G401) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U933 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U935 ( .A1(n839), .A2(n838), .ZN(G188) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  NOR2_X1 U938 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  INV_X1 U940 ( .A(n842), .ZN(G319) );
  XOR2_X1 U941 ( .A(KEYINPUT108), .B(G1981), .Z(n844) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U944 ( .A(n845), .B(KEYINPUT41), .Z(n847) );
  XNOR2_X1 U945 ( .A(G1971), .B(G1976), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U947 ( .A(G1956), .B(G1961), .Z(n849) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1966), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U950 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U951 ( .A(KEYINPUT107), .B(G2474), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(G229) );
  XOR2_X1 U953 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U954 ( .A(KEYINPUT105), .B(G2678), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U956 ( .A(KEYINPUT42), .B(G2090), .Z(n857) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U959 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U960 ( .A(G2096), .B(G2100), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n863) );
  XOR2_X1 U962 ( .A(G2078), .B(G2084), .Z(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(G227) );
  NAND2_X1 U964 ( .A1(G112), .A2(n897), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G100), .A2(n892), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n871) );
  NAND2_X1 U967 ( .A1(n895), .A2(G124), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G136), .A2(n891), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U971 ( .A(KEYINPUT109), .B(n869), .Z(n870) );
  NOR2_X1 U972 ( .A1(n871), .A2(n870), .ZN(G162) );
  XOR2_X1 U973 ( .A(KEYINPUT48), .B(KEYINPUT111), .Z(n874) );
  XNOR2_X1 U974 ( .A(n872), .B(KEYINPUT46), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n883) );
  NAND2_X1 U976 ( .A1(G118), .A2(n897), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G130), .A2(n895), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G142), .A2(n891), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G106), .A2(n892), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U982 ( .A(n879), .B(KEYINPUT45), .Z(n880) );
  NOR2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U984 ( .A(n883), .B(n882), .Z(n887) );
  XNOR2_X1 U985 ( .A(G160), .B(n884), .ZN(n885) );
  XNOR2_X1 U986 ( .A(n885), .B(n923), .ZN(n886) );
  XOR2_X1 U987 ( .A(n887), .B(n886), .Z(n890) );
  XNOR2_X1 U988 ( .A(G164), .B(n888), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n904) );
  NAND2_X1 U990 ( .A1(G139), .A2(n891), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G103), .A2(n892), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n902) );
  NAND2_X1 U993 ( .A1(n895), .A2(G127), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n896), .B(KEYINPUT110), .ZN(n899) );
  NAND2_X1 U995 ( .A1(G115), .A2(n897), .ZN(n898) );
  NAND2_X1 U996 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n900), .Z(n901) );
  NOR2_X1 U998 ( .A1(n902), .A2(n901), .ZN(n918) );
  XOR2_X1 U999 ( .A(n918), .B(G162), .Z(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1002 ( .A(G286), .B(n970), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1004 ( .A(n978), .B(G171), .Z(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G397) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n911), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1015 ( .A(G164), .B(G2078), .Z(n917) );
  XNOR2_X1 U1016 ( .A(KEYINPUT116), .B(n917), .ZN(n921) );
  XOR2_X1 U1017 ( .A(n918), .B(KEYINPUT115), .Z(n919) );
  XOR2_X1 U1018 ( .A(G2072), .B(n919), .Z(n920) );
  NOR2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1020 ( .A(KEYINPUT50), .B(n922), .Z(n942) );
  XNOR2_X1 U1021 ( .A(G160), .B(G2084), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(n927), .B(KEYINPUT112), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n935) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1028 ( .A(KEYINPUT113), .B(n932), .Z(n933) );
  XNOR2_X1 U1029 ( .A(n933), .B(KEYINPUT51), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1033 ( .A(KEYINPUT114), .B(n940), .Z(n941) );
  NOR2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n943), .ZN(n944) );
  XNOR2_X1 U1036 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n966) );
  NAND2_X1 U1037 ( .A1(n944), .A2(n966), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n945), .A2(G29), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(KEYINPUT118), .B(n946), .ZN(n1029) );
  XNOR2_X1 U1040 ( .A(G25), .B(n947), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n948), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1042 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(G2072), .B(G33), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(n951), .B(KEYINPUT119), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n958) );
  XNOR2_X1 U1047 ( .A(G1996), .B(G32), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(G27), .B(n954), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(n959), .B(KEYINPUT53), .ZN(n962) );
  XOR2_X1 U1052 ( .A(G2084), .B(G34), .Z(n960) );
  XNOR2_X1 U1053 ( .A(KEYINPUT54), .B(n960), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(G35), .B(G2090), .ZN(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(n966), .B(n965), .ZN(n967) );
  NOR2_X1 U1058 ( .A1(G29), .A2(n967), .ZN(n968) );
  XOR2_X1 U1059 ( .A(KEYINPUT120), .B(n968), .Z(n969) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n969), .ZN(n1027) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .ZN(n997) );
  XNOR2_X1 U1062 ( .A(n970), .B(G1348), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(n971), .B(KEYINPUT121), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(G1971), .A2(G303), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n985) );
  XNOR2_X1 U1066 ( .A(n974), .B(KEYINPUT122), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n975), .B(n1010), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(G1961), .B(G301), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n983) );
  XNOR2_X1 U1070 ( .A(n978), .B(G1341), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n979), .B(KEYINPUT123), .ZN(n981) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(KEYINPUT124), .B(n990), .ZN(n995) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G168), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(KEYINPUT57), .B(n993), .ZN(n994) );
  NAND2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1082 ( .A1(n997), .A2(n996), .ZN(n1025) );
  INV_X1 U1083 ( .A(G16), .ZN(n1023) );
  XOR2_X1 U1084 ( .A(G1986), .B(KEYINPUT127), .Z(n998) );
  XNOR2_X1 U1085 ( .A(G24), .B(n998), .ZN(n1003) );
  XNOR2_X1 U1086 ( .A(G1971), .B(G22), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(G1976), .B(G23), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(KEYINPUT126), .B(n1001), .Z(n1002) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(KEYINPUT58), .B(n1004), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(G1961), .B(G5), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1020) );
  XNOR2_X1 U1096 ( .A(KEYINPUT59), .B(G1348), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(n1009), .B(G4), .ZN(n1016) );
  XOR2_X1 U1098 ( .A(G1341), .B(G19), .Z(n1012) );
  XNOR2_X1 U1099 ( .A(n1010), .B(G20), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G6), .B(G1981), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1017), .Z(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT125), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1111 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

