//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  OAI21_X1  g0004(.A(G50), .B1(G58), .B2(G68), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n217), .A2(new_n218), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n210), .B(new_n214), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0026(.A(G238), .B(G244), .Z(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XOR2_X1   g0037(.A(G58), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n207), .B1(new_n211), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n208), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n251), .A2(new_n252), .B1(new_n208), .B2(G68), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n246), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n254), .B(KEYINPUT11), .Z(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT67), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n259), .A2(new_n256), .A3(G13), .A4(G20), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT74), .ZN(new_n262));
  INV_X1    g0062(.A(G68), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT12), .A4(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n246), .B1(new_n258), .B2(new_n260), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n256), .A2(G20), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT68), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n267), .A3(G68), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT74), .B(KEYINPUT12), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n258), .A2(new_n260), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n269), .B1(new_n270), .B2(G68), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n264), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n255), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT14), .ZN(new_n275));
  AND2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  OAI211_X1 g0077(.A(G232), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT72), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n281), .A2(KEYINPUT72), .A3(G232), .A4(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G97), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n281), .A2(G226), .A3(new_n284), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n280), .A2(new_n282), .A3(new_n283), .A4(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT13), .ZN(new_n291));
  INV_X1    g0091(.A(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  AOI21_X1  g0093(.A(G1), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(new_n288), .A3(G274), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT73), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT73), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n294), .A2(new_n288), .A3(new_n297), .A4(G274), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n289), .A2(new_n294), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n296), .A2(new_n298), .B1(new_n299), .B2(G238), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n290), .A2(new_n291), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n291), .B1(new_n290), .B2(new_n300), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n275), .B(G169), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n290), .A2(new_n300), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT13), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G179), .A3(new_n301), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n306), .B2(new_n301), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT75), .B1(new_n310), .B2(new_n275), .ZN(new_n311));
  OAI21_X1  g0111(.A(G169), .B1(new_n302), .B2(new_n303), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT75), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT14), .ZN(new_n314));
  AOI211_X1 g0114(.A(KEYINPUT76), .B(new_n308), .C1(new_n311), .C2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT76), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n311), .A2(new_n314), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n304), .A2(new_n307), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n274), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(G200), .B1(new_n302), .B2(new_n303), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n306), .A2(G190), .A3(new_n301), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(new_n273), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n324), .A2(KEYINPUT77), .ZN(new_n325));
  INV_X1    g0125(.A(new_n295), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(G226), .B2(new_n299), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n281), .A2(G1698), .ZN(new_n328));
  INV_X1    g0128(.A(G223), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n328), .A2(new_n329), .B1(new_n252), .B2(new_n281), .ZN(new_n330));
  OR2_X1    g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NAND2_X1  g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  AOI21_X1  g0132(.A(G1698), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(G222), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n327), .B1(new_n334), .B2(new_n288), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT10), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n335), .A2(new_n336), .B1(KEYINPUT71), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(G200), .B2(new_n335), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT9), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  INV_X1    g0141(.A(G150), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n341), .A2(new_n251), .B1(new_n342), .B2(new_n248), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G58), .A2(G68), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n208), .B1(new_n344), .B2(new_n249), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n246), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n265), .A2(new_n267), .A3(G50), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n346), .B(new_n347), .C1(G50), .C2(new_n270), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT70), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n339), .B1(new_n340), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n340), .B2(new_n349), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n337), .A2(KEYINPUT71), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n351), .B(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n335), .A2(new_n309), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n354), .B(new_n348), .C1(G179), .C2(new_n335), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n333), .A2(G223), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n281), .A2(G226), .A3(G1698), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G87), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n289), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n326), .B1(G232), .B2(new_n299), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n361), .A2(G190), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G200), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n361), .B2(new_n362), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n246), .ZN(new_n367));
  INV_X1    g0167(.A(G58), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(new_n263), .ZN(new_n369));
  OAI21_X1  g0169(.A(G20), .B1(new_n369), .B2(new_n344), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n247), .A2(G159), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n276), .A2(new_n277), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n208), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n263), .B1(new_n374), .B2(KEYINPUT7), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n281), .A2(G20), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n372), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n367), .B1(new_n379), .B2(KEYINPUT16), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT16), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n376), .A2(KEYINPUT7), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n374), .A2(new_n377), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n263), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n381), .B1(new_n384), .B2(new_n372), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n341), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n265), .A2(new_n267), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n261), .A2(new_n341), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT79), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT80), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n390), .B1(new_n388), .B2(new_n389), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n388), .A2(new_n389), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT79), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT80), .B1(new_n397), .B2(new_n391), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n366), .B(new_n386), .C1(new_n395), .C2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT81), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n400), .A2(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(KEYINPUT17), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n393), .B1(new_n392), .B2(new_n394), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n397), .A2(KEYINPUT80), .A3(new_n391), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n404), .A2(new_n405), .B1(new_n385), .B2(new_n380), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n361), .A2(new_n362), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G169), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n361), .A2(G179), .A3(new_n362), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT18), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n406), .A2(new_n400), .A3(KEYINPUT17), .A4(new_n366), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n386), .B1(new_n395), .B2(new_n398), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n415), .A3(new_n410), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n403), .A2(new_n412), .A3(new_n413), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n333), .A2(G232), .ZN(new_n418));
  INV_X1    g0218(.A(G107), .ZN(new_n419));
  INV_X1    g0219(.A(G238), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n418), .B1(new_n419), .B2(new_n281), .C1(new_n420), .C2(new_n328), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n289), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n326), .B1(G244), .B2(new_n299), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n336), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n265), .A2(new_n267), .A3(G77), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT69), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n341), .B1(new_n427), .B2(new_n248), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n427), .B2(new_n248), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT15), .B(G87), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n251), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n431), .A2(new_n432), .B1(G20), .B2(G77), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n426), .B1(G77), .B2(new_n270), .C1(new_n434), .C2(new_n367), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n424), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n436), .B1(new_n364), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G179), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n424), .A2(new_n309), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(new_n435), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NOR4_X1   g0243(.A1(new_n325), .A2(new_n356), .A3(new_n417), .A4(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n324), .A2(KEYINPUT77), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G283), .ZN(new_n447));
  INV_X1    g0247(.A(G97), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n447), .B(new_n208), .C1(G33), .C2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT87), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(G20), .B1(new_n245), .B2(G97), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(KEYINPUT87), .A3(new_n447), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n208), .A2(G116), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n367), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n454), .A2(KEYINPUT20), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT20), .B1(new_n454), .B2(new_n456), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n256), .A2(G33), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n459), .B1(new_n265), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n261), .A2(G116), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n457), .A2(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT83), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n293), .A2(G1), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(KEYINPUT82), .C1(KEYINPUT5), .C2(new_n292), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n256), .B(G45), .C1(new_n292), .C2(KEYINPUT5), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT82), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n292), .A2(KEYINPUT5), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n288), .A2(G274), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n465), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n473), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(KEYINPUT83), .A3(new_n467), .A4(new_n470), .ZN(new_n476));
  INV_X1    g0276(.A(new_n472), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(new_n468), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(new_n289), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n474), .A2(new_n476), .B1(G270), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n281), .A2(G257), .A3(new_n284), .ZN(new_n481));
  INV_X1    g0281(.A(G303), .ZN(new_n482));
  INV_X1    g0282(.A(G264), .ZN(new_n483));
  OAI221_X1 g0283(.A(new_n481), .B1(new_n482), .B2(new_n281), .C1(new_n328), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n289), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n309), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT21), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n480), .A2(G179), .A3(new_n485), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n464), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n480), .A2(new_n485), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G200), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n480), .A2(G190), .A3(new_n485), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n464), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT88), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n490), .A2(new_n463), .A3(new_n495), .A4(G169), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT21), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n495), .B1(new_n486), .B2(new_n463), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT89), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n490), .A2(new_n463), .A3(G169), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT88), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT89), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(new_n497), .A4(new_n496), .ZN(new_n504));
  AOI211_X1 g0304(.A(new_n489), .B(new_n494), .C1(new_n500), .C2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT23), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n208), .B2(G107), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n419), .A2(KEYINPUT23), .A3(G20), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n432), .A2(G116), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n208), .B(G87), .C1(new_n276), .C2(new_n277), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n511), .A2(KEYINPUT22), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(KEYINPUT22), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT24), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT24), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n516), .B(new_n510), .C1(new_n512), .C2(new_n513), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n367), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n270), .A2(G107), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT25), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n519), .A2(KEYINPUT25), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n265), .A2(new_n460), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n521), .A2(new_n522), .B1(new_n419), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n281), .A2(G257), .A3(G1698), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n281), .A2(G250), .A3(new_n284), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G294), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n529), .A2(new_n289), .B1(new_n479), .B2(G264), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n474), .A2(new_n476), .ZN(new_n531));
  AOI21_X1  g0331(.A(G200), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT92), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n531), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(G190), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n525), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n281), .A2(G250), .A3(G1698), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n281), .A2(G244), .A3(new_n284), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT4), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n447), .B(new_n538), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT4), .B1(new_n333), .B2(G244), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n289), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n479), .A2(G257), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n531), .A3(new_n544), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n545), .A2(G179), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n419), .B1(new_n382), .B2(new_n383), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n419), .A2(KEYINPUT6), .A3(G97), .ZN(new_n548));
  XOR2_X1   g0348(.A(G97), .B(G107), .Z(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(KEYINPUT6), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G20), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n252), .B2(new_n248), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n246), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n270), .A2(G97), .ZN(new_n554));
  INV_X1    g0354(.A(new_n523), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n554), .B1(new_n555), .B2(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n545), .A2(new_n309), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n546), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  OR2_X1    g0359(.A1(new_n545), .A2(new_n336), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n545), .A2(G200), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n560), .A2(new_n553), .A3(new_n556), .A4(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n537), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT90), .ZN(new_n564));
  INV_X1    g0364(.A(new_n522), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n565), .A2(new_n520), .B1(G107), .B2(new_n555), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n515), .A2(new_n517), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n564), .B(new_n566), .C1(new_n567), .C2(new_n367), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT90), .B1(new_n518), .B2(new_n524), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n534), .A2(KEYINPUT91), .A3(G169), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n530), .A2(new_n531), .A3(G179), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT91), .B1(new_n534), .B2(G169), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n568), .B(new_n569), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT85), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n281), .A2(G238), .A3(new_n284), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT84), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT84), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n333), .A2(new_n578), .A3(G238), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n245), .A2(new_n459), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n373), .A2(new_n284), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(new_n582), .B2(G244), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n288), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n466), .A2(G250), .ZN(new_n585));
  INV_X1    g0385(.A(G274), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n466), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n288), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n575), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(G244), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n328), .A2(new_n591), .B1(new_n245), .B2(new_n459), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n579), .B2(new_n577), .ZN(new_n593));
  OAI211_X1 g0393(.A(KEYINPUT85), .B(new_n588), .C1(new_n593), .C2(new_n288), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n309), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n281), .A2(new_n208), .A3(G68), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT19), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n208), .B1(new_n283), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(G87), .B2(new_n203), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n598), .B1(new_n251), .B2(new_n448), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n246), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n261), .A2(new_n430), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT86), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(KEYINPUT86), .A3(new_n604), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n555), .A2(new_n431), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n590), .A2(new_n594), .A3(new_n439), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n596), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n579), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n578), .B1(new_n333), .B2(G238), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n583), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n289), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT85), .B1(new_n617), .B2(new_n588), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n584), .A2(new_n575), .A3(new_n589), .ZN(new_n619));
  OAI21_X1  g0419(.A(G200), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n607), .A2(new_n608), .B1(G87), .B2(new_n555), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n590), .A2(new_n594), .A3(G190), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n574), .A2(new_n613), .A3(new_n623), .ZN(new_n624));
  NOR4_X1   g0424(.A1(new_n446), .A2(new_n506), .A3(new_n563), .A4(new_n624), .ZN(G372));
  OAI21_X1  g0425(.A(new_n588), .B1(new_n593), .B2(new_n288), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n309), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n627), .B(KEYINPUT93), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n611), .A2(new_n612), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(G200), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n622), .A2(new_n621), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n633), .A2(new_n559), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n559), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n613), .A3(new_n623), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT26), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n630), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n489), .B1(new_n500), .B2(new_n504), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n572), .A2(new_n573), .B1(new_n518), .B2(new_n524), .ZN(new_n642));
  AOI211_X1 g0442(.A(new_n563), .B(new_n633), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n444), .A2(new_n445), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n323), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n320), .B1(new_n646), .B2(new_n442), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n403), .A2(new_n413), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n412), .A2(new_n416), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n353), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(new_n355), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n645), .A2(new_n653), .ZN(G369));
  NAND3_X1  g0454(.A1(new_n256), .A2(new_n208), .A3(G13), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n464), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT94), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n506), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n505), .A2(KEYINPUT94), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n664), .A2(new_n665), .B1(new_n641), .B2(new_n662), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n568), .A2(new_n569), .A3(new_n660), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT95), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n670), .A2(new_n537), .A3(new_n574), .A4(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n574), .B2(new_n661), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n641), .A2(new_n660), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n672), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n642), .A2(new_n660), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n674), .A2(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n212), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G1), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT96), .ZN(new_n687));
  OAI22_X1  g0487(.A1(new_n686), .A2(new_n687), .B1(new_n205), .B2(new_n684), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n687), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT97), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT28), .Z(new_n691));
  NOR2_X1   g0491(.A1(new_n633), .A2(new_n563), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n641), .A2(new_n574), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT99), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n634), .A2(new_n635), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n630), .B1(new_n638), .B2(KEYINPUT26), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n660), .B1(new_n695), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n644), .A2(new_n661), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n480), .A2(G179), .A3(new_n485), .ZN(new_n706));
  AND4_X1   g0506(.A1(new_n531), .A2(new_n543), .A3(new_n530), .A4(new_n544), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n705), .B1(new_n708), .B2(new_n595), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n490), .A2(new_n626), .A3(new_n439), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n545), .A2(new_n534), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT98), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT98), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n545), .A2(new_n713), .A3(new_n534), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n710), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n543), .A2(new_n530), .A3(new_n531), .A4(new_n544), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n488), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n590), .A4(new_n594), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n709), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT31), .B1(new_n719), .B2(new_n660), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n624), .A2(new_n563), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n505), .A2(new_n723), .A3(new_n661), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G330), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n704), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(KEYINPUT100), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(KEYINPUT100), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n691), .B1(new_n734), .B2(G1), .ZN(G364));
  INV_X1    g0535(.A(G13), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n256), .B1(new_n737), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n683), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n667), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n666), .A2(G330), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n666), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n207), .B1(G20), .B2(new_n309), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n208), .A2(G179), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G190), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G159), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT32), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n208), .A2(new_n439), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n336), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n756), .A2(G190), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n754), .B1(new_n758), .B2(new_n249), .C1(new_n263), .C2(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n336), .A2(G179), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n208), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G97), .ZN(new_n765));
  OR3_X1    g0565(.A1(new_n752), .A2(KEYINPUT32), .A3(new_n753), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G87), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n750), .A2(new_n336), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G107), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n765), .A2(new_n766), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n755), .A2(new_n751), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n755), .A2(G190), .A3(new_n364), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n281), .B1(new_n774), .B2(new_n252), .C1(new_n368), .C2(new_n775), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n761), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G294), .A2(new_n764), .B1(new_n757), .B2(G326), .ZN(new_n778));
  INV_X1    g0578(.A(new_n775), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G322), .ZN(new_n780));
  INV_X1    g0580(.A(new_n774), .ZN(new_n781));
  INV_X1    g0581(.A(new_n752), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G311), .A2(new_n781), .B1(new_n782), .B2(G329), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n759), .A2(new_n784), .B1(new_n771), .B2(G283), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n778), .A2(new_n780), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n373), .B1(new_n767), .B2(new_n482), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT102), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n749), .B1(new_n777), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n740), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n746), .A2(new_n749), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n682), .A2(new_n373), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n793), .A2(G355), .B1(new_n459), .B2(new_n682), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n239), .A2(new_n293), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n373), .A2(new_n212), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(new_n293), .B2(new_n206), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT101), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n794), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n791), .B1(new_n792), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n741), .A2(new_n743), .B1(new_n748), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  INV_X1    g0602(.A(KEYINPUT105), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n442), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n435), .A2(new_n660), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n440), .A2(KEYINPUT105), .A3(new_n435), .A4(new_n441), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n804), .A2(new_n438), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n442), .A2(new_n661), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n701), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n804), .A2(new_n806), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n438), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n661), .B(new_n814), .C1(new_n640), .C2(new_n643), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n740), .B1(new_n816), .B2(new_n729), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n729), .B2(new_n816), .ZN(new_n818));
  INV_X1    g0618(.A(new_n740), .ZN(new_n819));
  INV_X1    g0619(.A(new_n749), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n779), .A2(G143), .B1(new_n781), .B2(G159), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n758), .B2(new_n822), .C1(new_n342), .C2(new_n760), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT103), .B(KEYINPUT34), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n823), .B(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n825), .A2(KEYINPUT104), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(KEYINPUT104), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n771), .A2(G68), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n281), .C1(new_n829), .C2(new_n752), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n763), .A2(new_n368), .B1(new_n767), .B2(new_n249), .ZN(new_n831));
  OR4_X1    g0631(.A1(new_n826), .A2(new_n827), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G87), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n758), .A2(new_n482), .B1(new_n770), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(G107), .B2(new_n768), .ZN(new_n835));
  INV_X1    g0635(.A(G294), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n775), .A2(new_n836), .B1(new_n774), .B2(new_n459), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n281), .B(new_n837), .C1(G311), .C2(new_n782), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n759), .A2(G283), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n835), .A2(new_n765), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n820), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n749), .A2(new_n744), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n819), .B(new_n841), .C1(new_n252), .C2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n809), .B2(new_n745), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n818), .A2(new_n844), .ZN(G384));
  NOR2_X1   g0645(.A1(new_n737), .A2(new_n256), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n446), .A2(new_n726), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT112), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n810), .B1(new_n722), .B2(new_n724), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n310), .A2(KEYINPUT75), .A3(new_n275), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n313), .B1(new_n312), .B2(KEYINPUT14), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n318), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT76), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n317), .A2(new_n316), .A3(new_n318), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n273), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n273), .A2(new_n661), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n855), .A2(new_n646), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n856), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n320), .B2(new_n323), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n849), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT110), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n414), .A2(new_n410), .ZN(new_n864));
  INV_X1    g0664(.A(new_n658), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n414), .A2(new_n865), .ZN(new_n866));
  AND4_X1   g0666(.A1(new_n863), .A2(new_n864), .A3(new_n866), .A4(new_n399), .ZN(new_n867));
  INV_X1    g0667(.A(new_n372), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT7), .ZN(new_n869));
  OAI21_X1  g0669(.A(G68), .B1(new_n376), .B2(new_n869), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n373), .A2(new_n377), .A3(new_n208), .ZN(new_n871));
  OAI211_X1 g0671(.A(KEYINPUT16), .B(new_n868), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n246), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n379), .A2(KEYINPUT16), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n391), .B(new_n397), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n410), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n399), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT108), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT108), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n399), .A2(new_n879), .A3(new_n876), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT107), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n875), .A2(new_n881), .A3(new_n865), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n881), .B1(new_n875), .B2(new_n865), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n878), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n867), .B1(new_n885), .B2(KEYINPUT37), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n875), .A2(new_n865), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT107), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n875), .A2(new_n881), .A3(new_n865), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n417), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n862), .B1(new_n886), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n879), .B1(new_n399), .B2(new_n876), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n863), .B1(new_n895), .B2(new_n880), .ZN(new_n896));
  OAI211_X1 g0696(.A(KEYINPUT38), .B(new_n891), .C1(new_n896), .C2(new_n867), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n856), .B1(new_n855), .B2(new_n646), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n320), .A2(new_n323), .A3(new_n858), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT110), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n903), .A3(new_n849), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n861), .A2(new_n899), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT111), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT111), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n905), .A2(new_n909), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT109), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n648), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n650), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n648), .A2(new_n912), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n414), .B(new_n865), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n864), .A2(new_n866), .A3(new_n399), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT37), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT38), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n897), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT40), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n911), .B1(new_n860), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n848), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n848), .A2(new_n922), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n923), .A2(new_n924), .A3(new_n727), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n919), .B2(new_n920), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n898), .A2(KEYINPUT39), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n320), .A2(new_n660), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n812), .A2(new_n660), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n815), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(new_n899), .A3(new_n902), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n651), .A2(new_n658), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n933), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n704), .A2(new_n446), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n653), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n939), .B(new_n941), .Z(new_n942));
  AOI21_X1  g0742(.A(new_n846), .B1(new_n926), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n942), .B2(new_n926), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n945), .A2(G116), .A3(new_n209), .A4(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT36), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n369), .A2(new_n205), .A3(new_n252), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n949), .A2(KEYINPUT106), .B1(new_n249), .B2(G68), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(KEYINPUT106), .B2(new_n949), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(G1), .A3(new_n736), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n944), .A2(new_n948), .A3(new_n952), .ZN(G367));
  INV_X1    g0753(.A(new_n733), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(new_n731), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n637), .A2(new_n660), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n557), .A2(new_n660), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n562), .A2(new_n559), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(KEYINPUT113), .B(KEYINPUT44), .Z(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OR3_X1    g0761(.A1(new_n680), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n961), .B1(new_n680), .B2(new_n959), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n680), .A2(new_n959), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT45), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT45), .B1(new_n680), .B2(new_n959), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n962), .B(new_n963), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n674), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT115), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n966), .A2(new_n967), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n962), .A2(new_n963), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT115), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n674), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n674), .A2(KEYINPUT114), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n968), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n674), .A2(KEYINPUT114), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n970), .A2(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n678), .B1(new_n673), .B2(new_n675), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n667), .B(new_n979), .Z(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n955), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n683), .B(KEYINPUT41), .Z(new_n983));
  OAI21_X1  g0783(.A(new_n738), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n677), .A2(new_n959), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n985), .A2(KEYINPUT42), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n559), .B1(new_n958), .B2(new_n574), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n985), .A2(KEYINPUT42), .B1(new_n661), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n621), .A2(new_n661), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n633), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n628), .A2(new_n629), .A3(new_n989), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n986), .A2(new_n988), .B1(KEYINPUT43), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n969), .A2(new_n959), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n984), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n234), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n792), .B1(new_n212), .B2(new_n430), .C1(new_n999), .C2(new_n796), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n1000), .A2(new_n740), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n759), .A2(G294), .B1(new_n771), .B2(G97), .ZN(new_n1002));
  XOR2_X1   g0802(.A(KEYINPUT116), .B(G311), .Z(new_n1003));
  OAI221_X1 g0803(.A(new_n1002), .B1(new_n419), .B2(new_n763), .C1(new_n758), .C2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n779), .A2(G303), .B1(new_n782), .B2(G317), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n768), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT46), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n767), .B2(new_n459), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n281), .B1(new_n781), .B2(G283), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n768), .A2(G58), .B1(new_n771), .B2(G77), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n263), .B2(new_n763), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n759), .A2(G159), .B1(new_n757), .B2(G143), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n373), .B1(new_n779), .B2(G150), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G50), .A2(new_n781), .B1(new_n782), .B2(G137), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n1004), .A2(new_n1010), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT47), .Z(new_n1018));
  OAI221_X1 g0818(.A(new_n1001), .B1(new_n820), .B2(new_n1018), .C1(new_n992), .C2(new_n747), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n998), .A2(new_n1019), .ZN(G387));
  NAND2_X1  g0820(.A1(new_n734), .A2(new_n981), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n955), .A2(new_n980), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1021), .A2(new_n1022), .A3(new_n683), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n793), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n1024), .A2(new_n685), .B1(G107), .B2(new_n212), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n231), .A2(G45), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n685), .ZN(new_n1027));
  AOI211_X1 g0827(.A(G45), .B(new_n1027), .C1(G68), .C2(G77), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n341), .A2(G50), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT50), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n796), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1025), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n792), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n740), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n774), .A2(new_n263), .B1(new_n752), .B2(new_n342), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n373), .B(new_n1035), .C1(G50), .C2(new_n779), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n768), .A2(G77), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n763), .A2(new_n430), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n387), .B2(new_n759), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n757), .A2(G159), .B1(new_n771), .B2(G97), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n779), .A2(G317), .B1(new_n781), .B2(G303), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n757), .A2(G322), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n760), .C2(new_n1003), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(G283), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n763), .A2(new_n1047), .B1(new_n767), .B2(new_n836), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1046), .A2(KEYINPUT49), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n281), .B1(new_n782), .B2(G326), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n459), .C2(new_n770), .ZN(new_n1052));
  AOI21_X1  g0852(.A(KEYINPUT49), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1041), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1034), .B1(new_n1054), .B2(new_n749), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n673), .B2(new_n747), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT117), .Z(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n981), .B2(new_n739), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1023), .A2(new_n1058), .ZN(G393));
  OAI221_X1 g0859(.A(new_n792), .B1(new_n448), .B2(new_n212), .C1(new_n243), .C2(new_n796), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n740), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n758), .A2(new_n342), .B1(new_n753), .B2(new_n775), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT51), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n763), .A2(new_n252), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n387), .B2(new_n781), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(new_n249), .C2(new_n760), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n373), .B1(new_n782), .B2(G143), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n263), .B2(new_n767), .C1(new_n833), .C2(new_n770), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT118), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G317), .A2(new_n757), .B1(new_n779), .B2(G311), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT52), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n772), .B1(new_n760), .B2(new_n482), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n281), .B1(new_n782), .B2(G322), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n836), .B2(new_n774), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n763), .A2(new_n459), .B1(new_n767), .B2(new_n1047), .ZN(new_n1075));
  OR3_X1    g0875(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1066), .A2(new_n1069), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1061), .B1(new_n1077), .B2(new_n749), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n959), .B2(new_n747), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n970), .A2(new_n974), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n968), .A2(new_n969), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1079), .B1(new_n1082), .B2(new_n738), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n955), .A2(new_n980), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n684), .B1(new_n1084), .B2(new_n978), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1021), .A2(new_n1082), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(G390));
  NAND3_X1  g0888(.A1(new_n444), .A2(new_n445), .A3(new_n728), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n940), .A2(new_n653), .A3(new_n1089), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n849), .A2(G330), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n902), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1093), .A2(KEYINPUT119), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n902), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n729), .A2(KEYINPUT120), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT120), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n809), .B1(new_n728), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1095), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n934), .B1(new_n699), .B2(new_n814), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1093), .A2(KEYINPUT119), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1094), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1091), .A2(new_n902), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n936), .B1(new_n1093), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1090), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n932), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n919), .B2(new_n920), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n1100), .B2(new_n1095), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n936), .A2(new_n902), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1112), .A2(new_n1107), .B1(new_n928), .B2(new_n929), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1093), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1113), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1115), .A2(new_n1110), .A3(new_n1094), .A4(new_n1101), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1106), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1090), .A2(new_n1114), .A3(new_n1116), .A4(new_n1105), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1118), .A2(new_n683), .A3(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n739), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n760), .A2(new_n419), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1064), .B(new_n1123), .C1(G283), .C2(new_n757), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n774), .A2(new_n448), .B1(new_n752), .B2(new_n836), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n281), .B(new_n1125), .C1(G116), .C2(new_n779), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1124), .A2(new_n769), .A3(new_n828), .A4(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n775), .A2(new_n829), .B1(new_n774), .B2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n373), .B(new_n1129), .C1(G125), .C2(new_n782), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n767), .A2(new_n342), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n759), .A2(G137), .B1(new_n771), .B2(G50), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G159), .A2(new_n764), .B1(new_n757), .B2(G128), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n820), .B1(new_n1127), .B2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n819), .B(new_n1136), .C1(new_n341), .C2(new_n842), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n931), .B2(new_n745), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1120), .A2(new_n1122), .A3(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(KEYINPUT121), .ZN(new_n1140));
  OAI21_X1  g0940(.A(G330), .B1(new_n921), .B2(new_n860), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n898), .B1(new_n860), .B2(KEYINPUT110), .ZN(new_n1143));
  AOI211_X1 g0943(.A(KEYINPUT111), .B(KEYINPUT40), .C1(new_n1143), .C2(new_n904), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n909), .B1(new_n905), .B2(new_n906), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1142), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n356), .A2(new_n349), .A3(new_n865), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n349), .A2(new_n865), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n353), .A2(new_n355), .A3(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1147), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1146), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1153), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n1142), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1154), .A2(new_n939), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n939), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1140), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n939), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1155), .B1(new_n911), .B2(new_n1142), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1141), .B(new_n1153), .C1(new_n908), .C2(new_n910), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1154), .A2(new_n939), .A3(new_n1156), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(KEYINPUT121), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1159), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n940), .A2(new_n653), .A3(new_n1089), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1121), .B2(new_n1105), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT57), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1106), .A2(new_n1117), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1171), .B(KEYINPUT57), .C1(new_n1167), .C2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n683), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1153), .A2(new_n744), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n758), .A2(new_n459), .B1(new_n770), .B2(new_n368), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G97), .B2(new_n759), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n373), .A2(new_n292), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G283), .B2(new_n782), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n779), .A2(G107), .B1(new_n781), .B2(new_n431), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n764), .A2(G68), .B1(new_n768), .B2(G77), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT58), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1179), .B(new_n249), .C1(G33), .C2(G41), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n757), .A2(G125), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n760), .B2(new_n829), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n779), .A2(G128), .B1(new_n781), .B2(G137), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n767), .B2(new_n1128), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1189), .B(new_n1191), .C1(G150), .C2(new_n764), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n771), .A2(G159), .ZN(new_n1195));
  AOI211_X1 g0995(.A(G33), .B(G41), .C1(new_n782), .C2(G124), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1187), .B1(new_n1184), .B2(new_n1183), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n749), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n819), .B1(new_n249), .B2(new_n842), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1176), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1166), .B2(new_n739), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1175), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(G375));
  INV_X1    g1007(.A(new_n1105), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(new_n738), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n819), .B1(new_n263), .B2(new_n842), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n760), .A2(new_n459), .B1(new_n758), .B2(new_n836), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G97), .B2(new_n768), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n281), .B1(new_n782), .B2(G303), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n419), .B2(new_n774), .C1(new_n1047), .C2(new_n775), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1038), .B(new_n1214), .C1(G77), .C2(new_n771), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n757), .A2(G132), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n822), .B2(new_n775), .C1(new_n760), .C2(new_n1128), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT123), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n368), .A2(new_n770), .B1(new_n767), .B2(new_n753), .ZN(new_n1219));
  INV_X1    g1019(.A(G128), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n281), .B1(new_n752), .B2(new_n1220), .C1(new_n342), .C2(new_n774), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G50), .C2(new_n764), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1212), .A2(new_n1215), .B1(new_n1218), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1210), .B1(new_n1223), .B2(new_n820), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1095), .A2(KEYINPUT122), .A3(new_n744), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT122), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n902), .B2(new_n745), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1224), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1209), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1208), .A2(new_n1167), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n983), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1231), .A3(new_n1106), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(G381));
  INV_X1    g1033(.A(G384), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1087), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1023), .A2(new_n801), .A3(new_n1058), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(new_n1235), .A2(G378), .A3(G381), .A4(new_n1236), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1206), .A2(new_n1237), .A3(new_n998), .A4(new_n1019), .ZN(G407));
  INV_X1    g1038(.A(G378), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n659), .A2(G213), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1206), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(G407), .A2(G213), .A3(new_n1242), .ZN(G409));
  INV_X1    g1043(.A(KEYINPUT127), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1236), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n801), .B1(new_n1023), .B2(new_n1058), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n998), .A2(new_n1019), .A3(new_n1087), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1087), .B1(new_n998), .B2(new_n1019), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1244), .B(new_n1247), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(G390), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT127), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1246), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n1244), .A3(new_n1236), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .A4(new_n1248), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1251), .A2(new_n1252), .A3(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G378), .B(new_n1204), .C1(new_n1170), .C2(new_n1174), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n983), .B(new_n1168), .C1(new_n1159), .C2(new_n1165), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1171), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1202), .B1(new_n1261), .B2(new_n738), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1239), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1241), .B1(new_n1259), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1106), .A2(new_n683), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT125), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1230), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT60), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1230), .A2(new_n1266), .A3(KEYINPUT60), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1265), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT126), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1229), .B1(G384), .B2(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1234), .A2(KEYINPUT126), .ZN(new_n1274));
  OR3_X1    g1074(.A1(new_n1271), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1258), .B1(new_n1264), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1259), .A2(new_n1263), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT124), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT124), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1259), .A2(new_n1263), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1240), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1241), .A2(G2897), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1277), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1275), .A2(G2897), .A3(new_n1241), .A4(new_n1276), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1286), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1283), .A2(new_n1240), .A3(new_n1277), .A4(new_n1285), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1279), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1281), .A2(new_n1290), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1252), .B1(new_n1294), .B2(new_n1264), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT62), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1291), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1264), .A2(KEYINPUT62), .A3(new_n1277), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1295), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1251), .A2(new_n1257), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1293), .B1(new_n1299), .B2(new_n1300), .ZN(G405));
  NOR2_X1   g1101(.A1(new_n1206), .A2(G378), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1259), .ZN(new_n1303));
  OR3_X1    g1103(.A1(new_n1302), .A2(new_n1278), .A3(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1278), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1304), .A2(new_n1300), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1300), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(G402));
endmodule


