//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n639, new_n640, new_n641, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n462), .A2(G2104), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n467));
  OR2_X1    g042(.A1(new_n467), .A2(new_n462), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n461), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n464), .A2(G136), .ZN(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G162));
  AND2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  OAI211_X1 g055(.A(G126), .B(G2105), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n479), .B2(new_n480), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n484), .B(new_n487), .C1(new_n480), .C2(new_n479), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n482), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  OAI21_X1  g065(.A(G2105), .B1(KEYINPUT67), .B2(G114), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT67), .A2(G114), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n494), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(KEYINPUT68), .C1(new_n492), .C2(new_n491), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n489), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT69), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT69), .A2(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT6), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT69), .B(G651), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n507), .A2(G50), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n516));
  INV_X1    g091(.A(new_n511), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  OR2_X1    g093(.A1(KEYINPUT69), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT69), .A2(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n517), .B(G88), .C1(new_n521), .C2(new_n505), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n515), .A2(new_n516), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g098(.A(G50), .B(G543), .C1(new_n521), .C2(new_n505), .ZN(new_n524));
  OR2_X1    g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n512), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n508), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n514), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n522), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT70), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n523), .A2(new_n531), .ZN(G166));
  AOI21_X1  g107(.A(new_n505), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n511), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT71), .B(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n517), .A2(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n507), .A2(G51), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  NAND2_X1  g120(.A1(new_n534), .A2(G90), .ZN(new_n546));
  XOR2_X1   g121(.A(KEYINPUT72), .B(G52), .Z(new_n547));
  NAND2_X1  g122(.A1(new_n507), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G64), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n511), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(new_n514), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n546), .A2(new_n548), .A3(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n511), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(new_n514), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT74), .B(G81), .Z(new_n559));
  NAND2_X1  g134(.A1(new_n534), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT73), .B(G43), .Z(new_n562));
  NAND2_X1  g137(.A1(new_n507), .A2(new_n562), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n561), .B1(new_n560), .B2(new_n563), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n558), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  OAI211_X1 g147(.A(G53), .B(G543), .C1(new_n521), .C2(new_n505), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n507), .B2(G53), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT76), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n507), .A2(new_n575), .A3(G53), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(new_n533), .B2(new_n511), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n517), .B(KEYINPUT77), .C1(new_n521), .C2(new_n505), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n584), .A2(G91), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G78), .A2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(KEYINPUT78), .B(G65), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n511), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n582), .A2(new_n591), .ZN(G299));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n516), .B1(new_n515), .B2(new_n522), .ZN(new_n594));
  AND4_X1   g169(.A1(new_n516), .A2(new_n522), .A3(new_n524), .A4(new_n529), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n523), .A2(new_n531), .A3(KEYINPUT79), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(G303));
  NAND3_X1  g173(.A1(new_n584), .A2(G87), .A3(new_n585), .ZN(new_n599));
  INV_X1    g174(.A(G651), .ZN(new_n600));
  INV_X1    g175(.A(G74), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n511), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n507), .B2(G49), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(G288));
  NAND3_X1  g179(.A1(new_n584), .A2(G86), .A3(new_n585), .ZN(new_n605));
  INV_X1    g180(.A(G61), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n525), .B2(new_n526), .ZN(new_n607));
  NAND2_X1  g182(.A1(G73), .A2(G543), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT80), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n610), .A2(G73), .A3(G543), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g187(.A(KEYINPUT81), .B(new_n514), .C1(new_n607), .C2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n514), .B1(new_n607), .B2(new_n612), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n614), .A2(new_n615), .B1(new_n507), .B2(G48), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n605), .A2(new_n613), .A3(new_n616), .ZN(G305));
  NAND2_X1  g192(.A1(G72), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G60), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n511), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(new_n514), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT83), .B(G47), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n534), .A2(G85), .B1(new_n507), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n625), .ZN(G290));
  NAND2_X1  g201(.A1(G301), .A2(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n507), .A2(G54), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n600), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g205(.A1(new_n584), .A2(new_n585), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G92), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n631), .A2(KEYINPUT10), .A3(G92), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n627), .B1(new_n636), .B2(G868), .ZN(G284));
  OAI21_X1  g212(.A(new_n627), .B1(new_n636), .B2(G868), .ZN(G321));
  NAND2_X1  g213(.A1(G286), .A2(G868), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT84), .ZN(new_n640));
  INV_X1    g215(.A(G299), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(G868), .B2(new_n641), .ZN(G297));
  OAI21_X1  g217(.A(new_n640), .B1(G868), .B2(new_n641), .ZN(G280));
  INV_X1    g218(.A(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n636), .B1(new_n644), .B2(G860), .ZN(G148));
  NAND2_X1  g220(.A1(new_n634), .A2(new_n635), .ZN(new_n646));
  INV_X1    g221(.A(new_n630), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n648), .A2(G559), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT85), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  MUX2_X1   g226(.A(new_n566), .B(new_n651), .S(G868), .Z(G323));
  XNOR2_X1  g227(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g228(.A1(new_n461), .A2(new_n465), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT12), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT13), .ZN(new_n656));
  INV_X1    g231(.A(G2100), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n464), .A2(G135), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n472), .A2(G123), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n462), .A2(G111), .ZN(new_n662));
  OAI21_X1  g237(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n660), .B(new_n661), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(G2096), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n658), .A2(new_n659), .A3(new_n666), .ZN(G156));
  XNOR2_X1  g242(.A(G2427), .B(G2438), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2430), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT15), .B(G2435), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(KEYINPUT14), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2451), .B(G2454), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT16), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2443), .B(G2446), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1341), .B(G1348), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  OAI21_X1  g256(.A(G14), .B1(new_n678), .B2(new_n679), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(G401));
  INV_X1    g258(.A(KEYINPUT18), .ZN(new_n684));
  XOR2_X1   g259(.A(G2084), .B(G2090), .Z(new_n685));
  XNOR2_X1  g260(.A(G2067), .B(G2678), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(KEYINPUT17), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n685), .A2(new_n686), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT87), .B(G2100), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G2072), .B(G2078), .Z(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n687), .B2(KEYINPUT18), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(new_n665), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n692), .B(new_n695), .ZN(G227));
  XOR2_X1   g271(.A(G1971), .B(G1976), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT19), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1956), .B(G2474), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1961), .B(G1966), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(new_n701), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT20), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n698), .A2(new_n702), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(KEYINPUT88), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(KEYINPUT88), .ZN(new_n708));
  AOI211_X1 g283(.A(new_n703), .B(new_n705), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1991), .B(G1996), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(G1981), .B(G1986), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(G229));
  MUX2_X1   g291(.A(G24), .B(G290), .S(G16), .Z(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G1986), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n472), .A2(G119), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n464), .A2(G131), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n462), .A2(G107), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n719), .B(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G25), .B(new_n723), .S(G29), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  MUX2_X1   g301(.A(G6), .B(G305), .S(G16), .Z(new_n727));
  XOR2_X1   g302(.A(KEYINPUT32), .B(G1981), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G16), .A2(G22), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G166), .B2(G16), .ZN(new_n731));
  INV_X1    g306(.A(G1971), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G16), .A2(G23), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT89), .Z(new_n735));
  INV_X1    g310(.A(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(G288), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT33), .B(G1976), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT90), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n737), .B(new_n739), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n729), .A2(new_n733), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n718), .B(new_n726), .C1(new_n742), .C2(KEYINPUT34), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT91), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(KEYINPUT34), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT36), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT31), .B(G11), .Z(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G28), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(KEYINPUT93), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n750), .B2(G28), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(KEYINPUT93), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n748), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G168), .A2(new_n736), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n736), .B2(G21), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT92), .B(G1966), .Z(new_n758));
  OAI221_X1 g333(.A(new_n755), .B1(new_n749), .B2(new_n664), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n736), .A2(G5), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G171), .B2(new_n736), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT94), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G1961), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n760), .A2(KEYINPUT95), .A3(new_n764), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT25), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n461), .A2(G127), .ZN(new_n774));
  NAND2_X1  g349(.A1(G115), .A2(G2104), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n462), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n773), .B(new_n776), .C1(G139), .C2(new_n464), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(new_n749), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n749), .B2(G33), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(G2072), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT24), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n782), .A2(G34), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n749), .B1(new_n782), .B2(G34), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n469), .A2(new_n749), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G2084), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n780), .A2(G2072), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n781), .A2(new_n787), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n763), .A2(G1961), .ZN(new_n791));
  NAND2_X1  g366(.A1(G164), .A2(G29), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G27), .B2(G29), .ZN(new_n793));
  INV_X1    g368(.A(G2078), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n749), .A2(G32), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n464), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n472), .A2(G129), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT26), .Z(new_n800));
  AND3_X1   g375(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n796), .B1(new_n801), .B2(new_n749), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT27), .B(G1996), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n793), .A2(new_n794), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n790), .A2(new_n791), .A3(new_n795), .A4(new_n806), .ZN(new_n807));
  AND3_X1   g382(.A1(new_n767), .A2(new_n768), .A3(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT96), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT96), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n749), .A2(G35), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G162), .B2(new_n749), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT29), .B(G2090), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n749), .A2(G26), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT28), .Z(new_n816));
  OR2_X1    g391(.A1(G104), .A2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n818));
  INV_X1    g393(.A(G140), .ZN(new_n819));
  INV_X1    g394(.A(G128), .ZN(new_n820));
  OAI221_X1 g395(.A(new_n818), .B1(new_n463), .B2(new_n819), .C1(new_n820), .C2(new_n471), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n816), .B1(new_n821), .B2(G29), .ZN(new_n822));
  INV_X1    g397(.A(G2067), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n567), .A2(G16), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G16), .B2(G19), .ZN(new_n826));
  INV_X1    g401(.A(G1341), .ZN(new_n827));
  AOI211_X1 g402(.A(new_n814), .B(new_n824), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n827), .B2(new_n826), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n736), .A2(G4), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n636), .B2(new_n736), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G1348), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n736), .A2(G20), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT23), .Z(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G299), .B2(G16), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT97), .B(G1956), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n829), .A2(new_n832), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n809), .A2(new_n810), .A3(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n747), .A2(new_n839), .ZN(G311));
  NAND2_X1  g415(.A1(new_n747), .A2(new_n839), .ZN(G150));
  NAND2_X1  g416(.A1(new_n636), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n534), .A2(G93), .ZN(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT98), .B(G55), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n507), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(G80), .A2(G543), .ZN(new_n847));
  INV_X1    g422(.A(G67), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n511), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(new_n514), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n844), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n566), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n851), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n853), .B(new_n558), .C1(new_n564), .C2(new_n565), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n843), .B(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n858), .A2(new_n859), .A3(G860), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n851), .A2(G860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT37), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n860), .A2(new_n862), .ZN(G145));
  XNOR2_X1  g438(.A(new_n821), .B(KEYINPUT99), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n499), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n801), .ZN(new_n866));
  OR3_X1    g441(.A1(new_n866), .A2(KEYINPUT101), .A3(new_n777), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT101), .B1(new_n866), .B2(new_n777), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n777), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n866), .A2(KEYINPUT100), .A3(new_n777), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n723), .B(new_n655), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n472), .A2(G130), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n464), .A2(G142), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n878), .A2(new_n462), .A3(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n462), .B2(G118), .ZN(new_n880));
  OR2_X1    g455(.A1(G106), .A2(G2105), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(G2104), .A3(new_n881), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n876), .B(new_n877), .C1(new_n879), .C2(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n875), .B(new_n883), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT103), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n869), .A2(new_n874), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n469), .B(new_n664), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n477), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n869), .A2(new_n874), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(new_n890), .B2(new_n884), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n885), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n892), .B2(new_n886), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n650), .A2(new_n856), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n650), .A2(new_n856), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n636), .A2(new_n641), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n636), .A2(new_n641), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n902), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n905), .B2(new_n906), .ZN(new_n910));
  INV_X1    g485(.A(new_n906), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(KEYINPUT41), .A3(new_n904), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n900), .A2(new_n901), .A3(new_n910), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n903), .B1(new_n902), .B2(new_n907), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n899), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n599), .A2(new_n603), .ZN(new_n917));
  XNOR2_X1  g492(.A(G290), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT105), .ZN(new_n919));
  XOR2_X1   g494(.A(G166), .B(G305), .Z(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n918), .A2(KEYINPUT105), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n918), .A2(KEYINPUT105), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n921), .B1(new_n924), .B2(new_n920), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(new_n897), .B2(new_n898), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n902), .A2(new_n907), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT104), .ZN(new_n929));
  INV_X1    g504(.A(new_n899), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n929), .A2(new_n930), .A3(new_n913), .A4(new_n908), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n916), .A2(new_n927), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n927), .B1(new_n916), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(G868), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n853), .A2(G868), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(G295));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n935), .ZN(G331));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n939));
  OAI21_X1  g514(.A(G171), .B1(G286), .B2(KEYINPUT107), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(G286), .A2(KEYINPUT107), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n566), .A2(new_n851), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(new_n854), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n854), .A3(new_n942), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n943), .A2(new_n854), .A3(new_n942), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n948), .A2(new_n944), .A3(new_n940), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n910), .B(new_n912), .C1(new_n947), .C2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(new_n941), .A3(new_n946), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n940), .B1(new_n948), .B2(new_n944), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n907), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n939), .B1(new_n954), .B2(new_n926), .ZN(new_n955));
  AOI211_X1 g530(.A(KEYINPUT109), .B(new_n925), .C1(new_n950), .C2(new_n953), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(KEYINPUT108), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n953), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n925), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n894), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n938), .B1(new_n962), .B2(KEYINPUT43), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n959), .B1(new_n950), .B2(new_n953), .ZN(new_n964));
  INV_X1    g539(.A(new_n960), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n926), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n961), .A2(new_n894), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(KEYINPUT43), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n957), .A2(new_n970), .A3(new_n894), .A4(new_n961), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT110), .B1(new_n972), .B2(new_n938), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n974), .B(KEYINPUT44), .C1(new_n969), .C2(new_n971), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n968), .B1(new_n973), .B2(new_n975), .ZN(G397));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n495), .A2(new_n497), .ZN(new_n978));
  INV_X1    g553(.A(new_n488), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n487), .B1(new_n461), .B2(new_n484), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n481), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT45), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n983), .B2(new_n982), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT112), .B(G40), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n466), .A2(new_n468), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n801), .B(G1996), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n821), .B(new_n823), .ZN(new_n991));
  INV_X1    g566(.A(new_n725), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n723), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n723), .A2(new_n992), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n990), .A2(new_n991), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(G290), .B(G1986), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n989), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n998));
  INV_X1    g573(.A(G8), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n982), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n489), .B2(new_n498), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT113), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n988), .B1(new_n982), .B2(KEYINPUT50), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT117), .B(G2084), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT45), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(new_n988), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT113), .B1(new_n499), .B2(new_n977), .ZN(new_n1014));
  AOI211_X1 g589(.A(new_n1000), .B(G1384), .C1(new_n489), .C2(new_n498), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n988), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(KEYINPUT116), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1011), .A2(new_n1012), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1008), .B1(new_n1019), .B2(new_n758), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n999), .B1(new_n1020), .B2(G168), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1012), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT116), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n758), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1008), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G286), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n998), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  AOI211_X1 g603(.A(KEYINPUT51), .B(new_n999), .C1(new_n1020), .C2(G168), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT62), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1024), .A2(G168), .A3(new_n1025), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G8), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1020), .A2(G168), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT51), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT62), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1021), .A2(new_n998), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT50), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1038));
  INV_X1    g613(.A(G2090), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n988), .B1(new_n1003), .B2(new_n1002), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n982), .A2(new_n1013), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(new_n1017), .A3(new_n1012), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n732), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n999), .B1(KEYINPUT114), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n596), .A2(new_n597), .A3(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(KEYINPUT114), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1049), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n596), .A2(new_n597), .A3(new_n1047), .A4(new_n1051), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1045), .A2(G8), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1001), .A2(new_n1017), .A3(new_n1004), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n917), .A2(G1976), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(G8), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT52), .ZN(new_n1057));
  INV_X1    g632(.A(G1976), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT52), .B1(G288), .B2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1054), .A2(G8), .A3(new_n1055), .A4(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1981), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n605), .A2(new_n1061), .A3(new_n616), .A4(new_n613), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n614), .A2(new_n615), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n507), .A2(G48), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n517), .B(G86), .C1(new_n521), .C2(new_n505), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1063), .A2(new_n1064), .A3(new_n613), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G1981), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT49), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1062), .A2(new_n1067), .A3(KEYINPUT49), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(G8), .A3(new_n1054), .A4(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1057), .A2(new_n1060), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1053), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1005), .A2(new_n1039), .A3(new_n1006), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n999), .B1(new_n1075), .B2(new_n1044), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1050), .A2(new_n1077), .A3(new_n1052), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n1043), .B2(G2078), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1083), .B(KEYINPUT125), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1082), .A2(G2078), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1011), .A2(new_n1012), .A3(new_n1085), .A4(new_n1018), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1088));
  INV_X1    g663(.A(G1961), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1086), .A2(new_n1087), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1087), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1084), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1081), .A2(G171), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1030), .A2(new_n1037), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n1096));
  NAND2_X1  g671(.A1(G168), .A2(G8), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1076), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1073), .A2(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1080), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1098), .A2(new_n1074), .A3(new_n1080), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1098), .A2(new_n1104), .B1(new_n1105), .B2(new_n1102), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1072), .A2(new_n1058), .A3(new_n917), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1062), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1054), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(new_n999), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1080), .B2(new_n1073), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1096), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1112), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1105), .A2(new_n1102), .ZN(new_n1115));
  AND4_X1   g690(.A1(new_n1080), .A2(new_n1098), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1116));
  OAI211_X1 g691(.A(KEYINPUT118), .B(new_n1114), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1095), .A2(new_n1113), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1956), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1002), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1040), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n578), .A2(new_n579), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(new_n586), .A3(new_n590), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n582), .A2(KEYINPUT57), .A3(new_n591), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1124), .A2(KEYINPUT119), .A3(new_n1125), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1042), .A2(new_n1017), .A3(new_n1012), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT56), .B(G2072), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1122), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(G1348), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1054), .A2(G2067), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1138), .A2(new_n648), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1131), .B1(new_n1122), .B2(new_n1134), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1135), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1122), .A2(new_n1134), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1131), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1135), .A2(KEYINPUT123), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1122), .A2(new_n1131), .A3(new_n1134), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1138), .A2(KEYINPUT60), .A3(new_n648), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n1151));
  INV_X1    g726(.A(G1996), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT58), .B(G1341), .Z(new_n1153));
  AOI22_X1  g728(.A1(new_n1132), .A2(new_n1152), .B1(new_n1054), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1151), .B1(new_n1154), .B2(new_n566), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1054), .A2(new_n1153), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1042), .A2(new_n1152), .A3(new_n1012), .A4(new_n1017), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1158), .A2(KEYINPUT121), .A3(new_n567), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1155), .A2(KEYINPUT120), .A3(KEYINPUT59), .A4(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1149), .A2(new_n1150), .A3(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n1162));
  AND3_X1   g737(.A1(new_n1122), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1163), .B2(new_n1140), .ZN(new_n1164));
  NAND2_X1  g739(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT121), .B1(new_n1158), .B2(new_n567), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n1151), .B(new_n566), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1137), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1088), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1169), .B(KEYINPUT60), .C1(new_n1170), .C2(G1348), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT60), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n636), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1164), .A2(new_n1168), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1141), .B1(new_n1161), .B2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1084), .B(G301), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1177));
  AND3_X1   g752(.A1(G160), .A2(G40), .A3(new_n1085), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n985), .A2(new_n1012), .A3(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1084), .A2(new_n1090), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(G171), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1177), .A2(new_n1181), .A3(KEYINPUT54), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1176), .A2(new_n1182), .A3(new_n1081), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1093), .A2(G171), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1084), .A2(G301), .A3(new_n1090), .A4(new_n1179), .ZN(new_n1185));
  AOI21_X1  g760(.A(KEYINPUT54), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1183), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n997), .B1(new_n1118), .B2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(G290), .A2(G1986), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n989), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1194));
  AOI211_X1 g769(.A(new_n1193), .B(new_n1194), .C1(new_n989), .C2(new_n995), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n991), .A2(new_n801), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n989), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT46), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1198), .B1(new_n989), .B2(new_n1152), .ZN(new_n1199));
  NOR4_X1   g774(.A1(new_n985), .A2(KEYINPUT46), .A3(G1996), .A4(new_n988), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1197), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT47), .Z(new_n1202));
  NAND2_X1  g777(.A1(new_n990), .A2(new_n991), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1203), .A2(new_n994), .B1(G2067), .B2(new_n821), .ZN(new_n1204));
  AOI211_X1 g779(.A(new_n1195), .B(new_n1202), .C1(new_n989), .C2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1189), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1189), .A2(KEYINPUT127), .A3(new_n1205), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g785(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1212));
  NAND3_X1  g786(.A1(new_n1212), .A2(new_n895), .A3(new_n972), .ZN(G225));
  INV_X1    g787(.A(G225), .ZN(G308));
endmodule


