//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G211gat), .A2(G218gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n205), .A2(KEYINPUT70), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT70), .B1(new_n205), .B2(new_n206), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n203), .B1(new_n210), .B2(KEYINPUT71), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(KEYINPUT71), .A3(new_n203), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT25), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT23), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G169gat), .B2(G176gat), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(G190gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n225), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n226), .A2(new_n229), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n216), .B1(new_n222), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n227), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(new_n226), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n235), .B2(new_n226), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n222), .A2(new_n216), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n233), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n217), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT26), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n219), .A2(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(KEYINPUT27), .B(G183gat), .Z(new_n243));
  INV_X1    g042(.A(KEYINPUT28), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n243), .A2(new_n244), .A3(G190gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G183gat), .ZN(new_n247));
  AOI21_X1  g046(.A(G190gat), .B1(new_n247), .B2(KEYINPUT27), .ZN(new_n248));
  OR3_X1    g047(.A1(new_n224), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT28), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI221_X1 g049(.A(new_n240), .B1(new_n217), .B2(new_n242), .C1(new_n245), .C2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT29), .B1(new_n239), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G226gat), .ZN(new_n253));
  INV_X1    g052(.A(G233gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n251), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n257), .A2(new_n255), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n215), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n255), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n260), .B(new_n214), .C1(new_n255), .C2(new_n252), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G8gat), .B(G36gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT72), .ZN(new_n264));
  XNOR2_X1  g063(.A(G64gat), .B(G92gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n259), .A2(new_n261), .A3(new_n266), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(KEYINPUT30), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n262), .A2(new_n271), .A3(new_n267), .ZN(new_n272));
  XOR2_X1   g071(.A(G141gat), .B(G148gat), .Z(new_n273));
  INV_X1    g072(.A(G155gat), .ZN(new_n274));
  INV_X1    g073(.A(G162gat), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT2), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G155gat), .B(G162gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n273), .A2(new_n278), .A3(new_n276), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G113gat), .B(G120gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n287));
  XNOR2_X1  g086(.A(G127gat), .B(G134gat), .ZN(new_n288));
  INV_X1    g087(.A(G120gat), .ZN(new_n289));
  OR3_X1    g088(.A1(new_n289), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n286), .A2(new_n287), .A3(new_n288), .A4(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n288), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(KEYINPUT1), .B2(new_n285), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT3), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n284), .B(new_n294), .C1(new_n295), .C2(new_n282), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n297));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT4), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n281), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(new_n294), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n301), .A2(new_n294), .A3(new_n300), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT74), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n294), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n282), .A2(new_n306), .A3(KEYINPUT4), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n302), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n296), .A2(new_n302), .A3(new_n307), .A4(new_n298), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n301), .B(new_n294), .ZN(new_n312));
  INV_X1    g111(.A(new_n298), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n297), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n299), .A2(new_n310), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G1gat), .B(G29gat), .Z(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT0), .ZN(new_n317));
  XNOR2_X1  g116(.A(G57gat), .B(G85gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n319), .B(KEYINPUT79), .Z(new_n320));
  OR2_X1    g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n270), .A2(new_n272), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT82), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(KEYINPUT40), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n309), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n308), .B1(new_n307), .B2(new_n302), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n296), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n313), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n329), .B(KEYINPUT39), .C1(new_n313), .C2(new_n312), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT80), .B(KEYINPUT39), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(new_n313), .A3(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n332), .A2(KEYINPUT81), .A3(new_n320), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT81), .B1(new_n332), .B2(new_n320), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n325), .B(new_n330), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n322), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(new_n320), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n332), .A2(KEYINPUT81), .A3(new_n320), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n325), .B1(new_n341), .B2(new_n330), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n315), .A2(new_n319), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n344), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n346), .B1(new_n315), .B2(new_n319), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n345), .B1(new_n347), .B2(new_n321), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT37), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n259), .A2(new_n349), .A3(new_n261), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n349), .B1(new_n259), .B2(new_n261), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n266), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT38), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT38), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n354), .B(new_n266), .C1(new_n350), .C2(new_n351), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n348), .A2(new_n268), .A3(new_n353), .A4(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G78gat), .B(G106gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT31), .B(G50gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT77), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n212), .A2(new_n361), .A3(new_n213), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n282), .B1(new_n362), .B2(new_n295), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n284), .A2(new_n361), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n364), .A2(new_n214), .ZN(new_n365));
  OAI211_X1 g164(.A(G228gat), .B(G233gat), .C1(new_n363), .C2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G22gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n214), .ZN(new_n368));
  NAND2_X1  g167(.A1(G228gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n283), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n210), .A2(new_n203), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT29), .B1(new_n210), .B2(new_n203), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n368), .B(new_n369), .C1(new_n282), .C2(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n366), .A2(new_n367), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n367), .B1(new_n366), .B2(new_n374), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n360), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n359), .A2(KEYINPUT77), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n378), .B(KEYINPUT78), .Z(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n360), .B(new_n379), .C1(new_n375), .C2(new_n376), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n356), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT83), .B1(new_n343), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT69), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT36), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(KEYINPUT69), .A2(KEYINPUT36), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n257), .A2(new_n294), .ZN(new_n390));
  INV_X1    g189(.A(G227gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(new_n254), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n239), .A2(new_n306), .A3(new_n251), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n390), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n395), .B(KEYINPUT34), .Z(new_n396));
  INV_X1    g195(.A(new_n394), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n306), .B1(new_n239), .B2(new_n251), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n392), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT68), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n393), .B1(new_n390), .B2(new_n394), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT68), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT33), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G15gat), .B(G43gat), .Z(new_n405));
  XNOR2_X1  g204(.A(G71gat), .B(G99gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n396), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n402), .A2(KEYINPUT68), .ZN(new_n410));
  AOI211_X1 g209(.A(new_n400), .B(new_n393), .C1(new_n390), .C2(new_n394), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT32), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT33), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n410), .B2(new_n411), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n395), .B(KEYINPUT34), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n407), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n409), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n409), .B2(new_n418), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n388), .B(new_n389), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n409), .A2(new_n418), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT32), .B1(new_n410), .B2(new_n411), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n414), .A3(new_n418), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n424), .A2(new_n386), .A3(new_n387), .A4(new_n425), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n345), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n299), .A2(new_n310), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n311), .A2(new_n314), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n319), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n344), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI22_X1  g232(.A1(new_n433), .A2(KEYINPUT76), .B1(new_n319), .B2(new_n315), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n433), .A2(KEYINPUT76), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n428), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n270), .A2(new_n272), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n383), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n330), .B1(new_n333), .B2(new_n334), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n324), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(new_n335), .A3(new_n322), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n443), .A2(new_n444), .A3(new_n383), .A4(new_n356), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n385), .A2(new_n427), .A3(new_n440), .A4(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n419), .A2(new_n420), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n383), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT35), .B1(new_n448), .B2(new_n438), .ZN(new_n449));
  INV_X1    g248(.A(new_n437), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT84), .B(KEYINPUT35), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n450), .A2(new_n348), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(new_n447), .A3(new_n383), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT85), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n446), .A2(KEYINPUT85), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(G50gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n460), .A2(G43gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(G43gat), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n461), .B1(KEYINPUT88), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(KEYINPUT88), .B2(new_n462), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT15), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G43gat), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(G50gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(new_n461), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n465), .B1(new_n469), .B2(KEYINPUT86), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(new_n468), .B2(new_n461), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G29gat), .A2(G36gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT89), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n476));
  OR3_X1    g275(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n466), .A2(new_n473), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT87), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n476), .A2(new_n480), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n477), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n474), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n472), .A3(new_n470), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT16), .ZN(new_n490));
  AOI21_X1  g289(.A(G1gat), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n489), .B(new_n492), .C1(new_n490), .C2(G1gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT91), .B(G8gat), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G8gat), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n494), .A2(new_n495), .B1(KEYINPUT91), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n479), .A2(KEYINPUT17), .A3(new_n485), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n486), .B1(new_n499), .B2(new_n501), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT18), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n504), .A2(KEYINPUT18), .A3(new_n505), .A4(new_n506), .ZN(new_n510));
  INV_X1    g309(.A(new_n501), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n511), .A2(new_n479), .A3(new_n485), .A4(new_n498), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n506), .A2(KEYINPUT92), .A3(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n505), .B(KEYINPUT13), .Z(new_n514));
  INV_X1    g313(.A(KEYINPUT92), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n502), .A2(new_n515), .A3(new_n485), .A4(new_n479), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n509), .A2(new_n510), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G113gat), .B(G141gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(G197gat), .ZN(new_n520));
  XOR2_X1   g319(.A(KEYINPUT11), .B(G169gat), .Z(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT12), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n509), .A2(new_n523), .A3(new_n510), .A4(new_n517), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(G85gat), .A3(G92gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533));
  INV_X1    g332(.A(G85gat), .ZN(new_n534));
  INV_X1    g333(.A(G92gat), .ZN(new_n535));
  AOI22_X1  g334(.A1(KEYINPUT8), .A2(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G99gat), .B(G106gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n532), .A2(new_n536), .A3(new_n538), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n486), .A2(new_n543), .B1(KEYINPUT41), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n503), .A2(new_n542), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT17), .B1(new_n479), .B2(new_n485), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G190gat), .B(G218gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT98), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n544), .A2(KEYINPUT41), .ZN(new_n552));
  XNOR2_X1  g351(.A(G134gat), .B(G162gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n550), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n545), .B(new_n555), .C1(new_n546), .C2(new_n547), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n551), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n554), .B1(new_n551), .B2(new_n556), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT93), .B1(G71gat), .B2(G78gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(KEYINPUT93), .A2(G71gat), .A3(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(G71gat), .ZN(new_n565));
  INV_X1    g364(.A(G78gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n563), .A2(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G57gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT94), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT94), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(G57gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n571), .A3(G64gat), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(G64gat), .B1(new_n569), .B2(new_n571), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n567), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(new_n568), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(G64gat), .ZN(new_n581));
  INV_X1    g380(.A(G64gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(KEYINPUT96), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT9), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(new_n565), .B2(new_n566), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(KEYINPUT96), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n580), .A2(G64gat), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n587), .B(new_n588), .C1(new_n578), .C2(new_n568), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n584), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n577), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  OAI21_X1  g394(.A(new_n502), .B1(new_n592), .B2(new_n591), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT97), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G183gat), .B(G211gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n597), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n561), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G120gat), .B(G148gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(G176gat), .B(G204gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n565), .A2(new_n566), .ZN(new_n609));
  INV_X1    g408(.A(new_n564), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(new_n562), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT94), .B(G57gat), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n573), .B1(new_n612), .B2(G64gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n569), .A2(new_n571), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n582), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n611), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n584), .A2(new_n589), .A3(new_n586), .ZN(new_n617));
  INV_X1    g416(.A(new_n541), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n538), .B1(new_n532), .B2(new_n536), .ZN(new_n619));
  OAI22_X1  g418(.A1(new_n616), .A2(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n577), .A2(new_n590), .A3(new_n541), .A4(new_n540), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n591), .A2(KEYINPUT99), .A3(new_n542), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n622), .A2(new_n626), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n631), .B(KEYINPUT100), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n625), .A2(new_n631), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n608), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT10), .B1(new_n623), .B2(new_n624), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n631), .B1(new_n638), .B2(new_n628), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n639), .A2(new_n636), .A3(new_n608), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n605), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n459), .A2(new_n527), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n643), .A2(new_n436), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT101), .B(G1gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1324gat));
  NOR2_X1   g445(.A1(new_n643), .A2(new_n437), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT102), .B1(new_n647), .B2(new_n500), .ZN(new_n648));
  OR3_X1    g447(.A1(new_n647), .A2(KEYINPUT102), .A3(new_n500), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n651), .A2(KEYINPUT42), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(KEYINPUT42), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n648), .B(new_n649), .C1(new_n652), .C2(new_n653), .ZN(G1325gat));
  OAI21_X1  g453(.A(G15gat), .B1(new_n643), .B2(new_n427), .ZN(new_n655));
  INV_X1    g454(.A(new_n447), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(G15gat), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n655), .B1(new_n643), .B2(new_n657), .ZN(G1326gat));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n383), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT43), .B(G22gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  NOR3_X1   g460(.A1(new_n561), .A2(new_n604), .A3(new_n641), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n459), .A2(new_n527), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n436), .ZN(new_n664));
  INV_X1    g463(.A(G29gat), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OR3_X1    g465(.A1(new_n663), .A2(KEYINPUT103), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT103), .B1(new_n663), .B2(new_n666), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT45), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n637), .A2(new_n640), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(KEYINPUT104), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(KEYINPUT104), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n527), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n676), .A2(new_n677), .A3(new_n604), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n446), .A2(KEYINPUT85), .A3(new_n454), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT85), .B1(new_n446), .B2(new_n454), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n560), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT44), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n560), .A2(KEYINPUT106), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n558), .B2(new_n559), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n455), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n679), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n664), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G29gat), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n667), .A2(KEYINPUT45), .A3(new_n668), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n671), .A2(new_n692), .A3(new_n693), .ZN(G1328gat));
  INV_X1    g493(.A(G36gat), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n696), .B2(KEYINPUT107), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n663), .A2(new_n437), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(KEYINPUT107), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n682), .A2(KEYINPUT44), .B1(new_n455), .B2(new_n688), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(new_n437), .A3(new_n679), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n702), .B2(new_n695), .ZN(G1329gat));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704));
  INV_X1    g503(.A(new_n427), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n467), .B1(new_n690), .B2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n663), .A2(G43gat), .A3(new_n656), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n707), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n701), .A2(new_n427), .A3(new_n679), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n709), .B(KEYINPUT47), .C1(new_n710), .C2(new_n467), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(G1330gat));
  NOR4_X1   g511(.A1(new_n701), .A2(new_n460), .A3(new_n383), .A4(new_n679), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n460), .B1(new_n663), .B2(new_n383), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT48), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n690), .A2(G50gat), .A3(new_n439), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n718), .A3(new_n714), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(G1331gat));
  NOR3_X1   g519(.A1(new_n675), .A2(new_n527), .A3(new_n605), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n455), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n436), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(new_n568), .ZN(G1332gat));
  XNOR2_X1  g523(.A(new_n437), .B(KEYINPUT108), .ZN(new_n725));
  AOI211_X1 g524(.A(new_n725), .B(new_n722), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1333gat));
  NOR3_X1   g527(.A1(new_n722), .A2(new_n565), .A3(new_n427), .ZN(new_n729));
  INV_X1    g528(.A(new_n722), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT109), .B1(new_n730), .B2(new_n447), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(G71gat), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(KEYINPUT109), .A3(new_n447), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1334gat));
  NOR2_X1   g535(.A1(new_n722), .A2(new_n383), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(new_n566), .ZN(G1335gat));
  INV_X1    g537(.A(new_n604), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n677), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT111), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n641), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n701), .A2(new_n436), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n455), .A2(KEYINPUT51), .A3(new_n560), .A4(new_n741), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n455), .A2(new_n560), .A3(new_n741), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n746), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n664), .A2(new_n534), .A3(new_n641), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n743), .A2(new_n534), .B1(new_n752), .B2(new_n753), .ZN(G1336gat));
  NOR3_X1   g553(.A1(new_n725), .A2(G92gat), .A3(new_n675), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT52), .B1(new_n751), .B2(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n701), .A2(new_n725), .A3(new_n742), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(new_n535), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n683), .A2(new_n689), .ZN(new_n759));
  INV_X1    g558(.A(new_n742), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n450), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n750), .A2(new_n744), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n761), .A2(G92gat), .B1(new_n762), .B2(new_n755), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n758), .B1(new_n763), .B2(new_n764), .ZN(G1337gat));
  NOR3_X1   g564(.A1(new_n701), .A2(new_n427), .A3(new_n742), .ZN(new_n766));
  INV_X1    g565(.A(G99gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n447), .A2(new_n767), .A3(new_n641), .ZN(new_n768));
  OAI22_X1  g567(.A1(new_n766), .A2(new_n767), .B1(new_n752), .B2(new_n768), .ZN(G1338gat));
  NOR3_X1   g568(.A1(new_n675), .A2(new_n383), .A3(G106gat), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT53), .B1(new_n751), .B2(new_n770), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n701), .A2(new_n383), .A3(new_n742), .ZN(new_n772));
  INV_X1    g571(.A(G106gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n439), .A3(new_n760), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n775), .A2(G106gat), .B1(new_n762), .B2(new_n770), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(G1339gat));
  NAND2_X1  g577(.A1(new_n685), .A2(new_n687), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n780), .B(new_n633), .C1(new_n638), .C2(new_n628), .ZN(new_n781));
  INV_X1    g580(.A(new_n608), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n780), .B1(new_n630), .B2(new_n631), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n627), .A2(new_n632), .A3(new_n629), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT114), .B1(new_n786), .B2(KEYINPUT55), .ZN(new_n787));
  INV_X1    g586(.A(new_n783), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n785), .A2(KEYINPUT54), .A3(new_n639), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n787), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n789), .A2(KEYINPUT55), .A3(new_n782), .A4(new_n781), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n788), .A2(KEYINPUT113), .A3(new_n789), .A4(KEYINPUT55), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n640), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n794), .A2(new_n799), .A3(new_n527), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n514), .B1(new_n513), .B2(new_n516), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n522), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n526), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n641), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n779), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  AND4_X1   g605(.A1(new_n779), .A2(new_n794), .A3(new_n799), .A4(new_n804), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n739), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n642), .A2(new_n677), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n439), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n664), .A3(new_n447), .A4(new_n725), .ZN(new_n811));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n677), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n436), .B1(new_n808), .B2(new_n809), .ZN(new_n813));
  INV_X1    g612(.A(new_n448), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n813), .A2(new_n814), .A3(new_n725), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n677), .A2(G113gat), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT115), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n812), .A2(new_n818), .ZN(G1340gat));
  AOI21_X1  g618(.A(G120gat), .B1(new_n815), .B2(new_n641), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n811), .A2(new_n289), .A3(new_n675), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(G1341gat));
  INV_X1    g621(.A(G127gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n815), .A2(new_n823), .A3(new_n604), .ZN(new_n824));
  OAI21_X1  g623(.A(G127gat), .B1(new_n811), .B2(new_n739), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(G1342gat));
  NOR3_X1   g625(.A1(new_n450), .A2(G134gat), .A3(new_n561), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n813), .A2(new_n814), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(KEYINPUT56), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT116), .Z(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(KEYINPUT56), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT117), .Z(new_n832));
  OAI21_X1  g631(.A(G134gat), .B1(new_n811), .B2(new_n561), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(G1343gat));
  NAND2_X1  g633(.A1(new_n427), .A2(new_n439), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT121), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n813), .A2(KEYINPUT120), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n813), .A2(KEYINPUT120), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n725), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  OR3_X1    g638(.A1(new_n839), .A2(G141gat), .A3(new_n677), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n427), .A2(new_n664), .A3(new_n725), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n808), .A2(new_n809), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT57), .B1(new_n843), .B2(new_n439), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n439), .A2(KEYINPUT57), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n846), .B1(new_n804), .B2(new_n641), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n526), .A2(new_n803), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n672), .A2(new_n848), .A3(KEYINPUT118), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n790), .A2(new_n792), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n799), .A2(new_n527), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n560), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n739), .B1(new_n853), .B2(new_n807), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n845), .B1(new_n854), .B2(new_n809), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n842), .B1(new_n844), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G141gat), .B1(new_n856), .B2(new_n677), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g659(.A(KEYINPUT119), .B(new_n842), .C1(new_n844), .C2(new_n855), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n527), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(G141gat), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n863), .A2(new_n840), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n858), .B1(new_n864), .B2(new_n841), .ZN(G1344gat));
  NAND2_X1  g664(.A1(new_n842), .A2(new_n641), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  INV_X1    g666(.A(new_n809), .ZN(new_n868));
  AND4_X1   g667(.A1(new_n560), .A2(new_n794), .A3(new_n799), .A4(new_n804), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n853), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n868), .B1(new_n870), .B2(new_n739), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n439), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI211_X1 g672(.A(KEYINPUT123), .B(new_n868), .C1(new_n870), .C2(new_n739), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n867), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n843), .A2(KEYINPUT57), .A3(new_n439), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n866), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(G148gat), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT59), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n860), .A2(new_n641), .A3(new_n861), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n878), .A2(KEYINPUT59), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n880), .A2(KEYINPUT122), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT122), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OR3_X1    g683(.A1(new_n839), .A2(G148gat), .A3(new_n672), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1345gat));
  NAND4_X1  g685(.A1(new_n860), .A2(G155gat), .A3(new_n604), .A4(new_n861), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n274), .B1(new_n839), .B2(new_n739), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT124), .ZN(G1346gat));
  NOR3_X1   g689(.A1(new_n450), .A2(G162gat), .A3(new_n561), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n836), .B(new_n891), .C1(new_n837), .C2(new_n838), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n860), .A2(new_n779), .A3(new_n861), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n275), .ZN(G1347gat));
  NAND2_X1  g693(.A1(new_n436), .A2(new_n450), .ZN(new_n895));
  XOR2_X1   g694(.A(new_n895), .B(KEYINPUT125), .Z(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n656), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n810), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n899), .A2(G169gat), .A3(new_n527), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n664), .B1(new_n808), .B2(new_n809), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n448), .A2(new_n725), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(G169gat), .B1(new_n903), .B2(new_n527), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n900), .A2(new_n904), .ZN(G1348gat));
  OAI21_X1  g704(.A(G176gat), .B1(new_n898), .B2(new_n675), .ZN(new_n906));
  INV_X1    g705(.A(new_n903), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n672), .A2(G176gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(G1349gat));
  NOR3_X1   g708(.A1(new_n907), .A2(new_n243), .A3(new_n739), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n224), .B1(new_n899), .B2(new_n604), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT126), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT60), .Z(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n898), .B2(new_n561), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT61), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n903), .A2(new_n225), .A3(new_n779), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1351gat));
  INV_X1    g716(.A(G197gat), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n896), .A2(new_n705), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n919), .B1(new_n875), .B2(new_n876), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n918), .B1(new_n920), .B2(new_n527), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n835), .A2(new_n725), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n901), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n918), .A3(new_n527), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT127), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927));
  AOI211_X1 g726(.A(new_n677), .B(new_n919), .C1(new_n875), .C2(new_n876), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n927), .B(new_n924), .C1(new_n928), .C2(new_n918), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n926), .A2(new_n929), .ZN(G1352gat));
  INV_X1    g729(.A(G204gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n923), .A2(new_n931), .A3(new_n641), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT62), .Z(new_n933));
  AND2_X1   g732(.A1(new_n920), .A2(new_n676), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(new_n931), .ZN(G1353gat));
  INV_X1    g734(.A(G211gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n923), .A2(new_n936), .A3(new_n604), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n875), .A2(new_n876), .ZN(new_n938));
  INV_X1    g737(.A(new_n919), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n604), .A3(new_n939), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n940), .B2(G211gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(G1354gat));
  INV_X1    g742(.A(G218gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n923), .A2(new_n944), .A3(new_n779), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n920), .A2(new_n560), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n944), .ZN(G1355gat));
endmodule


