

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774;

  NOR2_X1 U367 ( .A1(n745), .A2(n744), .ZN(n422) );
  AND2_X1 U368 ( .A1(n416), .A2(n375), .ZN(n376) );
  NAND2_X1 U369 ( .A1(n414), .A2(n378), .ZN(n354) );
  XNOR2_X2 U370 ( .A(n508), .B(G469), .ZN(n414) );
  XNOR2_X2 U371 ( .A(n345), .B(KEYINPUT40), .ZN(n613) );
  NAND2_X2 U372 ( .A1(n584), .A2(n672), .ZN(n345) );
  XNOR2_X2 U373 ( .A(n414), .B(KEYINPUT1), .ZN(n585) );
  NOR2_X2 U374 ( .A1(n450), .A2(n449), .ZN(n642) );
  XNOR2_X1 U375 ( .A(n635), .B(n434), .ZN(n433) );
  INV_X1 U376 ( .A(G953), .ZN(n767) );
  INV_X1 U377 ( .A(n394), .ZN(n635) );
  XNOR2_X1 U378 ( .A(KEYINPUT63), .B(KEYINPUT86), .ZN(n346) );
  XOR2_X1 U379 ( .A(n652), .B(KEYINPUT62), .Z(n347) );
  XOR2_X1 U380 ( .A(n625), .B(n624), .Z(n348) );
  AND2_X1 U381 ( .A1(n647), .A2(n646), .ZN(n397) );
  AND2_X1 U382 ( .A1(n746), .A2(n766), .ZN(n644) );
  XNOR2_X2 U383 ( .A(n532), .B(n480), .ZN(n437) );
  XNOR2_X2 U384 ( .A(n534), .B(n464), .ZN(n751) );
  XNOR2_X2 U385 ( .A(n472), .B(n471), .ZN(n534) );
  XNOR2_X2 U386 ( .A(n608), .B(n607), .ZN(n715) );
  NOR2_X2 U387 ( .A1(n688), .A2(n687), .ZN(n608) );
  NAND2_X1 U388 ( .A1(n364), .A2(n349), .ZN(n363) );
  XNOR2_X1 U389 ( .A(n358), .B(KEYINPUT42), .ZN(n774) );
  INV_X1 U390 ( .A(KEYINPUT97), .ZN(n353) );
  INV_X1 U391 ( .A(KEYINPUT68), .ZN(n470) );
  NOR2_X1 U392 ( .A1(n736), .A2(n744), .ZN(n420) );
  NOR2_X1 U393 ( .A1(n730), .A2(n744), .ZN(n731) );
  XNOR2_X1 U394 ( .A(n365), .B(n347), .ZN(n364) );
  NAND2_X1 U395 ( .A1(n397), .A2(G472), .ZN(n365) );
  NAND2_X1 U396 ( .A1(n415), .A2(n458), .ZN(n419) );
  NOR2_X1 U397 ( .A1(n772), .A2(n663), .ZN(n605) );
  XNOR2_X1 U398 ( .A(n360), .B(KEYINPUT84), .ZN(n582) );
  NAND2_X1 U399 ( .A1(n613), .A2(n774), .ZN(n401) );
  INV_X1 U400 ( .A(n361), .ZN(n705) );
  NAND2_X1 U401 ( .A1(n715), .A2(n623), .ZN(n358) );
  AND2_X1 U402 ( .A1(n413), .A2(n615), .ZN(n601) );
  XNOR2_X1 U403 ( .A(n423), .B(KEYINPUT99), .ZN(n362) );
  XNOR2_X1 U404 ( .A(n440), .B(n380), .ZN(n413) );
  XNOR2_X1 U405 ( .A(n589), .B(n588), .ZN(n684) );
  BUF_X1 U406 ( .A(n594), .Z(n596) );
  NAND2_X1 U407 ( .A1(n355), .A2(n429), .ZN(n423) );
  AND2_X1 U408 ( .A1(n412), .A2(n439), .ZN(n411) );
  NOR2_X1 U409 ( .A1(n674), .A2(n672), .ZN(n689) );
  NOR2_X1 U410 ( .A1(n727), .A2(n640), .ZN(n539) );
  XNOR2_X1 U411 ( .A(n463), .B(n465), .ZN(n727) );
  XNOR2_X1 U412 ( .A(n350), .B(n751), .ZN(n463) );
  OR2_X1 U413 ( .A1(n742), .A2(G902), .ZN(n526) );
  XNOR2_X1 U414 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U415 ( .A(n536), .B(n466), .ZN(n465) );
  XOR2_X1 U416 ( .A(KEYINPUT69), .B(n752), .Z(n535) );
  INV_X1 U417 ( .A(n744), .ZN(n349) );
  INV_X1 U418 ( .A(n386), .ZN(n371) );
  XNOR2_X1 U419 ( .A(n520), .B(G902), .ZN(n640) );
  INV_X1 U420 ( .A(n510), .ZN(n386) );
  XNOR2_X1 U421 ( .A(n438), .B(n470), .ZN(n472) );
  XNOR2_X1 U422 ( .A(G146), .B(G125), .ZN(n531) );
  XNOR2_X1 U423 ( .A(G119), .B(G116), .ZN(n438) );
  XNOR2_X1 U424 ( .A(KEYINPUT24), .B(G128), .ZN(n513) );
  INV_X1 U425 ( .A(n532), .ZN(n350) );
  NAND2_X1 U426 ( .A1(n351), .A2(n600), .ZN(n393) );
  NOR2_X1 U427 ( .A1(n468), .A2(n599), .ZN(n351) );
  NAND2_X1 U428 ( .A1(n411), .A2(n409), .ZN(n594) );
  XNOR2_X2 U429 ( .A(n352), .B(n541), .ZN(n584) );
  NAND2_X1 U430 ( .A1(n455), .A2(n454), .ZN(n352) );
  XNOR2_X2 U431 ( .A(n354), .B(n353), .ZN(n653) );
  XNOR2_X2 U432 ( .A(n448), .B(n462), .ZN(n773) );
  NAND2_X1 U433 ( .A1(n587), .A2(n355), .ZN(n589) );
  XNOR2_X2 U434 ( .A(n586), .B(KEYINPUT73), .ZN(n355) );
  NAND2_X1 U435 ( .A1(n356), .A2(n637), .ZN(n405) );
  NAND2_X1 U436 ( .A1(n357), .A2(n417), .ZN(n356) );
  NAND2_X1 U437 ( .A1(n419), .A2(KEYINPUT81), .ZN(n357) );
  NAND2_X1 U438 ( .A1(n601), .A2(n620), .ZN(n360) );
  NAND2_X1 U439 ( .A1(n362), .A2(n596), .ZN(n595) );
  OR2_X1 U440 ( .A1(n704), .A2(n362), .ZN(n361) );
  XNOR2_X1 U441 ( .A(n363), .B(n346), .ZN(G57) );
  INV_X1 U442 ( .A(n773), .ZN(n366) );
  INV_X1 U443 ( .A(n366), .ZN(n367) );
  BUF_X1 U444 ( .A(n599), .Z(n368) );
  BUF_X1 U445 ( .A(n437), .Z(n369) );
  XNOR2_X2 U446 ( .A(n572), .B(n571), .ZN(n622) );
  NAND2_X1 U447 ( .A1(n437), .A2(n386), .ZN(n372) );
  NAND2_X1 U448 ( .A1(n370), .A2(n371), .ZN(n373) );
  NAND2_X1 U449 ( .A1(n373), .A2(n372), .ZN(n395) );
  INV_X1 U450 ( .A(n437), .ZN(n370) );
  XNOR2_X2 U451 ( .A(n401), .B(n382), .ZN(n461) );
  INV_X1 U452 ( .A(G134), .ZN(n479) );
  NOR2_X1 U453 ( .A1(G902), .A2(G237), .ZN(n490) );
  XOR2_X1 U454 ( .A(G137), .B(KEYINPUT5), .Z(n482) );
  XNOR2_X1 U455 ( .A(G146), .B(G101), .ZN(n484) );
  INV_X1 U456 ( .A(KEYINPUT81), .ZN(n403) );
  XOR2_X1 U457 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n558) );
  XNOR2_X1 U458 ( .A(G107), .B(G134), .ZN(n557) );
  INV_X1 U459 ( .A(G902), .ZN(n507) );
  XNOR2_X1 U460 ( .A(KEYINPUT16), .B(G122), .ZN(n464) );
  XNOR2_X1 U461 ( .A(G140), .B(G137), .ZN(n510) );
  XNOR2_X1 U462 ( .A(KEYINPUT93), .B(KEYINPUT23), .ZN(n509) );
  NOR2_X1 U463 ( .A1(n430), .A2(G953), .ZN(n515) );
  XNOR2_X1 U464 ( .A(n533), .B(n377), .ZN(n436) );
  XNOR2_X1 U465 ( .A(n531), .B(KEYINPUT18), .ZN(n435) );
  NAND2_X1 U466 ( .A1(n444), .A2(n626), .ZN(n443) );
  NAND2_X1 U467 ( .A1(n594), .A2(n469), .ZN(n440) );
  XNOR2_X1 U468 ( .A(n651), .B(KEYINPUT87), .ZN(n744) );
  NAND2_X1 U469 ( .A1(n348), .A2(n424), .ZN(n460) );
  NOR2_X1 U470 ( .A1(n668), .A2(n677), .ZN(n424) );
  INV_X1 U471 ( .A(KEYINPUT44), .ZN(n391) );
  INV_X1 U472 ( .A(KEYINPUT15), .ZN(n520) );
  NAND2_X1 U473 ( .A1(G237), .A2(G234), .ZN(n493) );
  INV_X1 U474 ( .A(n433), .ZN(n432) );
  INV_X1 U475 ( .A(n610), .ZN(n431) );
  NAND2_X1 U476 ( .A1(n596), .A2(n447), .ZN(n446) );
  INV_X1 U477 ( .A(KEYINPUT34), .ZN(n447) );
  NAND2_X1 U478 ( .A1(n410), .A2(n374), .ZN(n409) );
  XNOR2_X1 U479 ( .A(n486), .B(n456), .ZN(n453) );
  NAND2_X1 U480 ( .A1(n405), .A2(n402), .ZN(n766) );
  NAND2_X1 U481 ( .A1(n404), .A2(n376), .ZN(n402) );
  XNOR2_X1 U482 ( .A(G101), .B(G104), .ZN(n500) );
  XNOR2_X1 U483 ( .A(G116), .B(G122), .ZN(n556) );
  XOR2_X1 U484 ( .A(G143), .B(G104), .Z(n549) );
  XNOR2_X1 U485 ( .A(G140), .B(G122), .ZN(n548) );
  XOR2_X1 U486 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n544) );
  XNOR2_X1 U487 ( .A(n653), .B(KEYINPUT105), .ZN(n454) );
  AND2_X1 U488 ( .A1(n499), .A2(n610), .ZN(n452) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n425) );
  INV_X1 U490 ( .A(KEYINPUT28), .ZN(n426) );
  NAND2_X1 U491 ( .A1(n429), .A2(n428), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n519), .B(n518), .ZN(n742) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n466) );
  XNOR2_X1 U494 ( .A(KEYINPUT35), .B(KEYINPUT80), .ZN(n462) );
  XNOR2_X1 U495 ( .A(n408), .B(n602), .ZN(n772) );
  AND2_X1 U496 ( .A1(n568), .A2(n697), .ZN(n467) );
  NAND2_X1 U497 ( .A1(n623), .A2(n410), .ZN(n669) );
  NOR2_X1 U498 ( .A1(n580), .A2(n379), .ZN(n374) );
  AND2_X1 U499 ( .A1(n637), .A2(n403), .ZN(n375) );
  XNOR2_X1 U500 ( .A(KEYINPUT88), .B(KEYINPUT17), .ZN(n377) );
  XNOR2_X1 U501 ( .A(n526), .B(n525), .ZN(n697) );
  NOR2_X1 U502 ( .A1(n697), .A2(n696), .ZN(n378) );
  INV_X1 U503 ( .A(G234), .ZN(n430) );
  XOR2_X1 U504 ( .A(KEYINPUT66), .B(KEYINPUT0), .Z(n379) );
  XNOR2_X1 U505 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n380) );
  XNOR2_X1 U506 ( .A(n398), .B(n648), .ZN(n381) );
  XOR2_X1 U507 ( .A(KEYINPUT82), .B(KEYINPUT46), .Z(n382) );
  INV_X1 U508 ( .A(KEYINPUT48), .ZN(n631) );
  NOR2_X1 U509 ( .A1(KEYINPUT79), .A2(n639), .ZN(n383) );
  AND2_X1 U510 ( .A1(KEYINPUT48), .A2(KEYINPUT81), .ZN(n384) );
  XNOR2_X1 U511 ( .A(n395), .B(n385), .ZN(n649) );
  INV_X1 U512 ( .A(n506), .ZN(n385) );
  XNOR2_X2 U513 ( .A(n387), .B(KEYINPUT45), .ZN(n746) );
  NAND2_X1 U514 ( .A1(n392), .A2(n388), .ZN(n387) );
  NAND2_X1 U515 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U516 ( .A1(n605), .A2(n367), .ZN(n389) );
  XNOR2_X1 U517 ( .A(n605), .B(n391), .ZN(n390) );
  XNOR2_X1 U518 ( .A(n393), .B(KEYINPUT85), .ZN(n392) );
  BUF_X1 U519 ( .A(n570), .Z(n394) );
  INV_X1 U520 ( .A(n395), .ZN(n396) );
  AND2_X2 U521 ( .A1(n647), .A2(n646), .ZN(n400) );
  NAND2_X1 U522 ( .A1(n397), .A2(G469), .ZN(n399) );
  XNOR2_X1 U523 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U524 ( .A1(n590), .A2(KEYINPUT34), .ZN(n444) );
  XNOR2_X1 U525 ( .A(n396), .B(n506), .ZN(n398) );
  BUF_X1 U526 ( .A(n684), .Z(n716) );
  XNOR2_X1 U527 ( .A(n399), .B(n381), .ZN(n407) );
  NAND2_X1 U528 ( .A1(n400), .A2(G217), .ZN(n743) );
  NAND2_X1 U529 ( .A1(n400), .A2(G210), .ZN(n729) );
  NAND2_X1 U530 ( .A1(n400), .A2(G475), .ZN(n735) );
  NAND2_X1 U531 ( .A1(n397), .A2(G478), .ZN(n740) );
  INV_X1 U532 ( .A(n419), .ZN(n404) );
  XNOR2_X1 U533 ( .A(n406), .B(KEYINPUT117), .ZN(G54) );
  NAND2_X1 U534 ( .A1(n407), .A2(n349), .ZN(n406) );
  NAND2_X1 U535 ( .A1(n601), .A2(n467), .ZN(n408) );
  INV_X1 U536 ( .A(n622), .ZN(n410) );
  NAND2_X1 U537 ( .A1(n622), .A2(n379), .ZN(n412) );
  NAND2_X1 U538 ( .A1(n413), .A2(n620), .ZN(n604) );
  AND2_X1 U539 ( .A1(n414), .A2(n425), .ZN(n623) );
  NAND2_X1 U540 ( .A1(n461), .A2(n457), .ZN(n415) );
  NAND2_X1 U541 ( .A1(n418), .A2(KEYINPUT48), .ZN(n416) );
  NAND2_X1 U542 ( .A1(n418), .A2(n384), .ZN(n417) );
  INV_X1 U543 ( .A(n461), .ZN(n418) );
  XNOR2_X1 U544 ( .A(n420), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U545 ( .A(KEYINPUT4), .ZN(n474) );
  NAND2_X1 U546 ( .A1(n421), .A2(n643), .ZN(n647) );
  NOR2_X1 U547 ( .A1(n642), .A2(n641), .ZN(n421) );
  XNOR2_X1 U548 ( .A(n422), .B(KEYINPUT120), .ZN(G66) );
  NOR2_X2 U549 ( .A1(n675), .A2(n597), .ZN(n598) );
  XNOR2_X2 U550 ( .A(n595), .B(KEYINPUT31), .ZN(n675) );
  NOR2_X1 U551 ( .A1(n582), .A2(n697), .ZN(n599) );
  INV_X1 U552 ( .A(n460), .ZN(n630) );
  NOR2_X1 U553 ( .A1(n612), .A2(n616), .ZN(n428) );
  INV_X1 U554 ( .A(n700), .ZN(n429) );
  NOR2_X1 U555 ( .A1(n433), .A2(n431), .ZN(n451) );
  NAND2_X1 U556 ( .A1(n432), .A2(n685), .ZN(n688) );
  AND2_X1 U557 ( .A1(n433), .A2(n491), .ZN(n686) );
  INV_X1 U558 ( .A(KEYINPUT38), .ZN(n434) );
  XNOR2_X1 U559 ( .A(n369), .B(n453), .ZN(n652) );
  NAND2_X1 U560 ( .A1(n580), .A2(n379), .ZN(n439) );
  NAND2_X1 U561 ( .A1(n442), .A2(n441), .ZN(n448) );
  NAND2_X1 U562 ( .A1(n684), .A2(KEYINPUT34), .ZN(n441) );
  NOR2_X1 U563 ( .A1(n445), .A2(n443), .ZN(n442) );
  NOR2_X1 U564 ( .A1(n684), .A2(n446), .ZN(n445) );
  INV_X1 U565 ( .A(n746), .ZN(n449) );
  NAND2_X1 U566 ( .A1(n766), .A2(n383), .ZN(n450) );
  INV_X1 U567 ( .A(n645), .ZN(n681) );
  AND2_X1 U568 ( .A1(n499), .A2(n451), .ZN(n455) );
  AND2_X1 U569 ( .A1(n454), .A2(n452), .ZN(n629) );
  XNOR2_X2 U570 ( .A(n478), .B(KEYINPUT64), .ZN(n532) );
  XNOR2_X2 U571 ( .A(n502), .B(n501), .ZN(n752) );
  INV_X1 U572 ( .A(n535), .ZN(n536) );
  XNOR2_X1 U573 ( .A(n489), .B(n488), .ZN(n569) );
  AND2_X1 U574 ( .A1(n459), .A2(n679), .ZN(n458) );
  INV_X1 U575 ( .A(n534), .ZN(n456) );
  AND2_X1 U576 ( .A1(n630), .A2(n631), .ZN(n457) );
  NAND2_X1 U577 ( .A1(n460), .A2(KEYINPUT48), .ZN(n459) );
  NOR2_X1 U578 ( .A1(n598), .A2(n689), .ZN(n468) );
  NOR2_X1 U579 ( .A1(n696), .A2(n687), .ZN(n469) );
  XNOR2_X1 U580 ( .A(n479), .B(G131), .ZN(n480) );
  INV_X1 U581 ( .A(KEYINPUT19), .ZN(n571) );
  XNOR2_X1 U582 ( .A(n487), .B(G472), .ZN(n488) );
  XNOR2_X1 U583 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U584 ( .A(n740), .B(n739), .ZN(n741) );
  XOR2_X1 U585 ( .A(KEYINPUT3), .B(G113), .Z(n471) );
  XNOR2_X2 U586 ( .A(G128), .B(KEYINPUT77), .ZN(n473) );
  XNOR2_X2 U587 ( .A(n473), .B(G143), .ZN(n555) );
  INV_X1 U588 ( .A(n555), .ZN(n475) );
  NAND2_X1 U589 ( .A1(n475), .A2(n474), .ZN(n477) );
  NAND2_X1 U590 ( .A1(n555), .A2(KEYINPUT4), .ZN(n476) );
  NAND2_X1 U591 ( .A1(n477), .A2(n476), .ZN(n478) );
  NOR2_X2 U592 ( .A1(G953), .A2(G237), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n542), .A2(G210), .ZN(n481) );
  XNOR2_X1 U594 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U595 ( .A(n483), .B(KEYINPUT75), .Z(n485) );
  XNOR2_X1 U596 ( .A(n485), .B(n484), .ZN(n486) );
  NOR2_X1 U597 ( .A1(G902), .A2(n652), .ZN(n489) );
  XNOR2_X1 U598 ( .A(KEYINPUT72), .B(KEYINPUT98), .ZN(n487) );
  BUF_X2 U599 ( .A(n569), .Z(n700) );
  XOR2_X1 U600 ( .A(KEYINPUT74), .B(n490), .Z(n537) );
  NAND2_X1 U601 ( .A1(n537), .A2(G214), .ZN(n685) );
  INV_X1 U602 ( .A(n685), .ZN(n491) );
  NOR2_X1 U603 ( .A1(n700), .A2(n491), .ZN(n492) );
  XNOR2_X1 U604 ( .A(n492), .B(KEYINPUT30), .ZN(n499) );
  XOR2_X1 U605 ( .A(KEYINPUT14), .B(KEYINPUT89), .Z(n494) );
  XNOR2_X1 U606 ( .A(n494), .B(n493), .ZN(n496) );
  NAND2_X1 U607 ( .A1(n496), .A2(G952), .ZN(n495) );
  XOR2_X1 U608 ( .A(KEYINPUT90), .B(n495), .Z(n713) );
  NAND2_X1 U609 ( .A1(n713), .A2(n767), .ZN(n573) );
  NAND2_X1 U610 ( .A1(G902), .A2(n496), .ZN(n574) );
  NOR2_X1 U611 ( .A1(G900), .A2(n574), .ZN(n497) );
  NAND2_X1 U612 ( .A1(n497), .A2(G953), .ZN(n498) );
  NAND2_X1 U613 ( .A1(n573), .A2(n498), .ZN(n610) );
  INV_X1 U614 ( .A(n500), .ZN(n502) );
  XNOR2_X1 U615 ( .A(G110), .B(G107), .ZN(n501) );
  XOR2_X1 U616 ( .A(G146), .B(KEYINPUT76), .Z(n504) );
  NAND2_X1 U617 ( .A1(G227), .A2(n767), .ZN(n503) );
  XNOR2_X1 U618 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U619 ( .A(n535), .B(n505), .ZN(n506) );
  NAND2_X1 U620 ( .A1(n649), .A2(n507), .ZN(n508) );
  XNOR2_X1 U621 ( .A(n531), .B(KEYINPUT10), .ZN(n759) );
  XNOR2_X1 U622 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U623 ( .A(n759), .B(n511), .ZN(n519) );
  INV_X1 U624 ( .A(G119), .ZN(n512) );
  XNOR2_X1 U625 ( .A(n512), .B(G110), .ZN(n514) );
  XNOR2_X1 U626 ( .A(n514), .B(n513), .ZN(n517) );
  XNOR2_X1 U627 ( .A(KEYINPUT8), .B(n515), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n561), .A2(G221), .ZN(n516) );
  XNOR2_X1 U629 ( .A(n517), .B(n516), .ZN(n518) );
  OR2_X1 U630 ( .A1(n640), .A2(n430), .ZN(n521) );
  XNOR2_X1 U631 ( .A(n521), .B(KEYINPUT20), .ZN(n527) );
  AND2_X1 U632 ( .A1(n527), .A2(G217), .ZN(n524) );
  XNOR2_X1 U633 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n522) );
  XNOR2_X1 U634 ( .A(n522), .B(KEYINPUT25), .ZN(n523) );
  XNOR2_X1 U635 ( .A(n524), .B(n523), .ZN(n525) );
  NAND2_X1 U636 ( .A1(n527), .A2(G221), .ZN(n530) );
  INV_X1 U637 ( .A(KEYINPUT96), .ZN(n528) );
  XNOR2_X1 U638 ( .A(n528), .B(KEYINPUT21), .ZN(n529) );
  XNOR2_X1 U639 ( .A(n530), .B(n529), .ZN(n609) );
  INV_X1 U640 ( .A(n609), .ZN(n696) );
  NAND2_X1 U641 ( .A1(G224), .A2(n767), .ZN(n533) );
  NAND2_X1 U642 ( .A1(G210), .A2(n537), .ZN(n538) );
  XNOR2_X1 U643 ( .A(n539), .B(n538), .ZN(n570) );
  XNOR2_X1 U644 ( .A(KEYINPUT83), .B(KEYINPUT39), .ZN(n540) );
  XNOR2_X1 U645 ( .A(n540), .B(KEYINPUT71), .ZN(n541) );
  NAND2_X1 U646 ( .A1(n542), .A2(G214), .ZN(n543) );
  XNOR2_X1 U647 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U648 ( .A(n545), .B(KEYINPUT11), .Z(n547) );
  XNOR2_X1 U649 ( .A(G113), .B(G131), .ZN(n546) );
  XNOR2_X1 U650 ( .A(n547), .B(n546), .ZN(n552) );
  XNOR2_X1 U651 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U652 ( .A(n759), .B(n550), .ZN(n551) );
  XNOR2_X1 U653 ( .A(n552), .B(n551), .ZN(n733) );
  OR2_X1 U654 ( .A1(n733), .A2(G902), .ZN(n554) );
  XOR2_X1 U655 ( .A(KEYINPUT13), .B(G475), .Z(n553) );
  XNOR2_X1 U656 ( .A(n554), .B(n553), .ZN(n592) );
  INV_X1 U657 ( .A(n592), .ZN(n567) );
  XNOR2_X1 U658 ( .A(n556), .B(KEYINPUT101), .ZN(n560) );
  XNOR2_X1 U659 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U660 ( .A(n560), .B(n559), .Z(n563) );
  NAND2_X1 U661 ( .A1(G217), .A2(n561), .ZN(n562) );
  XNOR2_X1 U662 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U663 ( .A(n555), .B(n564), .ZN(n738) );
  NOR2_X1 U664 ( .A1(G902), .A2(n738), .ZN(n566) );
  INV_X1 U665 ( .A(G478), .ZN(n565) );
  XNOR2_X1 U666 ( .A(n566), .B(n565), .ZN(n591) );
  AND2_X1 U667 ( .A1(n567), .A2(n591), .ZN(n674) );
  NAND2_X1 U668 ( .A1(n584), .A2(n674), .ZN(n637) );
  XNOR2_X1 U669 ( .A(n637), .B(G134), .ZN(G36) );
  BUF_X1 U670 ( .A(n585), .Z(n568) );
  INV_X1 U671 ( .A(n568), .ZN(n620) );
  XOR2_X1 U672 ( .A(n569), .B(KEYINPUT6), .Z(n615) );
  INV_X1 U673 ( .A(n615), .ZN(n587) );
  NAND2_X1 U674 ( .A1(n570), .A2(n685), .ZN(n572) );
  INV_X1 U675 ( .A(n573), .ZN(n578) );
  INV_X1 U676 ( .A(n574), .ZN(n575) );
  NOR2_X1 U677 ( .A1(G898), .A2(n767), .ZN(n754) );
  NAND2_X1 U678 ( .A1(n575), .A2(n754), .ZN(n576) );
  XNOR2_X1 U679 ( .A(KEYINPUT91), .B(n576), .ZN(n577) );
  NOR2_X1 U680 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U681 ( .A(n579), .B(KEYINPUT92), .ZN(n580) );
  NOR2_X1 U682 ( .A1(n591), .A2(n592), .ZN(n581) );
  XOR2_X1 U683 ( .A(KEYINPUT102), .B(n581), .Z(n687) );
  XOR2_X1 U684 ( .A(n368), .B(G101), .Z(G3) );
  INV_X1 U685 ( .A(n591), .ZN(n583) );
  AND2_X1 U686 ( .A1(n583), .A2(n592), .ZN(n672) );
  XNOR2_X1 U687 ( .A(n613), .B(G131), .ZN(G33) );
  NAND2_X1 U688 ( .A1(n585), .A2(n378), .ZN(n586) );
  XOR2_X1 U689 ( .A(KEYINPUT33), .B(KEYINPUT70), .Z(n588) );
  INV_X1 U690 ( .A(n596), .ZN(n590) );
  NAND2_X1 U691 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U692 ( .A(n593), .B(KEYINPUT103), .ZN(n626) );
  NAND2_X1 U693 ( .A1(n773), .A2(KEYINPUT44), .ZN(n600) );
  NAND2_X1 U694 ( .A1(n596), .A2(n700), .ZN(n656) );
  NOR2_X1 U695 ( .A1(n656), .A2(n653), .ZN(n597) );
  INV_X1 U696 ( .A(n697), .ZN(n612) );
  INV_X1 U697 ( .A(KEYINPUT32), .ZN(n602) );
  NAND2_X1 U698 ( .A1(n700), .A2(n697), .ZN(n603) );
  NOR2_X1 U699 ( .A1(n604), .A2(n603), .ZN(n663) );
  XNOR2_X1 U700 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n606) );
  XNOR2_X1 U701 ( .A(n606), .B(KEYINPUT41), .ZN(n607) );
  NAND2_X1 U702 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U703 ( .A(n611), .B(KEYINPUT67), .Z(n616) );
  NAND2_X1 U704 ( .A1(n697), .A2(n685), .ZN(n614) );
  NOR2_X1 U705 ( .A1(n615), .A2(n614), .ZN(n618) );
  INV_X1 U706 ( .A(n672), .ZN(n670) );
  NOR2_X1 U707 ( .A1(n670), .A2(n616), .ZN(n617) );
  NAND2_X1 U708 ( .A1(n618), .A2(n617), .ZN(n632) );
  NOR2_X1 U709 ( .A1(n635), .A2(n632), .ZN(n619) );
  XOR2_X1 U710 ( .A(KEYINPUT36), .B(n619), .Z(n621) );
  NOR2_X1 U711 ( .A1(n621), .A2(n620), .ZN(n677) );
  NOR2_X1 U712 ( .A1(n669), .A2(n689), .ZN(n625) );
  INV_X1 U713 ( .A(KEYINPUT47), .ZN(n624) );
  INV_X1 U714 ( .A(n626), .ZN(n627) );
  NOR2_X1 U715 ( .A1(n635), .A2(n627), .ZN(n628) );
  AND2_X1 U716 ( .A1(n629), .A2(n628), .ZN(n668) );
  OR2_X1 U717 ( .A1(n632), .A2(n568), .ZN(n634) );
  XNOR2_X1 U718 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n633) );
  XNOR2_X1 U719 ( .A(n634), .B(n633), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n636), .A2(n635), .ZN(n679) );
  NAND2_X1 U721 ( .A1(n644), .A2(n640), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n638), .A2(KEYINPUT79), .ZN(n643) );
  INV_X1 U723 ( .A(n640), .ZN(n639) );
  AND2_X1 U724 ( .A1(n640), .A2(KEYINPUT2), .ZN(n641) );
  BUF_X1 U725 ( .A(n644), .Z(n645) );
  NAND2_X1 U726 ( .A1(n645), .A2(KEYINPUT2), .ZN(n646) );
  XOR2_X1 U727 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n648) );
  INV_X1 U728 ( .A(G952), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n650), .A2(G953), .ZN(n651) );
  NOR2_X1 U730 ( .A1(n656), .A2(n670), .ZN(n654) );
  INV_X1 U731 ( .A(n653), .ZN(n657) );
  NAND2_X1 U732 ( .A1(n654), .A2(n657), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n655), .B(G104), .ZN(G6) );
  XNOR2_X1 U734 ( .A(G107), .B(KEYINPUT27), .ZN(n662) );
  XOR2_X1 U735 ( .A(KEYINPUT108), .B(KEYINPUT26), .Z(n660) );
  INV_X1 U736 ( .A(n674), .ZN(n664) );
  NOR2_X1 U737 ( .A1(n656), .A2(n664), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U739 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U740 ( .A(n662), .B(n661), .ZN(G9) );
  XOR2_X1 U741 ( .A(G110), .B(n663), .Z(G12) );
  NOR2_X1 U742 ( .A1(n664), .A2(n669), .ZN(n666) );
  XNOR2_X1 U743 ( .A(KEYINPUT109), .B(KEYINPUT29), .ZN(n665) );
  XNOR2_X1 U744 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U745 ( .A(G128), .B(n667), .Z(G30) );
  XOR2_X1 U746 ( .A(G143), .B(n668), .Z(G45) );
  NOR2_X1 U747 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U748 ( .A(G146), .B(n671), .Z(G48) );
  NAND2_X1 U749 ( .A1(n675), .A2(n672), .ZN(n673) );
  XNOR2_X1 U750 ( .A(n673), .B(G113), .ZN(G15) );
  NAND2_X1 U751 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U752 ( .A(n676), .B(G116), .ZN(G18) );
  XNOR2_X1 U753 ( .A(G125), .B(n677), .ZN(n678) );
  XNOR2_X1 U754 ( .A(n678), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U755 ( .A(G140), .B(KEYINPUT110), .ZN(n680) );
  XNOR2_X1 U756 ( .A(n680), .B(n679), .ZN(G42) );
  AND2_X1 U757 ( .A1(KEYINPUT2), .A2(KEYINPUT78), .ZN(n682) );
  NAND2_X1 U758 ( .A1(n681), .A2(n682), .ZN(n724) );
  XNOR2_X1 U759 ( .A(n681), .B(KEYINPUT78), .ZN(n683) );
  NOR2_X1 U760 ( .A1(n683), .A2(KEYINPUT2), .ZN(n722) );
  NOR2_X1 U761 ( .A1(n687), .A2(n686), .ZN(n691) );
  NOR2_X1 U762 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U763 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U764 ( .A(n692), .B(KEYINPUT114), .ZN(n693) );
  NOR2_X1 U765 ( .A1(n716), .A2(n693), .ZN(n694) );
  XNOR2_X1 U766 ( .A(KEYINPUT115), .B(n694), .ZN(n710) );
  XNOR2_X1 U767 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n695) );
  XNOR2_X1 U768 ( .A(n695), .B(KEYINPUT51), .ZN(n706) );
  NAND2_X1 U769 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U770 ( .A(KEYINPUT49), .B(n698), .Z(n699) );
  NAND2_X1 U771 ( .A1(n700), .A2(n699), .ZN(n703) );
  NOR2_X1 U772 ( .A1(n568), .A2(n378), .ZN(n701) );
  XNOR2_X1 U773 ( .A(n701), .B(KEYINPUT50), .ZN(n702) );
  NOR2_X1 U774 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U775 ( .A(n706), .B(n705), .Z(n707) );
  NAND2_X1 U776 ( .A1(n715), .A2(n707), .ZN(n708) );
  XOR2_X1 U777 ( .A(KEYINPUT113), .B(n708), .Z(n709) );
  NAND2_X1 U778 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U779 ( .A(n711), .B(KEYINPUT116), .ZN(n712) );
  XNOR2_X1 U780 ( .A(KEYINPUT52), .B(n712), .ZN(n714) );
  NAND2_X1 U781 ( .A1(n714), .A2(n713), .ZN(n720) );
  INV_X1 U782 ( .A(n715), .ZN(n717) );
  NOR2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U784 ( .A1(G953), .A2(n718), .ZN(n719) );
  NAND2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U786 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U787 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U788 ( .A(KEYINPUT53), .B(n725), .Z(G75) );
  XOR2_X1 U789 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n726) );
  XNOR2_X1 U790 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U791 ( .A(n731), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U792 ( .A(KEYINPUT59), .B(KEYINPUT118), .Z(n732) );
  XNOR2_X1 U793 ( .A(n735), .B(n734), .ZN(n736) );
  INV_X1 U794 ( .A(KEYINPUT119), .ZN(n737) );
  NOR2_X1 U795 ( .A1(n744), .A2(n741), .ZN(G63) );
  XNOR2_X1 U796 ( .A(n743), .B(n742), .ZN(n745) );
  NAND2_X1 U797 ( .A1(n767), .A2(n746), .ZN(n750) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n747) );
  XNOR2_X1 U799 ( .A(KEYINPUT61), .B(n747), .ZN(n748) );
  NAND2_X1 U800 ( .A1(n748), .A2(G898), .ZN(n749) );
  NAND2_X1 U801 ( .A1(n750), .A2(n749), .ZN(n757) );
  XOR2_X1 U802 ( .A(n751), .B(n752), .Z(n753) );
  NOR2_X1 U803 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U804 ( .A(KEYINPUT121), .B(n755), .Z(n756) );
  XNOR2_X1 U805 ( .A(n757), .B(n756), .ZN(G69) );
  XNOR2_X1 U806 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n758) );
  XNOR2_X1 U807 ( .A(n759), .B(n758), .ZN(n760) );
  XNOR2_X1 U808 ( .A(n396), .B(n760), .ZN(n765) );
  XNOR2_X1 U809 ( .A(G227), .B(n765), .ZN(n761) );
  NAND2_X1 U810 ( .A1(n761), .A2(G900), .ZN(n762) );
  XOR2_X1 U811 ( .A(KEYINPUT124), .B(n762), .Z(n763) );
  NOR2_X1 U812 ( .A1(n767), .A2(n763), .ZN(n764) );
  XNOR2_X1 U813 ( .A(n764), .B(KEYINPUT125), .ZN(n770) );
  XOR2_X1 U814 ( .A(n766), .B(n765), .Z(n768) );
  NAND2_X1 U815 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U816 ( .A1(n770), .A2(n769), .ZN(G72) );
  XOR2_X1 U817 ( .A(G119), .B(KEYINPUT126), .Z(n771) );
  XNOR2_X1 U818 ( .A(n772), .B(n771), .ZN(G21) );
  XOR2_X1 U819 ( .A(n367), .B(G122), .Z(G24) );
  XNOR2_X1 U820 ( .A(n774), .B(G137), .ZN(G39) );
endmodule

