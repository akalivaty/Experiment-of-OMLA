//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n211, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1376, new_n1377;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(KEYINPUT64), .A3(G50), .ZN(new_n204));
  INV_X1    g0004(.A(KEYINPUT64), .ZN(new_n205));
  NOR2_X1   g0005(.A1(G58), .A2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  AOI21_X1  g0007(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NOR3_X1   g0008(.A1(new_n204), .A2(G77), .A3(new_n208), .ZN(G353));
  NOR2_X1   g0009(.A1(G97), .A2(G107), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G87), .ZN(G355));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n219), .B(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n218), .B1(new_n225), .B2(KEYINPUT0), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT65), .B(G77), .Z(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT66), .B(G244), .Z(new_n228));
  AND2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G87), .A2(G250), .ZN(new_n233));
  NAND4_X1  g0033(.A1(new_n230), .A2(new_n231), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n220), .B1(new_n229), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT1), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n226), .B(new_n236), .C1(KEYINPUT0), .C2(new_n225), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT68), .B(G50), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G226), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n257), .B(new_n260), .C1(G232), .C2(new_n259), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G97), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n256), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n264), .B(G274), .C1(G41), .C2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT69), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n270), .A2(KEYINPUT69), .A3(new_n264), .A4(G274), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT73), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n256), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G238), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n273), .B1(new_n256), .B2(new_n274), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n272), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT74), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(KEYINPUT74), .B(new_n272), .C1(new_n276), .C2(new_n277), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n263), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI211_X1 g0085(.A(new_n283), .B(new_n263), .C1(new_n280), .C2(new_n281), .ZN(new_n286));
  OAI21_X1  g0086(.A(G200), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n202), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT12), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT11), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n215), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n216), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(G77), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n295), .A2(new_n296), .B1(new_n216), .B2(G68), .ZN(new_n297));
  INV_X1    g0097(.A(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n216), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(new_n207), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n294), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n294), .B1(new_n264), .B2(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n291), .B1(new_n292), .B2(new_n301), .C1(new_n202), .C2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n301), .A2(new_n292), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n280), .A2(new_n281), .ZN(new_n307));
  INV_X1    g0107(.A(new_n263), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n284), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT13), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n309), .B(G190), .C1(new_n310), .C2(new_n282), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n287), .A2(new_n306), .A3(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n309), .B(G179), .C1(new_n310), .C2(new_n282), .ZN(new_n313));
  NAND2_X1  g0113(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(G169), .B1(new_n285), .B2(new_n286), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI221_X1 g0118(.A(G169), .B1(KEYINPUT76), .B2(KEYINPUT14), .C1(new_n285), .C2(new_n286), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n315), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n312), .B1(new_n320), .B2(new_n306), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT8), .B(G58), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n288), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n302), .B2(new_n322), .ZN(new_n324));
  INV_X1    g0124(.A(G159), .ZN(new_n325));
  OR3_X1    g0125(.A1(new_n299), .A2(KEYINPUT78), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT78), .B1(new_n299), .B2(new_n325), .ZN(new_n327));
  XNOR2_X1  g0127(.A(G58), .B(G68), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n326), .A2(new_n327), .B1(G20), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT7), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT3), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT77), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT77), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT3), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n298), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n330), .B(new_n216), .C1(new_n335), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G68), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n336), .B1(new_n340), .B2(new_n298), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n330), .B1(new_n341), .B2(new_n216), .ZN(new_n342));
  OAI211_X1 g0142(.A(KEYINPUT16), .B(new_n329), .C1(new_n339), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n294), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n216), .A2(KEYINPUT7), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n332), .A2(new_n334), .A3(new_n298), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n331), .A2(G33), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n336), .A2(new_n347), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT7), .B1(new_n349), .B2(new_n216), .ZN(new_n350));
  OAI21_X1  g0150(.A(G68), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT16), .B1(new_n351), .B2(new_n329), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n324), .B1(new_n344), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT17), .ZN(new_n355));
  NOR2_X1   g0155(.A1(G223), .A2(G1698), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n258), .B2(G1698), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(new_n336), .C1(new_n298), .C2(new_n340), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G87), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n256), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n256), .A2(G232), .A3(new_n274), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT79), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT79), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n256), .A2(new_n274), .A3(new_n363), .A4(G232), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n272), .A3(new_n364), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n360), .A2(new_n365), .A3(G190), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT81), .ZN(new_n367));
  INV_X1    g0167(.A(new_n256), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n258), .A2(G1698), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(G223), .B2(G1698), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n335), .A2(new_n370), .A3(new_n337), .ZN(new_n371));
  INV_X1    g0171(.A(new_n359), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n362), .A2(new_n272), .A3(new_n364), .ZN(new_n374));
  INV_X1    g0174(.A(G190), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT81), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n360), .B2(new_n365), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n367), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n354), .A2(new_n355), .A3(new_n381), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n351), .A2(new_n329), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n343), .B(new_n294), .C1(new_n383), .C2(KEYINPUT16), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n380), .B1(new_n366), .B2(KEYINPUT81), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n376), .A2(new_n377), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n384), .B(new_n324), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT17), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n360), .A2(new_n365), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G179), .ZN(new_n391));
  INV_X1    g0191(.A(G169), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(new_n390), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT18), .B1(new_n353), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT80), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n353), .A2(KEYINPUT18), .A3(new_n393), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI211_X1 g0197(.A(KEYINPUT80), .B(KEYINPUT18), .C1(new_n353), .C2(new_n393), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n389), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n256), .A2(new_n274), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n272), .B1(new_n258), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n227), .A2(new_n349), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n259), .A2(G222), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT70), .B1(new_n349), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT70), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n257), .A2(new_n405), .A3(G222), .A4(new_n259), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n257), .A2(G223), .A3(G1698), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n402), .A2(new_n404), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n401), .B1(new_n408), .B2(new_n368), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n379), .ZN(new_n410));
  AOI211_X1 g0210(.A(new_n375), .B(new_n401), .C1(new_n368), .C2(new_n408), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n288), .A2(G50), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n302), .B2(G50), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(G150), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n322), .A2(new_n295), .B1(new_n416), .B2(new_n299), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT71), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT71), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n419), .B1(new_n416), .B2(new_n299), .C1(new_n322), .C2(new_n295), .ZN(new_n420));
  OAI21_X1  g0220(.A(G20), .B1(new_n204), .B2(new_n208), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n415), .B1(new_n422), .B2(new_n294), .ZN(new_n423));
  OR2_X1    g0223(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n424));
  NAND2_X1  g0224(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n423), .B2(new_n424), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n412), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT10), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT10), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n412), .B(new_n430), .C1(new_n426), .C2(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n409), .A2(G169), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n422), .A2(new_n294), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n414), .ZN(new_n435));
  INV_X1    g0235(.A(G179), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n409), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(G232), .A2(G1698), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n259), .A2(G238), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n257), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n368), .C1(G107), .C2(new_n257), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n228), .A2(new_n256), .A3(new_n274), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n442), .A2(new_n272), .A3(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n444), .A2(G169), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n436), .ZN(new_n446));
  INV_X1    g0246(.A(new_n227), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n302), .A2(G77), .B1(new_n447), .B2(new_n289), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n447), .A2(new_n216), .B1(new_n322), .B2(new_n299), .ZN(new_n449));
  INV_X1    g0249(.A(new_n295), .ZN(new_n450));
  XOR2_X1   g0250(.A(KEYINPUT15), .B(G87), .Z(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n293), .A2(new_n215), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n445), .A2(new_n446), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(G190), .B2(new_n444), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n379), .B2(new_n444), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n432), .A2(new_n438), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n321), .A2(new_n399), .A3(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n299), .A2(new_n296), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT6), .ZN(new_n461));
  INV_X1    g0261(.A(G97), .ZN(new_n462));
  INV_X1    g0262(.A(G107), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n461), .B1(new_n464), .B2(new_n210), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n463), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(G97), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT82), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT6), .A2(G97), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n467), .B1(new_n468), .B2(G107), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n465), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n460), .B1(new_n470), .B2(G20), .ZN(new_n471));
  OAI21_X1  g0271(.A(G107), .B1(new_n348), .B2(new_n350), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n294), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n288), .A2(G97), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n264), .A2(G33), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n453), .A2(new_n288), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n475), .B1(new_n477), .B2(G97), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G244), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G1698), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n336), .B(new_n481), .C1(new_n340), .C2(new_n298), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n336), .A2(new_n347), .A3(G250), .A4(G1698), .ZN(new_n485));
  AND2_X1   g0285(.A1(KEYINPUT4), .A2(G244), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n336), .A2(new_n347), .A3(new_n486), .A4(new_n259), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n256), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n268), .A2(KEYINPUT5), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT5), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G41), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n264), .A2(G45), .A3(G274), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g0296(.A(KEYINPUT5), .B(G41), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n269), .A2(G1), .ZN(new_n498));
  INV_X1    g0298(.A(new_n215), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n255), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n496), .B1(new_n500), .B2(G257), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n490), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n436), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n483), .B2(new_n482), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n501), .B1(new_n506), .B2(new_n256), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n392), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n479), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT83), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n490), .B2(new_n502), .ZN(new_n511));
  OAI211_X1 g0311(.A(KEYINPUT83), .B(new_n501), .C1(new_n506), .C2(new_n256), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n511), .A2(G200), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n478), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n473), .B2(new_n294), .ZN(new_n515));
  OAI211_X1 g0315(.A(G190), .B(new_n501), .C1(new_n506), .C2(new_n256), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(KEYINPUT84), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n511), .A2(new_n512), .A3(G200), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT84), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n519), .A2(new_n520), .A3(new_n515), .A4(new_n516), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n509), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(G87), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(G20), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT22), .B1(new_n257), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n463), .A2(KEYINPUT23), .A3(G20), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT23), .B1(new_n463), .B2(G20), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G116), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n526), .A2(new_n527), .B1(G20), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g0330(.A(KEYINPUT88), .B(KEYINPUT24), .Z(new_n531));
  NAND2_X1  g0331(.A1(new_n332), .A2(new_n334), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G33), .ZN(new_n533));
  AND2_X1   g0333(.A1(KEYINPUT22), .A2(G87), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n533), .A2(new_n216), .A3(new_n336), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n530), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n531), .B1(new_n530), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(KEYINPUT89), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT89), .ZN(new_n539));
  AOI211_X1 g0339(.A(new_n539), .B(new_n531), .C1(new_n530), .C2(new_n535), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n294), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n494), .A2(new_n256), .ZN(new_n542));
  INV_X1    g0342(.A(new_n498), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n256), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n224), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(G294), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n298), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G250), .A2(G1698), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n223), .B2(G1698), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n548), .B1(new_n341), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n545), .B1(new_n552), .B2(new_n368), .ZN(new_n553));
  INV_X1    g0353(.A(new_n495), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n497), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n379), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n550), .B(new_n336), .C1(new_n298), .C2(new_n340), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n256), .B1(new_n557), .B2(new_n548), .ZN(new_n558));
  NOR4_X1   g0358(.A1(new_n558), .A2(new_n375), .A3(new_n545), .A4(new_n496), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n289), .A2(new_n463), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT90), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT25), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n477), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(new_n463), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT90), .B1(new_n561), .B2(new_n563), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n561), .A2(new_n563), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n541), .A2(new_n560), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n451), .A2(new_n288), .ZN(new_n572));
  INV_X1    g0372(.A(new_n451), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n565), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n216), .B(new_n336), .C1(new_n340), .C2(new_n298), .ZN(new_n575));
  OAI21_X1  g0375(.A(KEYINPUT86), .B1(new_n575), .B2(new_n202), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n450), .A2(new_n577), .A3(G97), .ZN(new_n578));
  AOI21_X1  g0378(.A(G20), .B1(G33), .B2(G97), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n523), .A2(KEYINPUT85), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT85), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G87), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n579), .B1(new_n583), .B2(new_n210), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n578), .B1(new_n584), .B2(new_n577), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n337), .B1(new_n532), .B2(G33), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT86), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n216), .A4(G68), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n576), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  AOI211_X1 g0389(.A(new_n572), .B(new_n574), .C1(new_n589), .C2(new_n294), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n495), .B1(new_n544), .B2(new_n219), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n528), .ZN(new_n593));
  NOR2_X1   g0393(.A1(G238), .A2(G1698), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n480), .B2(G1698), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n593), .B1(new_n586), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n592), .B1(new_n596), .B2(new_n256), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n392), .ZN(new_n598));
  INV_X1    g0398(.A(new_n595), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n528), .B1(new_n341), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n591), .B1(new_n600), .B2(new_n368), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n436), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n589), .A2(new_n294), .ZN(new_n604));
  INV_X1    g0404(.A(new_n572), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n477), .A2(G87), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n597), .A2(G200), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n592), .B(G190), .C1(new_n596), .C2(new_n256), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI22_X1  g0410(.A1(new_n590), .A2(new_n603), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n571), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n500), .A2(G264), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n547), .B1(new_n586), .B2(new_n550), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n555), .B(new_n613), .C1(new_n614), .C2(new_n256), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n392), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n553), .A2(new_n436), .A3(new_n555), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n541), .B2(new_n570), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n488), .B(new_n216), .C1(G33), .C2(new_n462), .ZN(new_n620));
  INV_X1    g0420(.A(G116), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G20), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n620), .A2(KEYINPUT20), .A3(new_n294), .A4(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT87), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n293), .A2(new_n215), .B1(G20), .B2(new_n621), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n620), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n626), .A2(KEYINPUT87), .A3(new_n620), .A4(KEYINPUT20), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n625), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n288), .A2(G116), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n477), .B2(G116), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n496), .B1(new_n500), .B2(G270), .ZN(new_n635));
  INV_X1    g0435(.A(G303), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n257), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n224), .A2(G1698), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(G257), .B2(G1698), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n586), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n635), .B1(new_n641), .B2(new_n256), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n634), .A2(new_n642), .A3(G169), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT21), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n634), .A2(new_n642), .A3(KEYINPUT21), .A4(G169), .ZN(new_n646));
  OAI211_X1 g0446(.A(G270), .B(new_n256), .C1(new_n494), .C2(new_n543), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n555), .ZN(new_n648));
  OAI22_X1  g0448(.A1(new_n341), .A2(new_n639), .B1(new_n636), .B2(new_n257), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(new_n368), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n634), .A2(new_n650), .A3(G179), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n645), .A2(new_n646), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n650), .A2(new_n379), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n642), .A2(new_n375), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n653), .A2(new_n654), .A3(new_n634), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n619), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  AND4_X1   g0456(.A1(new_n459), .A2(new_n522), .A3(new_n612), .A4(new_n656), .ZN(G372));
  INV_X1    g0457(.A(new_n438), .ZN(new_n658));
  INV_X1    g0458(.A(new_n394), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n396), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n318), .A2(new_n319), .ZN(new_n661));
  INV_X1    g0461(.A(new_n315), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n306), .ZN(new_n664));
  INV_X1    g0464(.A(new_n455), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n663), .A2(new_n664), .B1(new_n312), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n389), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n660), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n658), .B1(new_n668), .B2(new_n432), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n646), .A2(new_n651), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n335), .A2(new_n639), .A3(new_n337), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n368), .B1(new_n671), .B2(new_n637), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n392), .B1(new_n672), .B2(new_n635), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT21), .B1(new_n673), .B2(new_n634), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT91), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT91), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n645), .A2(new_n676), .A3(new_n646), .A4(new_n651), .ZN(new_n677));
  INV_X1    g0477(.A(new_n570), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n530), .A2(new_n535), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n539), .B1(new_n679), .B2(new_n531), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n537), .A2(KEYINPUT89), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n536), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n678), .B1(new_n682), .B2(new_n294), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n675), .B(new_n677), .C1(new_n683), .C2(new_n618), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n522), .A2(new_n684), .A3(new_n612), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n604), .A2(new_n605), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n598), .B(new_n602), .C1(new_n686), .C2(new_n574), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n479), .A2(new_n504), .A3(new_n508), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n611), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n572), .B1(new_n589), .B2(new_n294), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(new_n606), .A3(new_n608), .A4(new_n609), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n509), .A2(new_n687), .A3(KEYINPUT26), .A4(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n688), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n685), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n459), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n669), .A2(new_n697), .ZN(G369));
  INV_X1    g0498(.A(G13), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G20), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT27), .B1(new_n701), .B2(G1), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT27), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n700), .A2(new_n703), .A3(new_n264), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(G213), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G343), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT92), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n634), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n655), .B1(new_n710), .B2(new_n652), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n675), .A2(new_n677), .A3(new_n634), .A4(new_n709), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(G330), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n541), .A2(new_n570), .ZN(new_n714));
  INV_X1    g0514(.A(new_n618), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n708), .B1(new_n541), .B2(new_n570), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n571), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n619), .A2(new_n708), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n716), .A2(new_n709), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n652), .A2(new_n708), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n723), .B1(new_n718), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n722), .A2(new_n726), .ZN(G399));
  INV_X1    g0527(.A(new_n583), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n728), .A2(G116), .A3(new_n211), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n222), .A2(G41), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(new_n731), .A3(G1), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n213), .B2(new_n731), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n522), .A2(new_n656), .A3(new_n612), .A4(new_n708), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n672), .A2(G179), .A3(new_n635), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n507), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT93), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n613), .B1(new_n614), .B2(new_n256), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n738), .B1(new_n597), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n601), .A2(new_n553), .A3(KEYINPUT93), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n737), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(KEYINPUT94), .B(KEYINPUT30), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n650), .A2(new_n601), .A3(G179), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT95), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n507), .A2(new_n746), .A3(new_n615), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(new_n507), .B2(new_n615), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n737), .A2(new_n740), .A3(KEYINPUT30), .A4(new_n741), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n744), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n709), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT31), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n735), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n708), .A2(new_n753), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n750), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n744), .A2(new_n749), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n758), .B1(new_n759), .B2(KEYINPUT96), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT96), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n744), .A2(new_n749), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n757), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(G330), .B1(new_n755), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n652), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n716), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n522), .A2(new_n612), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n709), .B1(new_n767), .B2(new_n695), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n768), .A2(KEYINPUT29), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n709), .B1(new_n685), .B2(new_n695), .ZN(new_n770));
  XNOR2_X1  g0570(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n764), .B1(new_n769), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n734), .B1(new_n775), .B2(G1), .ZN(G364));
  NOR2_X1   g0576(.A1(new_n216), .A2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G179), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n325), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT32), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n436), .A2(new_n379), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n216), .A2(new_n375), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n436), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G50), .A2(new_n785), .B1(new_n788), .B2(G58), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n777), .A2(new_n786), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n781), .B(new_n789), .C1(new_n447), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n379), .A2(G179), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n777), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n463), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n783), .A2(new_n792), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n794), .B1(new_n728), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n216), .B1(new_n778), .B2(G190), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G97), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n782), .A2(new_n777), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n349), .B1(new_n802), .B2(G68), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n797), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n779), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G303), .A2(new_n796), .B1(new_n805), .B2(G329), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n785), .A2(G326), .ZN(new_n807));
  XOR2_X1   g0607(.A(KEYINPUT33), .B(G317), .Z(new_n808));
  OAI211_X1 g0608(.A(new_n806), .B(new_n807), .C1(new_n801), .C2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n793), .ZN(new_n810));
  INV_X1    g0610(.A(new_n790), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G283), .A2(new_n810), .B1(new_n811), .B2(G311), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n257), .B1(new_n788), .B2(G322), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(new_n546), .C2(new_n798), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n791), .A2(new_n804), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n499), .B1(new_n216), .B2(G169), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT98), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(KEYINPUT98), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G13), .A2(G33), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(G20), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n586), .A2(new_n222), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(G45), .B2(new_n213), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n250), .B2(G45), .ZN(new_n827));
  INV_X1    g0627(.A(G355), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n257), .A2(new_n221), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n828), .A2(new_n829), .B1(G116), .B2(new_n221), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n824), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n264), .B1(new_n700), .B2(G45), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n730), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n820), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n711), .A2(new_n712), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n823), .ZN(new_n837));
  INV_X1    g0637(.A(new_n713), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(new_n834), .ZN(new_n839));
  INV_X1    g0639(.A(G330), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n837), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G396));
  NOR2_X1   g0643(.A1(new_n819), .A2(new_n821), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n834), .B1(new_n845), .B2(G77), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n810), .A2(G87), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n463), .B2(new_n795), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n257), .B(new_n848), .C1(G283), .C2(new_n802), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G294), .A2(new_n788), .B1(new_n811), .B2(G116), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n785), .A2(G303), .B1(new_n805), .B2(G311), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n849), .A2(new_n800), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(G143), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n853), .A2(new_n787), .B1(new_n801), .B2(new_n416), .ZN(new_n854));
  INV_X1    g0654(.A(G137), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n784), .A2(new_n855), .B1(new_n790), .B2(new_n325), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n857), .A2(KEYINPUT34), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n795), .A2(new_n207), .B1(new_n793), .B2(new_n202), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(G132), .B2(new_n805), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n341), .B1(G58), .B2(new_n799), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n860), .B(new_n861), .C1(new_n857), .C2(KEYINPUT34), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n852), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n846), .B1(new_n863), .B2(new_n819), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n709), .A2(new_n454), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n665), .B1(new_n457), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n665), .A2(new_n708), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n864), .B1(new_n869), .B2(new_n822), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n770), .B(new_n869), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n834), .B1(new_n871), .B2(new_n764), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n871), .A2(new_n764), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(G384));
  OAI211_X1 g0675(.A(G116), .B(new_n217), .C1(new_n470), .C2(KEYINPUT35), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT99), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n470), .A2(KEYINPUT35), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n877), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n881), .B(KEYINPUT36), .Z(new_n882));
  OAI211_X1 g0682(.A(new_n214), .B(new_n227), .C1(new_n201), .C2(new_n202), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n207), .A2(G68), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n264), .B(G13), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT101), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n751), .A2(KEYINPUT101), .A3(KEYINPUT31), .A4(new_n709), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n754), .A3(new_n735), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n459), .A3(G330), .ZN(new_n893));
  INV_X1    g0693(.A(new_n866), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n867), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n708), .A2(new_n306), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n312), .B(new_n897), .C1(new_n320), .C2(new_n306), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n663), .A2(new_n896), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n391), .B(new_n705), .C1(new_n392), .C2(new_n390), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n353), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n903), .A2(new_n387), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT7), .B1(new_n586), .B2(G20), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(G68), .A3(new_n338), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT16), .B1(new_n909), .B2(new_n329), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n324), .B1(new_n344), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n902), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n907), .B1(new_n912), .B2(new_n387), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n706), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n901), .B(new_n914), .C1(new_n399), .C2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n355), .B1(new_n354), .B2(new_n381), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n387), .A2(KEYINPUT17), .ZN(new_n919));
  INV_X1    g0719(.A(new_n396), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n918), .A2(new_n919), .B1(new_n920), .B2(new_n394), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n354), .A2(new_n705), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n905), .B1(new_n903), .B2(new_n387), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n906), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT38), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n892), .B(new_n900), .C1(new_n917), .C2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n892), .A2(new_n928), .A3(new_n900), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n396), .A2(new_n395), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n659), .ZN(new_n931));
  INV_X1    g0731(.A(new_n398), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n915), .B1(new_n933), .B2(new_n389), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n901), .B1(new_n934), .B2(new_n914), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n914), .B1(new_n399), .B2(new_n916), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT38), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI22_X1  g0738(.A1(KEYINPUT40), .A2(new_n927), .B1(new_n929), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n893), .B1(new_n939), .B2(new_n840), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n929), .A2(new_n938), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n926), .B1(KEYINPUT38), .B2(new_n936), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n892), .A2(new_n900), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT40), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n459), .A3(new_n892), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n768), .A2(KEYINPUT29), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n459), .B(new_n948), .C1(new_n770), .C2(new_n772), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n669), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n947), .B(new_n950), .Z(new_n951));
  AOI21_X1  g0751(.A(new_n868), .B1(new_n770), .B2(new_n869), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n898), .A2(new_n899), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n938), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n660), .B2(new_n706), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n663), .A2(new_n664), .A3(new_n708), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n399), .A2(new_n916), .ZN(new_n959));
  INV_X1    g0759(.A(new_n914), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT38), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT39), .B1(new_n961), .B2(new_n917), .ZN(new_n962));
  INV_X1    g0762(.A(new_n926), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT39), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n937), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n958), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n957), .A2(new_n966), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n951), .A2(new_n967), .B1(new_n264), .B2(new_n700), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n951), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n886), .B1(new_n968), .B2(new_n969), .ZN(G367));
  AOI21_X1  g0770(.A(new_n708), .B1(new_n692), .B2(new_n606), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(new_n611), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n823), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n245), .A2(new_n222), .A3(new_n586), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n824), .B1(new_n221), .B2(new_n573), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n834), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(KEYINPUT105), .B(G311), .Z(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n341), .B1(new_n462), .B2(new_n793), .C1(new_n978), .C2(new_n784), .ZN(new_n979));
  INV_X1    g0779(.A(G317), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n787), .A2(new_n636), .B1(new_n779), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(G283), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n801), .A2(new_n546), .B1(new_n790), .B2(new_n982), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n979), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n796), .A2(KEYINPUT46), .A3(G116), .ZN(new_n985));
  AOI21_X1  g0785(.A(KEYINPUT46), .B1(new_n796), .B2(G116), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(G107), .B2(new_n799), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n257), .B1(new_n447), .B2(new_n793), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G143), .B2(new_n785), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n787), .A2(new_n416), .B1(new_n798), .B2(new_n202), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT106), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(KEYINPUT106), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n801), .A2(new_n325), .B1(new_n790), .B2(new_n207), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(KEYINPUT107), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n990), .A2(new_n992), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n795), .A2(new_n201), .B1(new_n779), .B2(new_n855), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT108), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(KEYINPUT107), .B2(new_n994), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n988), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT47), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n819), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n976), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n973), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT45), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n714), .A2(new_n709), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n541), .A2(new_n560), .A3(new_n570), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n619), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n719), .B1(new_n1010), .B2(new_n724), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n709), .A2(new_n479), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n522), .A2(new_n1012), .B1(new_n509), .B2(new_n709), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1007), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n518), .A2(new_n521), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1015), .A2(new_n690), .A3(new_n1012), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n509), .A2(new_n709), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1018), .A2(new_n726), .A3(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n1021));
  NAND3_X1  g0821(.A1(new_n1011), .A2(new_n1013), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1021), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n1018), .B2(new_n726), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n722), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n1010), .A2(new_n723), .A3(new_n724), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n725), .B1(new_n718), .B2(new_n719), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n838), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n720), .A2(new_n724), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n718), .A2(new_n719), .A3(new_n725), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n713), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n764), .C1(new_n769), .C2(new_n773), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1026), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1020), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n721), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n774), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n730), .B(KEYINPUT41), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT104), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1034), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1042), .A2(new_n1037), .A3(new_n1025), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n775), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT104), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(new_n1045), .A3(new_n1039), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n833), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n722), .A2(new_n1013), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1027), .A2(new_n522), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT42), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n690), .B1(new_n1016), .B2(new_n716), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1049), .A2(KEYINPUT42), .B1(new_n708), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n972), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1053), .A2(KEYINPUT43), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1050), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT102), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1054), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1053), .A2(KEYINPUT43), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1048), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1056), .A2(new_n1048), .A3(new_n1060), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1006), .B1(new_n1047), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT109), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT109), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n1006), .C1(new_n1047), .C2(new_n1064), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1068), .ZN(G387));
  NOR2_X1   g0869(.A1(new_n1042), .A2(new_n731), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n775), .B2(new_n1033), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n825), .B1(new_n241), .B2(new_n269), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n729), .B2(new_n829), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n322), .A2(G50), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT50), .ZN(new_n1075));
  AOI21_X1  g0875(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n729), .A3(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1073), .A2(new_n1077), .B1(new_n463), .B2(new_n222), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n824), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n834), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT110), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n796), .A2(new_n227), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n416), .B2(new_n779), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT111), .Z(new_n1085));
  OAI22_X1  g0885(.A1(new_n573), .A2(new_n798), .B1(new_n207), .B2(new_n787), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT112), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n801), .A2(new_n322), .B1(new_n793), .B2(new_n462), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n784), .A2(new_n325), .B1(new_n790), .B2(new_n202), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1088), .A2(new_n1089), .A3(new_n341), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1085), .A2(new_n1087), .A3(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G116), .A2(new_n810), .B1(new_n805), .B2(G326), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G322), .A2(new_n785), .B1(new_n788), .B2(G317), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n636), .B2(new_n790), .C1(new_n801), .C2(new_n978), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT48), .Z(new_n1095));
  OAI22_X1  g0895(.A1(new_n795), .A2(new_n546), .B1(new_n798), .B2(new_n982), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n341), .B(new_n1092), .C1(new_n1097), .C2(KEYINPUT49), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1097), .A2(KEYINPUT49), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1091), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n819), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1082), .B(new_n1103), .C1(new_n720), .C2(new_n823), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n833), .B2(new_n1033), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1071), .A2(new_n1105), .ZN(G393));
  INV_X1    g0906(.A(KEYINPUT113), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1025), .A2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(new_n1037), .Z(new_n1109));
  OAI211_X1 g0909(.A(new_n730), .B(new_n1043), .C1(new_n1109), .C2(new_n1042), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G317), .A2(new_n785), .B1(new_n788), .B2(G311), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT52), .Z(new_n1112));
  AOI22_X1  g0912(.A1(G294), .A2(new_n811), .B1(new_n805), .B2(G322), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G283), .A2(new_n796), .B1(new_n802), .B2(G303), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n257), .B(new_n794), .C1(G116), .C2(new_n799), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n784), .A2(new_n416), .B1(new_n787), .B2(new_n325), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT51), .Z(new_n1118));
  OAI221_X1 g0918(.A(new_n847), .B1(new_n202), .B2(new_n795), .C1(new_n853), .C2(new_n779), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n798), .A2(new_n296), .ZN(new_n1120));
  OR4_X1    g0920(.A1(new_n341), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n801), .A2(new_n207), .B1(new_n790), .B2(new_n322), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT115), .Z(new_n1123));
  OAI21_X1  g0923(.A(new_n1116), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n819), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n825), .A2(new_n253), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n824), .B(new_n1126), .C1(new_n462), .C2(new_n221), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT114), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n834), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n1128), .B2(new_n1127), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n1013), .B2(new_n823), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n1109), .B2(new_n833), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1110), .A2(new_n1133), .ZN(G390));
  OAI21_X1  g0934(.A(new_n958), .B1(new_n952), .B2(new_n954), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n962), .A2(new_n1135), .A3(new_n965), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n763), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(new_n754), .A3(new_n735), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1138), .A2(G330), .A3(new_n869), .A4(new_n953), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n868), .B1(new_n768), .B2(new_n894), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n958), .B1(new_n917), .B2(new_n926), .C1(new_n954), .C2(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1136), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n892), .A2(G330), .A3(new_n900), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1136), .B2(new_n1141), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n669), .A2(new_n949), .A3(new_n893), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n768), .A2(new_n894), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n867), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n889), .A2(new_n890), .ZN(new_n1148));
  OAI211_X1 g0948(.A(G330), .B(new_n869), .C1(new_n1148), .C2(new_n755), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1147), .B1(new_n1149), .B2(new_n954), .ZN(new_n1150));
  OAI211_X1 g0950(.A(G330), .B(new_n869), .C1(new_n755), .C2(new_n763), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n954), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1143), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n952), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1139), .A2(new_n1150), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1142), .A2(new_n1144), .B1(new_n1145), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1136), .A2(new_n1141), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1143), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1149), .A2(new_n954), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1145), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1136), .A2(new_n1141), .A3(new_n1139), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1159), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1156), .A2(new_n1165), .A3(new_n730), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n962), .A2(new_n821), .A3(new_n965), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n730), .B(new_n833), .C1(new_n844), .C2(new_n322), .ZN(new_n1168));
  XOR2_X1   g0968(.A(KEYINPUT54), .B(G143), .Z(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n1170), .A2(new_n790), .B1(new_n855), .B2(new_n801), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G159), .B2(new_n799), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT117), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n795), .A2(new_n416), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT53), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n349), .B1(new_n788), .B2(G132), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n785), .A2(G128), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G50), .A2(new_n810), .B1(new_n805), .B2(G125), .ZN(new_n1179));
  AND4_X1   g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n349), .B1(new_n795), .B2(new_n523), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT118), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n784), .A2(new_n982), .B1(new_n787), .B2(new_n621), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n202), .A2(new_n793), .B1(new_n790), .B2(new_n462), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n801), .A2(new_n463), .B1(new_n779), .B2(new_n546), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1120), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1174), .A2(new_n1180), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1167), .B(new_n1168), .C1(new_n1003), .C2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT116), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n833), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1142), .A2(new_n1144), .A3(KEYINPUT116), .A4(new_n832), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1166), .B(new_n1188), .C1(new_n1191), .C2(new_n1192), .ZN(G378));
  NOR2_X1   g0993(.A1(new_n423), .A2(new_n705), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT55), .B1(new_n432), .B2(new_n438), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT55), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1196), .B(new_n658), .C1(new_n429), .C2(new_n431), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n431), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n435), .A2(KEYINPUT72), .A3(KEYINPUT9), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n430), .B1(new_n1203), .B2(new_n412), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n438), .B1(new_n1200), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1196), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1194), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n432), .A2(KEYINPUT55), .A3(new_n438), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1198), .A2(new_n1199), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1199), .B1(new_n1198), .B2(new_n1209), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n945), .B2(G330), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n840), .B(new_n1212), .C1(new_n941), .C2(new_n944), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n967), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1212), .B1(new_n939), .B2(new_n840), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n957), .A2(new_n966), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n945), .A2(G330), .A3(new_n1213), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1216), .A2(KEYINPUT121), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT121), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1217), .A2(new_n1219), .A3(new_n1218), .A4(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1165), .A2(new_n950), .A3(new_n893), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1221), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT57), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1216), .B2(new_n1220), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n731), .B1(new_n1228), .B2(new_n1224), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1221), .A2(new_n833), .A3(new_n1223), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1083), .B1(new_n201), .B2(new_n793), .C1(new_n982), .C2(new_n779), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1232), .A2(G41), .A3(new_n586), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT119), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n784), .A2(new_n621), .B1(new_n787), .B2(new_n463), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n573), .A2(new_n790), .B1(new_n462), .B2(new_n801), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(G68), .C2(new_n799), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(KEYINPUT58), .A3(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n341), .B2(new_n268), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G128), .A2(new_n788), .B1(new_n802), .B2(G132), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n796), .A2(new_n1169), .B1(new_n811), .B2(G137), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n785), .A2(G125), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n799), .A2(G150), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1246));
  AOI211_X1 g1046(.A(G33), .B(G41), .C1(new_n805), .C2(G124), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n325), .B2(new_n793), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1245), .B2(KEYINPUT59), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1240), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1238), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT58), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n819), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n730), .B(new_n833), .C1(new_n844), .C2(new_n207), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(new_n1213), .C2(new_n822), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1231), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1230), .A2(new_n1257), .ZN(G375));
  NOR2_X1   g1058(.A1(new_n1155), .A2(new_n832), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n954), .A2(new_n821), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n834), .B1(new_n845), .B2(G68), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G283), .A2(new_n788), .B1(new_n811), .B2(G107), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1262), .B1(new_n296), .B2(new_n793), .C1(new_n546), .C2(new_n784), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G116), .A2(new_n802), .B1(new_n805), .B2(G303), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n257), .B1(new_n796), .B2(G97), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n573), .C2(new_n798), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n341), .B1(G50), .B2(new_n799), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(G132), .A2(new_n785), .B1(new_n802), .B2(new_n1169), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G137), .A2(new_n788), .B1(new_n810), .B2(G58), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G159), .A2(new_n796), .B1(new_n805), .B2(G128), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n416), .B2(new_n790), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n1263), .A2(new_n1266), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1261), .B1(new_n1273), .B2(new_n819), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1259), .B1(new_n1260), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1163), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1155), .A2(new_n1145), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1039), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(G381));
  AOI21_X1  g1079(.A(new_n1256), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1280));
  INV_X1    g1080(.A(G378), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(G390), .ZN(new_n1283));
  INV_X1    g1083(.A(G384), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1071), .A2(new_n842), .A3(new_n1105), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1283), .A2(new_n1284), .A3(new_n1286), .ZN(new_n1287));
  OR4_X1    g1087(.A1(G387), .A2(new_n1282), .A3(G381), .A4(new_n1287), .ZN(G407));
  OAI211_X1 g1088(.A(G407), .B(G213), .C1(G343), .C2(new_n1282), .ZN(G409));
  INV_X1    g1089(.A(G213), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(G343), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT60), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1277), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1155), .A2(KEYINPUT60), .A3(new_n1145), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1293), .A2(new_n730), .A3(new_n1276), .A4(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(G384), .A3(new_n1275), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G384), .B1(new_n1295), .B2(new_n1275), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G2897), .B(new_n1291), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1298), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1291), .A2(G2897), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n1296), .A3(new_n1301), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1281), .B1(new_n1230), .B2(new_n1257), .ZN(new_n1304));
  OR2_X1    g1104(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1166), .A2(new_n1188), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1218), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n833), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1305), .A2(new_n1306), .A3(new_n1255), .A4(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1221), .A2(new_n1039), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  OAI22_X1  g1112(.A1(new_n1310), .A2(new_n1312), .B1(new_n1290), .B2(G343), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1303), .B1(new_n1304), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT122), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1006), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1045), .B1(new_n1044), .B2(new_n1039), .ZN(new_n1318));
  AOI211_X1 g1118(.A(KEYINPUT104), .B(new_n1040), .C1(new_n1043), .C2(new_n775), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n832), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1063), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1321), .A2(new_n1061), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1317), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1323), .A2(new_n1067), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1068), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1283), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n842), .B1(new_n1071), .B2(new_n1105), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1286), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT123), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1323), .A2(new_n1330), .A3(G390), .ZN(new_n1331));
  OAI21_X1  g1131(.A(KEYINPUT123), .B1(new_n1065), .B2(new_n1283), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1326), .A2(new_n1329), .A3(new_n1331), .A4(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1065), .A2(new_n1283), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1323), .A2(G390), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1328), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT61), .B1(new_n1333), .B2(new_n1336), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1303), .B(KEYINPUT122), .C1(new_n1304), .C2(new_n1313), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1316), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1309), .A2(new_n1255), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1340), .A2(G378), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1291), .B1(new_n1341), .B2(new_n1311), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1342), .B(new_n1343), .C1(new_n1280), .C2(new_n1281), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(KEYINPUT63), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(G375), .A2(G378), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT63), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1346), .A2(new_n1347), .A3(new_n1342), .A4(new_n1343), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1345), .A2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(KEYINPUT124), .B1(new_n1339), .B2(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1332), .A2(new_n1329), .A3(new_n1331), .ZN(new_n1351));
  AOI21_X1  g1151(.A(G390), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1336), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT61), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1355), .B1(new_n1315), .B2(new_n1314), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT124), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1345), .A2(new_n1348), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1356), .A2(new_n1357), .A3(new_n1358), .A4(new_n1338), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1350), .A2(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1353), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1344), .A2(KEYINPUT62), .ZN(new_n1362));
  OR2_X1    g1162(.A1(new_n1344), .A2(KEYINPUT62), .ZN(new_n1363));
  XNOR2_X1  g1163(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1346), .A2(new_n1342), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1364), .B1(new_n1365), .B2(new_n1303), .ZN(new_n1366));
  OAI211_X1 g1166(.A(new_n1362), .B(new_n1363), .C1(new_n1366), .C2(KEYINPUT126), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT126), .ZN(new_n1368));
  AOI211_X1 g1168(.A(new_n1368), .B(new_n1364), .C1(new_n1365), .C2(new_n1303), .ZN(new_n1369));
  OAI21_X1  g1169(.A(new_n1361), .B1(new_n1367), .B2(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1360), .A2(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1371), .A2(KEYINPUT127), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT127), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1360), .A2(new_n1370), .A3(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1372), .A2(new_n1374), .ZN(G405));
  NAND2_X1  g1175(.A1(new_n1346), .A2(new_n1282), .ZN(new_n1376));
  XNOR2_X1  g1176(.A(new_n1376), .B(new_n1343), .ZN(new_n1377));
  XNOR2_X1  g1177(.A(new_n1377), .B(new_n1353), .ZN(G402));
endmodule


