//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n460), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(G101), .A3(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n461), .A2(new_n462), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n460), .ZN(new_n475));
  MUX2_X1   g050(.A(G100), .B(G112), .S(G2105), .Z(new_n476));
  AOI22_X1  g051(.A1(new_n475), .A2(G124), .B1(G2104), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n474), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(G126), .ZN(new_n482));
  OR2_X1    g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  OAI21_X1  g061(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(KEYINPUT4), .A2(G138), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n483), .B2(new_n484), .ZN(new_n489));
  NAND2_X1  g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n460), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n487), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(KEYINPUT69), .A3(G543), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n500), .A2(new_n502), .B1(KEYINPUT5), .B2(new_n499), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n499), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n500), .A2(new_n502), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(new_n508), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n506), .A2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(new_n503), .A2(G89), .A3(new_n513), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n509), .A2(G51), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n518), .A2(new_n519), .A3(new_n520), .A4(new_n522), .ZN(G286));
  INV_X1    g098(.A(G286), .ZN(G168));
  AOI22_X1  g099(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n505), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n509), .A2(G52), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n514), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n526), .A2(new_n529), .ZN(G171));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n505), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n503), .A2(G81), .A3(new_n513), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n509), .A2(G43), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n531), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n503), .A2(G56), .ZN(new_n538));
  AND2_X1   g113(.A1(G68), .A2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(G651), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n534), .A2(new_n535), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT70), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(G188));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n514), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n503), .A2(KEYINPUT71), .A3(new_n513), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n551), .A2(G91), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n509), .A2(new_n556), .A3(G53), .ZN(new_n557));
  AND2_X1   g132(.A1(KEYINPUT6), .A2(G651), .ZN(new_n558));
  NOR2_X1   g133(.A1(KEYINPUT6), .A2(G651), .ZN(new_n559));
  OAI211_X1 g134(.A(G53), .B(G543), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n551), .A2(KEYINPUT72), .A3(G91), .A4(new_n552), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n503), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n505), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n555), .A2(new_n562), .A3(new_n563), .A4(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G166), .ZN(G303));
  AND2_X1   g143(.A1(new_n551), .A2(new_n552), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G87), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n503), .A2(G74), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n513), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n509), .A2(KEYINPUT73), .A3(G49), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n571), .A2(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n570), .A2(new_n577), .ZN(G288));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT76), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n509), .A2(new_n581), .A3(G48), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n569), .A2(G86), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n511), .A2(G61), .A3(new_n512), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT74), .B1(new_n503), .B2(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT75), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n591), .B(G651), .C1(new_n587), .C2(new_n588), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n583), .A2(new_n590), .A3(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n505), .ZN(new_n595));
  INV_X1    g170(.A(new_n514), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G85), .B1(G47), .B2(new_n509), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(G290));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(G301), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n509), .A2(G54), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n511), .A2(new_n512), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI211_X1 g179(.A(KEYINPUT77), .B(new_n602), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G651), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n503), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(KEYINPUT77), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n551), .A2(G92), .A3(new_n552), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n569), .A2(KEYINPUT10), .A3(G92), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n600), .B1(new_n614), .B2(new_n599), .ZN(G284));
  AOI21_X1  g190(.A(new_n600), .B1(new_n614), .B2(new_n599), .ZN(G321));
  NOR2_X1   g191(.A1(G286), .A2(new_n599), .ZN(new_n617));
  INV_X1    g192(.A(G299), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n599), .ZN(G297));
  AOI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(new_n599), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  AOI21_X1  g197(.A(new_n505), .B1(new_n607), .B2(KEYINPUT77), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n623), .A2(new_n626), .B1(G54), .B2(new_n509), .ZN(new_n627));
  INV_X1    g202(.A(new_n612), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n610), .A2(new_n611), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n627), .B(new_n621), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n630), .A2(new_n599), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n599), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g208(.A1(new_n468), .A2(new_n469), .ZN(new_n634));
  INV_X1    g209(.A(new_n474), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  MUX2_X1   g216(.A(G99), .B(G111), .S(G2105), .Z(new_n642));
  AOI22_X1  g217(.A1(new_n475), .A2(G123), .B1(G2104), .B2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT78), .ZN(new_n644));
  AND3_X1   g219(.A1(new_n478), .A2(new_n644), .A3(G135), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n644), .B1(new_n478), .B2(G135), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2096), .Z(new_n648));
  NAND3_X1  g223(.A1(new_n640), .A2(new_n641), .A3(new_n648), .ZN(G156));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT15), .B(G2435), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2427), .ZN(new_n653));
  INV_X1    g228(.A(G2430), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n654), .B2(new_n653), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G1341), .B(G1348), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n656), .A2(new_n663), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT80), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT17), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2084), .B(G2090), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n671), .B1(new_n668), .B2(new_n670), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n669), .B2(new_n670), .ZN(new_n674));
  INV_X1    g249(.A(new_n670), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n675), .A2(new_n671), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n672), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(G2096), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2100), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n684), .A2(new_n687), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT20), .Z(new_n691));
  AOI211_X1 g266(.A(new_n689), .B(new_n691), .C1(new_n684), .C2(new_n688), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G229));
  NOR2_X1   g274(.A1(G29), .A2(G33), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n635), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(new_n460), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT25), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n478), .A2(G139), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n700), .B1(new_n708), .B2(G29), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G2072), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n711), .A2(G32), .ZN(new_n712));
  AOI22_X1  g287(.A1(G129), .A2(new_n475), .B1(new_n478), .B2(G141), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT26), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G105), .B2(new_n634), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n712), .B1(new_n717), .B2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT27), .B(G1996), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n710), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G2084), .ZN(new_n721));
  NAND2_X1  g296(.A1(G160), .A2(G29), .ZN(new_n722));
  AND2_X1   g297(.A1(KEYINPUT24), .A2(G34), .ZN(new_n723));
  NOR2_X1   g298(.A1(KEYINPUT24), .A2(G34), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n711), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT88), .Z(new_n727));
  OAI21_X1  g302(.A(new_n720), .B1(new_n721), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT89), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n711), .A2(G35), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT91), .Z(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G162), .B2(new_n711), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT29), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G2090), .ZN(new_n734));
  NOR2_X1   g309(.A1(G27), .A2(G29), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G164), .B2(G29), .ZN(new_n736));
  INV_X1    g311(.A(G2078), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n711), .A2(G26), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT28), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n478), .A2(G140), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n475), .A2(G128), .ZN(new_n742));
  AND2_X1   g317(.A1(G116), .A2(G2105), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G104), .B2(new_n460), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n742), .C1(new_n467), .C2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT87), .B(G2067), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n738), .B(new_n748), .C1(new_n718), .C2(new_n719), .ZN(new_n749));
  INV_X1    g324(.A(G16), .ZN(new_n750));
  NOR2_X1   g325(.A1(G171), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G5), .B2(new_n750), .ZN(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n727), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G2084), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n734), .A2(new_n749), .A3(new_n756), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n729), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g333(.A1(KEYINPUT30), .A2(G28), .ZN(new_n759));
  NOR2_X1   g334(.A1(KEYINPUT30), .A2(G28), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n711), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT31), .B(G11), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n761), .B(new_n762), .C1(new_n647), .C2(new_n711), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n750), .A2(G21), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G168), .B2(new_n750), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n763), .B1(new_n765), .B2(G1966), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n766), .B1(G1966), .B2(new_n765), .C1(new_n752), .C2(new_n753), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT90), .ZN(new_n768));
  NOR2_X1   g343(.A1(G4), .A2(G16), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n614), .B2(G16), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT85), .B(G1348), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n750), .A2(G19), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n543), .B2(new_n750), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT86), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1341), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n750), .A2(G20), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT23), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n618), .B2(new_n750), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1956), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n758), .A2(new_n768), .A3(new_n772), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n750), .A2(G23), .ZN(new_n783));
  INV_X1    g358(.A(G288), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n750), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT33), .B(G1976), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G22), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G166), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1971), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(G6), .A2(G16), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G305), .B2(new_n750), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT84), .Z(new_n795));
  XOR2_X1   g370(.A(KEYINPUT32), .B(G1981), .Z(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n792), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT34), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G24), .B(G290), .S(G16), .Z(new_n802));
  XOR2_X1   g377(.A(KEYINPUT83), .B(G1986), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G25), .A2(G29), .ZN(new_n805));
  MUX2_X1   g380(.A(G95), .B(G107), .S(G2105), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G2104), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT81), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n475), .A2(G119), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n478), .A2(G131), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n805), .B1(new_n812), .B2(G29), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT35), .B(G1991), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT82), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n813), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n804), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n799), .B2(new_n800), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n801), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT36), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n801), .A2(new_n821), .A3(new_n818), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n782), .B1(new_n820), .B2(new_n822), .ZN(G311));
  NAND2_X1  g398(.A1(new_n820), .A2(new_n822), .ZN(new_n824));
  INV_X1    g399(.A(new_n782), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(G150));
  OAI21_X1  g401(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(new_n621), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  INV_X1    g405(.A(G67), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n603), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G651), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT92), .B(G93), .Z(new_n834));
  NAND3_X1  g409(.A1(new_n503), .A2(new_n513), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n509), .A2(G55), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n836), .B1(new_n835), .B2(new_n837), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n840), .A2(new_n537), .A3(new_n542), .ZN(new_n841));
  OAI221_X1 g416(.A(new_n833), .B1(new_n533), .B2(new_n536), .C1(new_n839), .C2(new_n838), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n829), .B(new_n843), .Z(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT94), .B(G860), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n847), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n840), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(G145));
  XNOR2_X1  g427(.A(new_n480), .B(G160), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n647), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n708), .A2(KEYINPUT95), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n717), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI22_X1  g432(.A1(G130), .A2(new_n475), .B1(new_n478), .B2(G142), .ZN(new_n858));
  NOR3_X1   g433(.A1(new_n460), .A2(KEYINPUT96), .A3(G118), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT96), .B1(new_n460), .B2(G118), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n860), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n858), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n637), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n812), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n812), .ZN(new_n866));
  XNOR2_X1  g441(.A(G164), .B(new_n745), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n863), .A2(new_n812), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n867), .B1(new_n870), .B2(new_n864), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n857), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n868), .B1(new_n865), .B2(new_n866), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n864), .A3(new_n867), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n856), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n854), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(G37), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n854), .A3(new_n875), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n878), .A2(KEYINPUT97), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(KEYINPUT97), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n877), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g458(.A(KEYINPUT98), .B(new_n877), .C1(new_n879), .C2(new_n880), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n883), .A2(KEYINPUT40), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT40), .B1(new_n883), .B2(new_n884), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(G395));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n843), .B(new_n630), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n614), .A2(new_n618), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n827), .A2(G299), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(KEYINPUT41), .A3(new_n891), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n889), .A2(new_n894), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n843), .A2(new_n621), .A3(new_n614), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n630), .A2(new_n842), .A3(new_n841), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n614), .A2(new_n618), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n827), .A2(G299), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n900), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n900), .B2(new_n903), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n897), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n896), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT41), .B1(new_n890), .B2(new_n891), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n895), .B1(new_n910), .B2(new_n889), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT42), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n906), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n900), .A2(new_n903), .A3(new_n904), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n894), .A2(new_n896), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT100), .B1(new_n916), .B2(new_n900), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n915), .A2(new_n917), .A3(new_n918), .A4(new_n897), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n592), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n585), .A2(new_n586), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n503), .A2(KEYINPUT74), .A3(G61), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n584), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n591), .B1(new_n924), .B2(G651), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(G166), .A3(new_n583), .ZN(new_n927));
  NAND2_X1  g502(.A1(G305), .A2(G303), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(G288), .B(G290), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n929), .A2(new_n932), .A3(new_n930), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n920), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n935), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n912), .A2(new_n919), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n599), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n840), .A2(G868), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n888), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n938), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n937), .B1(new_n912), .B2(new_n919), .ZN(new_n944));
  OAI21_X1  g519(.A(G868), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(KEYINPUT102), .A3(new_n940), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n942), .A2(new_n946), .ZN(G295));
  NOR2_X1   g522(.A1(new_n939), .A2(new_n941), .ZN(G331));
  NAND2_X1  g523(.A1(G171), .A2(G168), .ZN(new_n949));
  OAI21_X1  g524(.A(G286), .B1(new_n526), .B2(new_n529), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n842), .A3(new_n841), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n951), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n843), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT104), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n843), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n953), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n903), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n955), .A2(new_n961), .A3(new_n952), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n951), .A2(new_n841), .A3(KEYINPUT105), .A4(new_n842), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n960), .B1(new_n916), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n935), .A2(KEYINPUT108), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n967), .B(new_n931), .C1(new_n933), .C2(new_n934), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G37), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n965), .A2(new_n966), .A3(KEYINPUT109), .A4(new_n968), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n974), .B1(new_n964), .B2(new_n903), .ZN(new_n975));
  AOI211_X1 g550(.A(KEYINPUT106), .B(new_n892), .C1(new_n962), .C2(new_n963), .ZN(new_n976));
  OAI221_X1 g551(.A(new_n935), .B1(new_n916), .B2(new_n959), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n979));
  OAI22_X1  g554(.A1(new_n975), .A2(new_n976), .B1(new_n916), .B2(new_n959), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT107), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n982));
  OAI221_X1 g557(.A(new_n982), .B1(new_n916), .B2(new_n959), .C1(new_n975), .C2(new_n976), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n981), .A2(new_n983), .A3(new_n966), .A4(new_n968), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n977), .A2(new_n972), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n979), .A2(new_n987), .A3(KEYINPUT44), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n978), .A2(new_n986), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n984), .A2(new_n985), .A3(KEYINPUT43), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n992), .ZN(G397));
  AND2_X1   g568(.A1(KEYINPUT4), .A2(G138), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n461), .B2(new_n462), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n490), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n996), .A2(new_n460), .B1(new_n494), .B2(new_n493), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n997), .B2(new_n487), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT110), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n470), .A2(new_n471), .ZN(new_n1002));
  INV_X1    g577(.A(G125), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n483), .B2(new_n484), .ZN(new_n1004));
  INV_X1    g579(.A(new_n464), .ZN(new_n1005));
  OAI21_X1  g580(.A(G2105), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1006), .A3(G40), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT112), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n1009));
  NAND3_X1  g584(.A1(G160), .A2(new_n1009), .A3(G40), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1001), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G2067), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n745), .B(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1013), .B1(new_n717), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT126), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1012), .A2(G1996), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT46), .Z(new_n1021));
  AND3_X1   g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1019), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1023));
  OR2_X1    g598(.A1(G290), .A2(G1986), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1012), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT127), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT48), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n717), .B(G1996), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1016), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n812), .B(new_n814), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1029), .B1(new_n1012), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n1022), .A2(new_n1023), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n808), .A2(new_n811), .A3(new_n814), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n1012), .B2(new_n1031), .ZN(new_n1038));
  OR2_X1    g613(.A1(new_n745), .A2(G2067), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1040), .A2(KEYINPUT124), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1013), .B1(new_n1040), .B2(KEYINPUT124), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1043), .A2(KEYINPUT125), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(KEYINPUT125), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1036), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G166), .A2(new_n1047), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n1048), .A2(KEYINPUT55), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(KEYINPUT55), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1009), .B1(G160), .B2(G40), .ZN(new_n1051));
  AND4_X1   g626(.A1(new_n1009), .A2(new_n1002), .A3(G40), .A4(new_n1006), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  OAI22_X1  g628(.A1(new_n1051), .A2(new_n1052), .B1(new_n998), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT115), .ZN(new_n1055));
  INV_X1    g630(.A(G2090), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n998), .A2(new_n1053), .ZN(new_n1057));
  INV_X1    g632(.A(G1384), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n496), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT50), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1011), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1059), .A2(new_n1000), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n998), .A2(KEYINPUT45), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1011), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n790), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(KEYINPUT116), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G8), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT116), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1049), .B(new_n1050), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1976), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT52), .B1(G288), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1059), .B1(new_n1010), .B2(new_n1008), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(new_n1047), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1073), .B(new_n1075), .C1(new_n1072), .C2(G288), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1011), .A2(new_n998), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G8), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(G1976), .B2(new_n784), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1076), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n580), .A2(new_n582), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n596), .A2(G86), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT113), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1084), .A3(KEYINPUT113), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n590), .A2(new_n1087), .A3(new_n592), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G1981), .ZN(new_n1090));
  INV_X1    g665(.A(G1981), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n583), .A2(new_n590), .A3(new_n1091), .A4(new_n592), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1082), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT49), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1078), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1091), .B1(new_n1096), .B2(new_n926), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1092), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT114), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT49), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1081), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1010), .A2(new_n1008), .B1(new_n1059), .B2(KEYINPUT50), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1057), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1067), .B1(G2090), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n1105), .A3(G8), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1059), .A2(KEYINPUT45), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n998), .A2(new_n1000), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1107), .A2(new_n1108), .B1(new_n1010), .B2(new_n1008), .ZN(new_n1109));
  OAI22_X1  g684(.A1(new_n1103), .A2(G2084), .B1(new_n1109), .B2(G1966), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G8), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(G286), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1071), .A2(new_n1101), .A3(new_n1106), .A4(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT63), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1105), .B1(new_n1104), .B2(G8), .ZN(new_n1116));
  NOR4_X1   g691(.A1(new_n1116), .A2(new_n1111), .A3(new_n1114), .A4(G286), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(new_n1101), .A3(new_n1106), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1071), .A2(new_n1101), .A3(new_n1106), .ZN(new_n1120));
  NAND2_X1  g695(.A1(G286), .A2(G8), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT51), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1111), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(G8), .B(new_n1123), .C1(new_n1110), .C2(G286), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1110), .A2(G8), .A3(G286), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1125), .A2(KEYINPUT62), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(G1961), .B1(new_n1102), .B2(new_n1057), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1066), .B2(G2078), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1109), .A2(KEYINPUT53), .A3(new_n737), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1138), .A2(G171), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1120), .A2(new_n1132), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(new_n1072), .A3(new_n784), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1092), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1106), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1143), .A2(new_n1075), .B1(new_n1144), .B2(new_n1101), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1119), .A2(new_n1140), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n556), .B1(new_n509), .B2(G53), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n557), .A2(new_n561), .A3(KEYINPUT117), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n555), .A2(new_n563), .A3(new_n565), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT57), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT118), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1153), .A2(new_n1157), .A3(new_n1154), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n565), .A2(new_n563), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1159), .A2(KEYINPUT57), .A3(new_n562), .A4(new_n555), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1156), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1055), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1162));
  INV_X1    g737(.A(G1956), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(KEYINPUT56), .B(G2072), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT119), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1011), .A2(new_n1064), .A3(new_n1065), .A4(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1161), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1167), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1169), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1170), .A2(new_n1161), .ZN(new_n1171));
  INV_X1    g746(.A(G1348), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1103), .A2(new_n1172), .B1(new_n1074), .B2(new_n1014), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1173), .A2(new_n827), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1168), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(KEYINPUT58), .B(G1341), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1066), .A2(G1996), .B1(new_n1074), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n543), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT59), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1178), .B(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1157), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1102), .A2(new_n1061), .B1(new_n1053), .B2(new_n998), .ZN(new_n1185));
  AOI21_X1  g760(.A(G1956), .B1(new_n1185), .B2(new_n1055), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1186), .B2(new_n1169), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1181), .B1(new_n1187), .B2(new_n1168), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1180), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1161), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1191));
  OAI21_X1  g766(.A(KEYINPUT120), .B1(new_n1191), .B2(new_n1171), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(KEYINPUT61), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1190), .A2(new_n1193), .A3(KEYINPUT121), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n827), .B(KEYINPUT60), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1174), .A2(KEYINPUT60), .B1(new_n1195), .B2(new_n1173), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(KEYINPUT121), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1175), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  XOR2_X1   g774(.A(G171), .B(KEYINPUT54), .Z(new_n1200));
  INV_X1    g775(.A(new_n1001), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1002), .A2(KEYINPUT53), .A3(G40), .A4(new_n737), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1065), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n463), .A2(new_n464), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT123), .ZN(new_n1205));
  AOI211_X1 g780(.A(new_n1202), .B(new_n1203), .C1(G2105), .C2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g781(.A(new_n1200), .B(new_n1133), .C1(new_n1201), .C2(new_n1206), .ZN(new_n1207));
  AOI22_X1  g782(.A1(new_n1207), .A2(new_n1136), .B1(new_n1138), .B2(new_n1200), .ZN(new_n1208));
  AND3_X1   g783(.A1(new_n1120), .A2(new_n1128), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1146), .B1(new_n1199), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(G290), .A2(G1986), .ZN(new_n1211));
  NAND4_X1  g786(.A1(new_n1031), .A2(new_n1032), .A3(new_n1024), .A4(new_n1211), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1013), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1046), .B1(new_n1210), .B2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g789(.A1(G401), .A2(new_n458), .ZN(new_n1216));
  NAND3_X1  g790(.A1(new_n698), .A2(new_n681), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g791(.A(new_n1217), .B1(new_n883), .B2(new_n884), .ZN(new_n1218));
  AND3_X1   g792(.A1(new_n1218), .A2(new_n989), .A3(new_n990), .ZN(G308));
  NAND3_X1  g793(.A1(new_n1218), .A2(new_n989), .A3(new_n990), .ZN(G225));
endmodule


