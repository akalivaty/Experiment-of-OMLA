//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT88), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT89), .ZN(new_n209));
  NOR3_X1   g008(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n209), .B2(new_n210), .ZN(new_n212));
  NAND2_X1  g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n206), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n210), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n203), .B1(new_n217), .B2(new_n213), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT17), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n204), .B(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(new_n213), .A3(new_n212), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223));
  INV_X1    g022(.A(new_n218), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(G1gat), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  OAI221_X1 g029(.A(new_n229), .B1(KEYINPUT90), .B2(new_n230), .C1(G1gat), .C2(new_n227), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(KEYINPUT90), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n226), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n222), .A2(new_n224), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n233), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n236), .B(new_n233), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n238), .B(KEYINPUT13), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n235), .A2(KEYINPUT18), .A3(new_n237), .A4(new_n238), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n241), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT11), .B(G169gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G197gat), .ZN(new_n248));
  XOR2_X1   g047(.A(G113gat), .B(G141gat), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT12), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n241), .A2(new_n251), .A3(new_n244), .A4(new_n245), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G155gat), .A2(G162gat), .ZN(new_n257));
  INV_X1    g056(.A(G155gat), .ZN(new_n258));
  INV_X1    g057(.A(G162gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n257), .B1(new_n260), .B2(KEYINPUT2), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT80), .ZN(new_n262));
  INV_X1    g061(.A(G141gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(new_n263), .B2(G148gat), .ZN(new_n264));
  INV_X1    g063(.A(G148gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n265), .A2(KEYINPUT80), .A3(G141gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n265), .A2(G141gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n261), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT2), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n263), .A2(G148gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n270), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n260), .A2(new_n257), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G113gat), .B(G120gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT71), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n280));
  XNOR2_X1  g079(.A(G127gat), .B(G134gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n278), .A2(KEYINPUT71), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n281), .A2(KEYINPUT70), .ZN(new_n284));
  INV_X1    g083(.A(G134gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G127gat), .ZN(new_n286));
  OAI22_X1  g085(.A1(new_n278), .A2(KEYINPUT1), .B1(KEYINPUT70), .B2(new_n286), .ZN(new_n287));
  OAI22_X1  g086(.A1(new_n282), .A2(new_n283), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n277), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n288), .A2(new_n275), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT4), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n288), .A2(KEYINPUT4), .A3(new_n275), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n290), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OR3_X1    g096(.A1(new_n295), .A2(KEYINPUT5), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n288), .B(new_n275), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n297), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n291), .A2(new_n296), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT5), .B(new_n300), .C1(new_n295), .C2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G1gat), .B(G29gat), .Z(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT82), .ZN(new_n304));
  XNOR2_X1  g103(.A(G57gat), .B(G85gat), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n304), .B(new_n305), .Z(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n298), .A2(new_n302), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT6), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n308), .B1(new_n298), .B2(new_n302), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(G183gat), .A2(G190gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT68), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(KEYINPUT24), .ZN(new_n318));
  NAND2_X1  g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n319), .B2(new_n318), .ZN(new_n321));
  NOR2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT66), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n323), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n322), .B(KEYINPUT67), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n321), .B(new_n329), .C1(new_n326), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT25), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n316), .B1(new_n333), .B2(new_n319), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n333), .B2(new_n319), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT65), .B(G169gat), .ZN(new_n337));
  INV_X1    g136(.A(G176gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(KEYINPUT23), .A3(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n335), .A2(new_n329), .A3(new_n336), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n323), .A2(KEYINPUT26), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n324), .B(new_n341), .C1(new_n330), .C2(KEYINPUT26), .ZN(new_n342));
  XOR2_X1   g141(.A(KEYINPUT27), .B(G183gat), .Z(new_n343));
  OAI21_X1  g142(.A(KEYINPUT28), .B1(new_n343), .B2(G190gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT69), .ZN(new_n345));
  INV_X1    g144(.A(G183gat), .ZN(new_n346));
  OR3_X1    g145(.A1(new_n345), .A2(new_n346), .A3(KEYINPUT27), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348));
  INV_X1    g147(.A(G190gat), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT27), .B1(new_n345), .B2(new_n346), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n342), .A2(new_n319), .A3(new_n344), .A4(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n332), .A2(new_n340), .A3(new_n352), .ZN(new_n353));
  XOR2_X1   g152(.A(KEYINPUT77), .B(KEYINPUT29), .Z(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n315), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(new_n315), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n357), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G197gat), .B(G204gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT22), .ZN(new_n363));
  INV_X1    g162(.A(G211gat), .ZN(new_n364));
  INV_X1    g163(.A(G218gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(G211gat), .B(G218gat), .Z(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT75), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n367), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n368), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n374), .B(KEYINPUT76), .Z(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n353), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n359), .B1(new_n379), .B2(new_n315), .ZN(new_n380));
  INV_X1    g179(.A(new_n374), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383));
  INV_X1    g182(.A(G64gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G92gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n377), .A2(new_n382), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT38), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n361), .A2(new_n376), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT37), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n380), .A2(new_n381), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT37), .B1(new_n377), .B2(new_n382), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n390), .B(new_n387), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n314), .A2(new_n389), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n377), .A2(new_n382), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n392), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n377), .A2(KEYINPUT37), .A3(new_n382), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n388), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n398), .B1(new_n402), .B2(new_n390), .ZN(new_n403));
  INV_X1    g202(.A(new_n401), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n387), .B1(new_n404), .B2(new_n395), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(KEYINPUT87), .A3(KEYINPUT38), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n397), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n276), .A2(new_n354), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n374), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT83), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n367), .A2(new_n368), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n370), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT3), .B1(new_n414), .B2(new_n355), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(new_n274), .B2(new_n269), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n409), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n381), .A2(KEYINPUT29), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n275), .B1(new_n418), .B2(KEYINPUT3), .ZN(new_n419));
  INV_X1    g218(.A(new_n409), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n419), .B(new_n420), .C1(new_n375), .C2(new_n410), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(KEYINPUT85), .A2(G22gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G78gat), .B(G106gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT31), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(G50gat), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n417), .A2(new_n421), .A3(KEYINPUT85), .A4(G22gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT84), .ZN(new_n430));
  INV_X1    g229(.A(G22gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n422), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n427), .B1(KEYINPUT84), .B2(G22gat), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n417), .A2(new_n421), .A3(new_n430), .A4(new_n431), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n429), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n389), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n388), .B1(new_n377), .B2(new_n382), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n389), .A2(new_n438), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT79), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT79), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n389), .A2(new_n444), .A3(new_n438), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n312), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n295), .A2(new_n297), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n448), .B(KEYINPUT39), .C1(new_n297), .C2(new_n299), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT86), .B(KEYINPUT39), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n449), .B(new_n308), .C1(new_n448), .C2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(KEYINPUT40), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n446), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n408), .A2(new_n437), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n353), .A2(new_n288), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n455), .A2(KEYINPUT73), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(KEYINPUT73), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OR3_X1    g257(.A1(new_n353), .A2(KEYINPUT72), .A3(new_n288), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT72), .B1(new_n353), .B2(new_n288), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G227gat), .A2(G233gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT34), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n463), .B(KEYINPUT64), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n458), .A2(new_n466), .A3(new_n467), .A4(new_n461), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT32), .ZN(new_n470));
  INV_X1    g269(.A(new_n467), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n462), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G15gat), .B(G43gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(G71gat), .B(G99gat), .ZN(new_n475));
  XOR2_X1   g274(.A(new_n474), .B(new_n475), .Z(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n471), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(KEYINPUT32), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(new_n465), .A3(new_n468), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n473), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n480), .B1(new_n473), .B2(new_n482), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n473), .A2(new_n482), .ZN(new_n488));
  INV_X1    g287(.A(new_n480), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT36), .B1(new_n490), .B2(new_n483), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n441), .A2(new_n313), .A3(new_n443), .A4(new_n445), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n429), .A2(new_n436), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n454), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(new_n437), .A3(new_n483), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n497), .A2(KEYINPUT35), .A3(new_n493), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT35), .B1(new_n497), .B2(new_n493), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n256), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G127gat), .B(G155gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(G211gat), .ZN(new_n504));
  XOR2_X1   g303(.A(G71gat), .B(G78gat), .Z(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT9), .ZN(new_n507));
  INV_X1    g306(.A(G71gat), .ZN(new_n508));
  INV_X1    g307(.A(G78gat), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n384), .A2(G57gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT93), .ZN(new_n512));
  INV_X1    g311(.A(G57gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(G64gat), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n506), .B(new_n510), .C1(new_n512), .C2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n511), .B2(new_n514), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n513), .A2(G64gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n384), .A2(G57gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT91), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n510), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT92), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n521), .A2(new_n522), .A3(new_n505), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(new_n521), .B2(new_n505), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n515), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT21), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n527), .A2(new_n346), .A3(new_n234), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n346), .B1(new_n527), .B2(new_n234), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT95), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n234), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G183gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT95), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n527), .A2(new_n346), .A3(new_n234), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT94), .B(KEYINPUT21), .Z(new_n536));
  NOR2_X1   g335(.A1(new_n526), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n530), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n530), .B2(new_n535), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n504), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n530), .A2(new_n535), .ZN(new_n542));
  INV_X1    g341(.A(new_n537), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n504), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n538), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n547));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n547), .B(new_n548), .Z(new_n549));
  AND3_X1   g348(.A1(new_n541), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n549), .B1(new_n541), .B2(new_n546), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G85gat), .A2(G92gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT7), .ZN(new_n554));
  NAND2_X1  g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT96), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT96), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(G99gat), .A3(G106gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n558), .A3(KEYINPUT8), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT97), .ZN(new_n560));
  INV_X1    g359(.A(G85gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n386), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n560), .B1(new_n559), .B2(new_n562), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n554), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G99gat), .B(G106gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n566), .B(new_n554), .C1(new_n563), .C2(new_n564), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n568), .A2(KEYINPUT98), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT98), .B1(new_n568), .B2(new_n569), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n226), .A2(new_n572), .B1(KEYINPUT41), .B2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G190gat), .B(G218gat), .Z(new_n575));
  OAI21_X1  g374(.A(new_n236), .B1(new_n570), .B2(new_n571), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT99), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT99), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n574), .A2(new_n579), .A3(new_n575), .A4(new_n576), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT100), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n573), .A2(KEYINPUT41), .ZN(new_n582));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n575), .B1(new_n574), .B2(new_n576), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n578), .B2(new_n580), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  AOI221_X4 g389(.A(new_n587), .B1(KEYINPUT100), .B2(new_n584), .C1(new_n578), .C2(new_n580), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n552), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G230gat), .ZN(new_n595));
  INV_X1    g394(.A(G233gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n559), .A2(new_n562), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT97), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n566), .B1(new_n602), .B2(new_n554), .ZN(new_n603));
  INV_X1    g402(.A(new_n569), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n525), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n521), .A2(new_n505), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT92), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n521), .A2(new_n522), .A3(new_n505), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n609), .A2(new_n568), .A3(new_n569), .A4(new_n515), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n605), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n609), .A2(KEYINPUT10), .A3(new_n515), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n603), .B2(new_n604), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n568), .A2(KEYINPUT98), .A3(new_n569), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n598), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n605), .A2(new_n610), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(new_n598), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G148gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT102), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G120gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n620), .A2(new_n624), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OR3_X1    g427(.A1(new_n594), .A2(KEYINPUT103), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT103), .B1(new_n594), .B2(new_n628), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n502), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n314), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g434(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n228), .A2(new_n230), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n633), .A2(new_n446), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n446), .ZN(new_n641));
  OAI21_X1  g440(.A(G8gat), .B1(new_n632), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n639), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(new_n642), .A3(new_n643), .ZN(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n632), .A2(new_n645), .A3(new_n492), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n484), .A2(new_n485), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n645), .B1(new_n632), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n649), .A2(KEYINPUT104), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(KEYINPUT104), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(G1326gat));
  NOR2_X1   g451(.A1(new_n632), .A2(new_n437), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT43), .B(G22gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  INV_X1    g454(.A(new_n549), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n539), .A2(new_n540), .A3(new_n504), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n545), .B1(new_n544), .B2(new_n538), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n541), .A2(new_n546), .A3(new_n549), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n628), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n593), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n664), .A2(KEYINPUT105), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(KEYINPUT105), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n502), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n667), .A2(G29gat), .A3(new_n313), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT45), .Z(new_n669));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT35), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n484), .A2(new_n485), .A3(new_n494), .ZN(new_n672));
  INV_X1    g471(.A(new_n493), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n498), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n487), .A2(new_n491), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n494), .B1(new_n397), .B2(new_n407), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(new_n453), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n493), .A2(KEYINPUT106), .A3(new_n494), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT106), .B1(new_n493), .B2(new_n494), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n675), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n670), .B1(new_n682), .B2(new_n593), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n496), .A2(new_n501), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n588), .A2(new_n581), .A3(new_n585), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n591), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(KEYINPUT44), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n663), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n683), .A2(new_n687), .A3(new_n255), .A4(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G29gat), .B1(new_n689), .B2(new_n313), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n669), .A2(new_n690), .ZN(G1328gat));
  NOR3_X1   g490(.A1(new_n667), .A2(G36gat), .A3(new_n641), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G36gat), .B1(new_n689), .B2(new_n641), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(G1329gat));
  INV_X1    g495(.A(G43gat), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n689), .A2(new_n697), .A3(new_n492), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n667), .A2(new_n648), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(G43gat), .ZN(new_n700));
  OR3_X1    g499(.A1(new_n698), .A2(KEYINPUT47), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT47), .B1(new_n698), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(G1330gat));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705));
  INV_X1    g504(.A(G50gat), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n689), .A2(new_n706), .A3(new_n437), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n502), .A2(new_n494), .A3(new_n665), .A4(new_n666), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n706), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n704), .B(new_n705), .C1(new_n707), .C2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n454), .A2(new_n681), .A3(new_n492), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n593), .B1(new_n712), .B2(new_n501), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(KEYINPUT44), .ZN(new_n714));
  AOI211_X1 g513(.A(new_n670), .B(new_n593), .C1(new_n496), .C2(new_n501), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n714), .A2(new_n715), .A3(new_n663), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n716), .A2(G50gat), .A3(new_n255), .A4(new_n494), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n704), .A2(new_n705), .ZN(new_n718));
  NAND2_X1  g517(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .A4(new_n709), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n711), .A2(new_n720), .ZN(G1331gat));
  INV_X1    g520(.A(new_n682), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n594), .A2(new_n255), .A3(new_n662), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n313), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(new_n513), .ZN(G1332gat));
  NOR2_X1   g525(.A1(new_n724), .A2(new_n641), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  AND2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n727), .B2(new_n728), .ZN(G1333gat));
  OAI21_X1  g530(.A(new_n508), .B1(new_n724), .B2(new_n648), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n722), .A2(G71gat), .A3(new_n676), .A4(new_n723), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g534(.A1(new_n724), .A2(new_n437), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(new_n509), .ZN(G1335gat));
  NOR2_X1   g536(.A1(new_n552), .A2(new_n255), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n683), .A2(new_n687), .A3(new_n628), .A4(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n313), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n713), .A2(KEYINPUT51), .A3(new_n738), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT51), .B1(new_n713), .B2(new_n738), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n628), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n314), .A2(new_n561), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n740), .B1(new_n745), .B2(new_n746), .ZN(G1336gat));
  INV_X1    g546(.A(new_n738), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n714), .A2(new_n715), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n749), .A2(new_n750), .A3(new_n446), .A4(new_n628), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT111), .B1(new_n739), .B2(new_n641), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(new_n752), .A3(G92gat), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n446), .A2(new_n386), .A3(new_n628), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT109), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n743), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n753), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n739), .A2(new_n641), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n386), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n741), .B2(new_n742), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n742), .A2(new_n761), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n756), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT52), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n758), .A2(new_n765), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n739), .B2(new_n492), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n648), .A2(G99gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n745), .B2(new_n768), .ZN(G1338gat));
  OAI21_X1  g568(.A(G106gat), .B1(new_n739), .B2(new_n437), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n437), .A2(G106gat), .A3(new_n662), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n770), .B(new_n771), .C1(new_n743), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n762), .A2(new_n763), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n772), .B(KEYINPUT112), .Z(new_n776));
  NAND3_X1  g575(.A1(new_n749), .A2(new_n494), .A3(new_n628), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n775), .A2(new_n776), .B1(new_n777), .B2(G106gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n774), .B1(new_n778), .B2(new_n771), .ZN(G1339gat));
  NAND2_X1  g578(.A1(KEYINPUT117), .A2(G113gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n624), .B1(new_n618), .B2(KEYINPUT54), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT10), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n525), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n570), .B2(new_n571), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n605), .A2(new_n610), .A3(new_n611), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n785), .A2(new_n786), .A3(new_n597), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n597), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT114), .B1(new_n789), .B2(KEYINPUT54), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n785), .A2(new_n786), .A3(new_n597), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n618), .A2(KEYINPUT114), .A3(KEYINPUT54), .A4(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n782), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n625), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n618), .A2(KEYINPUT54), .A3(new_n791), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n792), .ZN(new_n800));
  AND4_X1   g599(.A1(KEYINPUT115), .A2(new_n800), .A3(KEYINPUT55), .A4(new_n782), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n781), .B1(new_n799), .B2(new_n792), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT115), .B1(new_n802), .B2(KEYINPUT55), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n796), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n796), .B(KEYINPUT116), .C1(new_n801), .C2(new_n803), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n255), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n238), .B1(new_n235), .B2(new_n237), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n242), .A2(new_n243), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n250), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n254), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n628), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n686), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n590), .A2(new_n592), .A3(new_n812), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n806), .A2(new_n807), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n661), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n686), .A2(new_n661), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n819), .A2(new_n820), .A3(new_n256), .A4(new_n662), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n552), .A2(new_n593), .A3(new_n256), .A4(new_n662), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT113), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n497), .B1(new_n818), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n314), .A3(new_n641), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n256), .ZN(new_n828));
  NOR2_X1   g627(.A1(KEYINPUT117), .A2(G113gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n780), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n828), .B2(new_n780), .ZN(G1340gat));
  XNOR2_X1  g630(.A(KEYINPUT118), .B(G120gat), .ZN(new_n832));
  NAND2_X1  g631(.A1(KEYINPUT118), .A2(G120gat), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n827), .A2(new_n662), .ZN(new_n834));
  MUX2_X1   g633(.A(new_n832), .B(new_n833), .S(new_n834), .Z(G1341gat));
  NOR2_X1   g634(.A1(new_n827), .A2(new_n661), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(G127gat), .Z(G1342gat));
  XOR2_X1   g636(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G134gat), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n827), .A2(new_n593), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n838), .A2(G134gat), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n841), .B(new_n842), .ZN(G1343gat));
  NOR2_X1   g642(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n437), .B1(new_n818), .B2(new_n825), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n676), .A2(new_n313), .A3(new_n446), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n845), .A2(new_n263), .A3(new_n255), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n818), .A2(new_n825), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT57), .B1(new_n850), .B2(new_n494), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n437), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n794), .A2(new_n854), .A3(new_n795), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT120), .B1(new_n802), .B2(KEYINPUT55), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n855), .A2(new_n856), .A3(new_n255), .A4(new_n626), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n801), .A2(new_n803), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n813), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n593), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n552), .B1(new_n860), .B2(new_n816), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n853), .B1(new_n861), .B2(new_n824), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT121), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n864), .B(new_n853), .C1(new_n861), .C2(new_n824), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n255), .B(new_n846), .C1(new_n851), .C2(new_n866), .ZN(new_n867));
  AOI211_X1 g666(.A(new_n844), .B(new_n849), .C1(G141gat), .C2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n844), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(G141gat), .ZN(new_n870));
  INV_X1    g669(.A(new_n849), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n868), .A2(new_n872), .ZN(G1344gat));
  AND2_X1   g672(.A1(new_n845), .A2(new_n846), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n265), .A3(new_n628), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n845), .A2(new_n852), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n629), .A2(new_n256), .A3(new_n630), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n815), .B(new_n796), .C1(new_n803), .C2(new_n801), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n552), .B1(new_n860), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n852), .B(new_n494), .C1(new_n878), .C2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n877), .A2(new_n628), .A3(new_n846), .A4(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n876), .B1(new_n882), .B2(G148gat), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n628), .B(new_n846), .C1(new_n851), .C2(new_n866), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n884), .A2(new_n876), .A3(G148gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n875), .B1(new_n883), .B2(new_n885), .ZN(G1345gat));
  OAI21_X1  g685(.A(new_n846), .B1(new_n851), .B2(new_n866), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(new_n258), .A3(new_n661), .ZN(new_n888));
  AOI21_X1  g687(.A(G155gat), .B1(new_n874), .B2(new_n552), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(G1346gat));
  OAI21_X1  g689(.A(G162gat), .B1(new_n887), .B2(new_n593), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n259), .A3(new_n686), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n641), .A2(new_n314), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n850), .A2(new_n672), .A3(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n826), .A2(KEYINPUT123), .A3(new_n894), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n897), .A2(new_n255), .A3(new_n337), .A4(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G169gat), .B1(new_n895), .B2(new_n256), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1348gat));
  NOR3_X1   g700(.A1(new_n895), .A2(new_n338), .A3(new_n662), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n897), .A2(new_n628), .A3(new_n898), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n338), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT124), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n903), .A2(new_n906), .A3(new_n338), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n902), .B1(new_n905), .B2(new_n907), .ZN(G1349gat));
  OAI21_X1  g707(.A(G183gat), .B1(new_n895), .B2(new_n661), .ZN(new_n909));
  INV_X1    g708(.A(new_n895), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n552), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n911), .B2(new_n343), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n686), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT61), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(G190gat), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n915), .A2(KEYINPUT61), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n897), .A2(new_n349), .A3(new_n686), .A4(new_n898), .ZN(new_n920));
  INV_X1    g719(.A(new_n918), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n914), .A2(G190gat), .A3(new_n921), .A4(new_n916), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(G1351gat));
  NAND2_X1  g722(.A1(new_n492), .A2(new_n894), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n881), .B(new_n925), .C1(new_n845), .C2(new_n852), .ZN(new_n926));
  OAI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n256), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n845), .A2(new_n925), .ZN(new_n928));
  OR3_X1    g727(.A1(new_n928), .A2(G197gat), .A3(new_n256), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT126), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n927), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1352gat));
  NOR3_X1   g733(.A1(new_n928), .A2(G204gat), .A3(new_n662), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT62), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n877), .A2(new_n628), .A3(new_n881), .ZN(new_n937));
  OAI21_X1  g736(.A(G204gat), .B1(new_n937), .B2(new_n924), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1353gat));
  OR2_X1    g738(.A1(new_n926), .A2(new_n661), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n940), .B2(G211gat), .ZN(new_n941));
  OAI211_X1 g740(.A(KEYINPUT63), .B(G211gat), .C1(new_n926), .C2(new_n661), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n552), .A2(new_n364), .ZN(new_n944));
  OAI22_X1  g743(.A1(new_n941), .A2(new_n943), .B1(new_n928), .B2(new_n944), .ZN(G1354gat));
  NAND4_X1  g744(.A1(new_n845), .A2(new_n365), .A3(new_n686), .A4(new_n925), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n926), .A2(KEYINPUT127), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n926), .A2(KEYINPUT127), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n947), .A2(new_n948), .A3(new_n593), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n949), .B2(new_n365), .ZN(G1355gat));
endmodule


