//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT88), .B(G469), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G137), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT11), .A3(G134), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n192), .A2(new_n194), .A3(new_n198), .A4(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT86), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  AOI21_X1  g019(.A(G128), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n201), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G143), .B(G146), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(new_n207), .A3(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n202), .A2(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n213), .B(KEYINPUT86), .C1(new_n210), .C2(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G104), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT82), .B(G107), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G101), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(G104), .B2(new_n216), .ZN(new_n222));
  INV_X1    g036(.A(G104), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT84), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT83), .B1(new_n216), .B2(G104), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT83), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n223), .A3(G107), .ZN(new_n229));
  AOI21_X1  g043(.A(G101), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n225), .A2(new_n226), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n226), .B1(new_n225), .B2(new_n230), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n215), .B(new_n220), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n203), .A2(new_n205), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n235), .A2(new_n236), .B1(KEYINPUT1), .B2(new_n212), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n211), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n216), .A2(KEYINPUT82), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G107), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n224), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G101), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n228), .B1(new_n223), .B2(G107), .ZN(new_n246));
  NOR3_X1   g060(.A1(new_n216), .A2(KEYINPUT83), .A3(G104), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT84), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n225), .A2(new_n226), .A3(new_n230), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n238), .B1(new_n251), .B2(new_n220), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n200), .B1(new_n234), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT12), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n249), .A2(new_n250), .B1(G101), .B2(new_n219), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n233), .B1(new_n256), .B2(new_n238), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT12), .A3(new_n200), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G140), .ZN(new_n260));
  INV_X1    g074(.A(G227), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(G953), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n260), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n227), .A2(new_n229), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n242), .A3(new_n243), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G101), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT0), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(new_n236), .ZN(new_n270));
  NOR2_X1   g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n235), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n210), .B1(new_n269), .B2(new_n236), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n267), .B1(new_n266), .B2(G101), .ZN(new_n277));
  OAI211_X1 g091(.A(KEYINPUT85), .B(new_n277), .C1(new_n231), .C2(new_n232), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT85), .B1(new_n251), .B2(new_n277), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n200), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT10), .ZN(new_n283));
  INV_X1    g097(.A(new_n238), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(new_n283), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n233), .A2(new_n283), .B1(new_n256), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n281), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n259), .A2(new_n264), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n277), .B1(new_n231), .B2(new_n232), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT85), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n275), .B1(new_n291), .B2(new_n278), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n233), .A2(new_n283), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n256), .A2(new_n285), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n292), .A2(new_n295), .A3(new_n200), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n282), .B1(new_n281), .B2(new_n286), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n263), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI211_X1 g112(.A(G902), .B(new_n189), .C1(new_n288), .C2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n257), .A2(KEYINPUT12), .A3(new_n200), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT12), .B1(new_n257), .B2(new_n200), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT87), .B1(new_n303), .B2(new_n296), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT87), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n287), .B(new_n305), .C1(new_n301), .C2(new_n302), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n264), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n287), .A2(new_n264), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(new_n297), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n300), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n299), .B1(new_n310), .B2(G469), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT9), .B(G234), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT80), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n300), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G221), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n315), .B(KEYINPUT81), .Z(new_n316));
  OAI21_X1  g130(.A(new_n187), .B1(new_n311), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n316), .ZN(new_n318));
  INV_X1    g132(.A(G469), .ZN(new_n319));
  INV_X1    g133(.A(new_n306), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n305), .B1(new_n259), .B2(new_n287), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n263), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n309), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n319), .B1(new_n324), .B2(new_n300), .ZN(new_n325));
  OAI211_X1 g139(.A(KEYINPUT89), .B(new_n318), .C1(new_n325), .C2(new_n299), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n317), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT2), .B(G113), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT64), .B(G119), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G116), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT65), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(G116), .ZN(new_n334));
  INV_X1    g148(.A(G116), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT65), .A3(G119), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n328), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n328), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n330), .A2(new_n339), .A3(new_n336), .A4(new_n334), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n191), .A2(G137), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n193), .A2(G134), .ZN(new_n343));
  OAI21_X1  g157(.A(G131), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n199), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(new_n237), .B2(new_n211), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n199), .A2(new_n197), .B1(new_n272), .B2(new_n273), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT30), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT30), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n200), .A2(new_n274), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n199), .A2(new_n344), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n238), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n349), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n341), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT68), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT67), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G237), .ZN(new_n359));
  INV_X1    g173(.A(G953), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G210), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n356), .B(KEYINPUT67), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n361), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT26), .B(G101), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n363), .A2(new_n365), .A3(new_n367), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n346), .A2(new_n347), .ZN(new_n372));
  INV_X1    g186(.A(new_n341), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n354), .A2(new_n355), .A3(new_n371), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT31), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n350), .A2(new_n352), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(new_n341), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT30), .B1(new_n346), .B2(new_n347), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n350), .A2(new_n352), .A3(new_n349), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n378), .B1(new_n381), .B2(new_n341), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT31), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n382), .A2(new_n355), .A3(new_n383), .A4(new_n371), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n369), .A2(new_n370), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT28), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n377), .A2(new_n341), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n386), .B1(new_n374), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT28), .B1(new_n372), .B2(new_n373), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n376), .A2(new_n384), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G472), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n300), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT32), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT70), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n391), .A2(KEYINPUT32), .A3(new_n392), .A4(new_n300), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n391), .A2(new_n392), .A3(new_n300), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n400));
  OR3_X1    g214(.A1(new_n388), .A2(new_n385), .A3(new_n389), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT69), .B1(new_n382), .B2(new_n371), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT69), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n373), .B1(new_n379), .B2(new_n380), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n385), .B(new_n404), .C1(new_n405), .C2(new_n378), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n401), .A2(new_n402), .A3(new_n403), .A4(new_n406), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n388), .A2(new_n385), .A3(new_n389), .ZN(new_n408));
  AOI21_X1  g222(.A(G902), .B1(new_n408), .B2(KEYINPUT29), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n398), .A2(new_n400), .B1(G472), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G217), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(G234), .B2(new_n300), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT74), .ZN(new_n415));
  INV_X1    g229(.A(G125), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(KEYINPUT74), .A2(G125), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n420), .A2(KEYINPUT16), .A3(G140), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT76), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT16), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT75), .ZN(new_n425));
  INV_X1    g239(.A(G140), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n425), .B1(G125), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n419), .B2(new_n426), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n417), .A2(new_n425), .A3(G140), .A4(new_n418), .ZN(new_n429));
  AOI211_X1 g243(.A(new_n423), .B(new_n424), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  AND2_X1   g244(.A1(KEYINPUT74), .A2(G125), .ZN(new_n431));
  NOR2_X1   g245(.A1(KEYINPUT74), .A2(G125), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n431), .A2(new_n432), .A3(new_n426), .ZN(new_n433));
  INV_X1    g247(.A(new_n427), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT76), .B1(new_n435), .B2(KEYINPUT16), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n422), .B1(new_n430), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n202), .ZN(new_n438));
  OAI211_X1 g252(.A(G146), .B(new_n422), .C1(new_n430), .C2(new_n436), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n236), .A2(G119), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT71), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n236), .A2(KEYINPUT71), .A3(G119), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n333), .A2(KEYINPUT64), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT64), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G119), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n448), .A3(G128), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT72), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n329), .A2(KEYINPUT72), .A3(G128), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n445), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT24), .B(G110), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT73), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT23), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n329), .B2(G128), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n236), .A2(KEYINPUT23), .A3(G119), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n449), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G110), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n440), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n426), .A2(G125), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n416), .A2(G140), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n202), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  XOR2_X1   g282(.A(KEYINPUT77), .B(G110), .Z(new_n469));
  NAND4_X1  g283(.A1(new_n458), .A2(new_n449), .A3(new_n459), .A4(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n453), .B2(new_n455), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n468), .B1(new_n471), .B2(KEYINPUT78), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT78), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n470), .B(new_n473), .C1(new_n453), .C2(new_n455), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n439), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT22), .B(G137), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n360), .A2(G221), .A3(G234), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n464), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n478), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n462), .B1(new_n438), .B2(new_n439), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n472), .A2(new_n474), .A3(new_n439), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n479), .A2(new_n483), .A3(new_n300), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT25), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n479), .A2(new_n483), .A3(KEYINPUT25), .A4(new_n300), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n414), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n479), .A2(new_n483), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n413), .A2(G902), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(KEYINPUT79), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n411), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G214), .B1(G237), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n272), .A2(new_n273), .A3(new_n419), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n238), .B2(new_n419), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n360), .A2(G224), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n341), .A2(new_n268), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n279), .B2(new_n280), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n251), .A2(new_n220), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT5), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n331), .A2(new_n506), .A3(new_n337), .ZN(new_n507));
  OAI21_X1  g321(.A(G113), .B1(new_n330), .B2(KEYINPUT5), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n340), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(G110), .B(G122), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT91), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT91), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n504), .A2(new_n514), .A3(new_n510), .A4(new_n511), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n513), .A2(KEYINPUT6), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT6), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n505), .A2(new_n509), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n291), .A2(new_n278), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n521), .B1(new_n522), .B2(new_n503), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n520), .B1(new_n523), .B2(new_n511), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n504), .A2(new_n510), .ZN(new_n525));
  INV_X1    g339(.A(new_n511), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n519), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n502), .B1(new_n516), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G210), .B1(G237), .B2(G902), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n513), .A2(new_n515), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT93), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n498), .A2(new_n532), .B1(KEYINPUT7), .B2(new_n500), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(new_n499), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n505), .B(new_n509), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT92), .B(KEYINPUT8), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n511), .B(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n534), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(G902), .B1(new_n531), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n529), .A2(new_n530), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n530), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n519), .B1(new_n525), .B2(new_n526), .ZN(new_n542));
  AOI211_X1 g356(.A(new_n511), .B(new_n520), .C1(new_n504), .C2(new_n510), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n513), .A2(KEYINPUT6), .A3(new_n515), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n501), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n514), .B1(new_n523), .B2(new_n511), .ZN(new_n547));
  INV_X1    g361(.A(new_n515), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n538), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n300), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n541), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n497), .B1(new_n540), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n359), .A2(new_n360), .A3(G214), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(KEYINPUT94), .B2(new_n204), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT94), .B(G143), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G131), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n554), .B(new_n198), .C1(new_n553), .C2(new_n555), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n559), .B1(new_n561), .B2(new_n558), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n438), .A2(new_n439), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(G113), .B(G122), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(new_n223), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n467), .B1(new_n435), .B2(new_n202), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT95), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g384(.A1(KEYINPUT18), .A2(G131), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n556), .B(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n563), .A2(new_n565), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n565), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n557), .A2(new_n560), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT19), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n465), .A2(new_n466), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n581), .B(new_n582), .C1(new_n435), .C2(new_n578), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n577), .B1(new_n583), .B2(G146), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n435), .A2(KEYINPUT16), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n423), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n435), .A2(KEYINPUT76), .A3(KEYINPUT16), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n421), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n584), .B1(new_n588), .B2(G146), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n572), .B1(new_n568), .B2(new_n569), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n576), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n575), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT20), .ZN(new_n593));
  NOR2_X1   g407(.A1(G475), .A2(G902), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n592), .A2(KEYINPUT97), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n575), .A2(new_n598), .A3(new_n591), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n594), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n596), .B1(new_n600), .B2(KEYINPUT20), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n563), .A2(new_n574), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n576), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n575), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n300), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G475), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n204), .A2(G128), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT13), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n236), .A2(G143), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n609), .A2(new_n610), .ZN(new_n614));
  OAI21_X1  g428(.A(G134), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n609), .A2(new_n612), .A3(new_n191), .ZN(new_n616));
  XNOR2_X1  g430(.A(G116), .B(G122), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n218), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n218), .A2(new_n617), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n615), .B(new_n616), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT14), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n335), .A2(KEYINPUT14), .A3(G122), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(G107), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT98), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n609), .A2(new_n612), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G134), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n627), .A2(new_n616), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n628), .A2(new_n619), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n620), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n313), .A2(G217), .A3(new_n360), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  AOI21_X1  g447(.A(G902), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(G478), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(KEYINPUT15), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(KEYINPUT15), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n635), .A2(new_n641), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n608), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(G234), .A2(G237), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n646), .A2(G952), .A3(new_n360), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n646), .A2(G902), .A3(G953), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT21), .B(G898), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n327), .A2(new_n495), .A3(new_n552), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G101), .ZN(G3));
  NAND2_X1  g467(.A1(KEYINPUT100), .A2(G472), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n391), .A2(new_n300), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n391), .B2(new_n300), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n494), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n327), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n630), .A2(new_n661), .ZN(new_n662));
  AND4_X1   g476(.A1(KEYINPUT33), .A2(new_n632), .A3(new_n633), .A4(new_n662), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n632), .A2(new_n633), .B1(KEYINPUT33), .B2(new_n662), .ZN(new_n664));
  OAI21_X1  g478(.A(G478), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n636), .A2(new_n300), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n634), .B2(new_n636), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n575), .A2(new_n598), .A3(new_n591), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n598), .B1(new_n575), .B2(new_n591), .ZN(new_n670));
  INV_X1    g484(.A(new_n594), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n595), .B1(new_n672), .B2(new_n593), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n668), .B1(new_n673), .B2(new_n606), .ZN(new_n674));
  INV_X1    g488(.A(new_n650), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n552), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n660), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT34), .B(G104), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G6));
  NAND2_X1  g494(.A1(new_n672), .A2(new_n593), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n600), .A2(KEYINPUT20), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n607), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n644), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n660), .A2(new_n677), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT35), .B(G107), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G9));
  NOR2_X1   g502(.A1(new_n480), .A2(KEYINPUT36), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n464), .A2(new_n475), .A3(new_n689), .ZN(new_n690));
  OAI22_X1  g504(.A1(new_n481), .A2(new_n482), .B1(KEYINPUT36), .B2(new_n480), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n491), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n488), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n658), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n327), .A2(new_n552), .A3(new_n651), .A4(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT37), .B(G110), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G12));
  INV_X1    g513(.A(new_n647), .ZN(new_n700));
  INV_X1    g514(.A(new_n648), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n700), .B1(new_n701), .B2(G900), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n683), .A2(new_n684), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n411), .A2(new_n695), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n327), .A2(new_n552), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G128), .ZN(G30));
  NAND2_X1  g520(.A1(new_n540), .A2(new_n551), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT38), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n382), .A2(new_n371), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n374), .A2(new_n387), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n709), .B(new_n710), .C1(new_n371), .C2(new_n711), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n385), .A2(new_n405), .A3(new_n378), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n371), .B1(new_n374), .B2(new_n387), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT102), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n712), .A2(new_n715), .A3(new_n300), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G472), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n716), .A2(KEYINPUT103), .A3(G472), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n400), .B2(new_n398), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n684), .B(new_n496), .C1(new_n601), .C2(new_n607), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n486), .A2(new_n487), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n413), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n693), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n708), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n702), .B(KEYINPUT39), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n317), .B2(new_n326), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT40), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n204), .ZN(G45));
  INV_X1    g551(.A(new_n668), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n738), .B(new_n702), .C1(new_n601), .C2(new_n607), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n327), .A2(new_n552), .A3(new_n704), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G146), .ZN(G48));
  INV_X1    g556(.A(new_n299), .ZN(new_n743));
  AOI21_X1  g557(.A(G902), .B1(new_n288), .B2(new_n298), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n743), .B(new_n315), .C1(new_n744), .C2(new_n319), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n411), .A2(new_n745), .A3(new_n494), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n677), .A3(new_n674), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT41), .B(G113), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G15));
  NAND3_X1  g563(.A1(new_n746), .A2(new_n677), .A3(new_n685), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G116), .ZN(G18));
  NOR2_X1   g565(.A1(new_n744), .A2(new_n319), .ZN(new_n752));
  INV_X1    g566(.A(new_n315), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n752), .A2(new_n299), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n707), .A2(new_n754), .A3(new_n496), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n755), .A2(new_n650), .A3(new_n645), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n704), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G119), .ZN(G21));
  AOI21_X1  g572(.A(new_n392), .B1(new_n391), .B2(new_n300), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n399), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n493), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n761), .A2(new_n745), .A3(new_n650), .ZN(new_n762));
  INV_X1    g576(.A(new_n707), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n724), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G122), .ZN(G24));
  INV_X1    g580(.A(KEYINPUT104), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n391), .A2(new_n300), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(G472), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n393), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n726), .B2(new_n693), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n674), .A3(new_n702), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n767), .B1(new_n772), .B2(new_n755), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n760), .B1(new_n488), .B2(new_n694), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n739), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(KEYINPUT104), .A3(new_n552), .A4(new_n754), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G125), .ZN(G27));
  NAND3_X1  g592(.A1(new_n540), .A2(new_n551), .A3(new_n496), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT106), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n540), .A2(new_n551), .A3(KEYINPUT106), .A4(new_n496), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT105), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n311), .B2(new_n753), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT105), .B(new_n315), .C1(new_n325), .C2(new_n299), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n410), .A2(G472), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n395), .A3(new_n397), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n493), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT42), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n790), .A2(new_n739), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n783), .A2(new_n787), .A3(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n783), .A2(new_n787), .A3(new_n495), .A4(new_n740), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT107), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G131), .ZN(G33));
  NAND4_X1  g614(.A1(new_n783), .A2(new_n787), .A3(new_n495), .A4(new_n703), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  NAND2_X1  g616(.A1(new_n781), .A2(new_n782), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n673), .A2(new_n606), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT43), .B1(new_n804), .B2(new_n668), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT43), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n608), .A2(new_n806), .A3(new_n738), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT108), .B1(new_n727), .B2(new_n658), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n695), .A2(new_n809), .A3(new_n657), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n805), .B(new_n807), .C1(new_n808), .C2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT44), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n803), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT45), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n307), .B2(new_n309), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n322), .A2(KEYINPUT45), .A3(new_n323), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n816), .A3(G469), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n319), .A2(new_n300), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT46), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n818), .A2(new_n821), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n299), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n753), .B(new_n731), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n805), .A2(new_n807), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n810), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n809), .B1(new_n695), .B2(new_n657), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n827), .A2(new_n830), .A3(KEYINPUT44), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n813), .A2(new_n825), .A3(new_n831), .ZN(new_n832));
  XOR2_X1   g646(.A(KEYINPUT109), .B(G137), .Z(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(G39));
  NAND2_X1  g648(.A1(new_n817), .A2(new_n823), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n743), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT46), .B1(new_n817), .B2(new_n819), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n315), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n319), .B1(new_n324), .B2(new_n814), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n818), .B1(new_n842), .B2(new_n816), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n824), .B1(new_n843), .B2(KEYINPUT46), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n315), .A3(new_n839), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n740), .A2(new_n494), .A3(new_n411), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n803), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n841), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(G140), .ZN(G42));
  NAND3_X1  g663(.A1(new_n493), .A2(new_n318), .A3(new_n496), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT111), .Z(new_n851));
  NOR2_X1   g665(.A1(new_n752), .A2(new_n299), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n668), .B(new_n804), .C1(new_n853), .C2(KEYINPUT49), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT112), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n853), .A2(KEYINPUT49), .ZN(new_n857));
  NOR4_X1   g671(.A1(new_n856), .A2(new_n723), .A3(new_n708), .A4(new_n857), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT113), .Z(new_n859));
  NAND3_X1  g673(.A1(new_n783), .A2(new_n647), .A3(new_n754), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n826), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n790), .B1(KEYINPUT119), .B2(KEYINPUT48), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n863), .B(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n708), .A2(new_n496), .A3(new_n745), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n826), .A2(new_n700), .A3(new_n761), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT50), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n866), .A2(KEYINPUT50), .A3(new_n867), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n870), .A2(new_n871), .B1(new_n771), .B2(new_n861), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n722), .A2(new_n493), .ZN(new_n873));
  OR3_X1    g687(.A1(new_n860), .A2(KEYINPUT117), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT117), .B1(new_n860), .B2(new_n873), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n608), .A3(new_n668), .A4(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n841), .A2(new_n845), .B1(new_n316), .B2(new_n852), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n867), .A2(new_n783), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT51), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n865), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n874), .A2(new_n674), .A3(new_n875), .ZN(new_n884));
  INV_X1    g698(.A(G952), .ZN(new_n885));
  INV_X1    g699(.A(new_n755), .ZN(new_n886));
  AOI211_X1 g700(.A(new_n885), .B(G953), .C1(new_n867), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT118), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n880), .A2(KEYINPUT116), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n877), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(KEYINPUT116), .B2(new_n880), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n883), .B(new_n889), .C1(new_n892), .C2(KEYINPUT51), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n645), .B1(new_n608), .B2(new_n738), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n676), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n327), .A3(new_n659), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n757), .A3(new_n765), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n746), .B(new_n677), .C1(new_n685), .C2(new_n674), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n652), .A2(new_n697), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n783), .A2(new_n787), .A3(new_n775), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n801), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n683), .A2(new_n644), .A3(new_n702), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n317), .B2(new_n326), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n704), .A3(new_n783), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT114), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT114), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n905), .A2(new_n908), .A3(new_n704), .A4(new_n783), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n903), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n799), .A2(new_n901), .A3(new_n910), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n722), .A2(new_n763), .A3(new_n724), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n311), .A2(new_n753), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n726), .A2(new_n693), .A3(new_n702), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n913), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NOR4_X1   g731(.A1(new_n311), .A2(new_n915), .A3(KEYINPUT115), .A4(new_n753), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n919), .A2(new_n705), .A3(new_n741), .A4(new_n777), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT52), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n894), .B1(new_n911), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n910), .A2(new_n901), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT52), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n920), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n705), .A2(new_n777), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT52), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n894), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n923), .A2(new_n925), .A3(new_n799), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT54), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n894), .B1(new_n926), .B2(KEYINPUT52), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n923), .A2(new_n925), .A3(new_n799), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n922), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n931), .B1(KEYINPUT54), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n893), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(G952), .A2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n859), .B1(new_n936), .B2(new_n937), .ZN(G75));
  NAND3_X1  g752(.A1(new_n934), .A2(G210), .A3(G902), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n516), .A2(new_n528), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n502), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT55), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n939), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n939), .B2(new_n940), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n360), .A2(G952), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G51));
  XNOR2_X1  g761(.A(new_n818), .B(KEYINPUT57), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n934), .A2(KEYINPUT54), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT54), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n922), .B2(new_n933), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n948), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n288), .A2(new_n298), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n934), .A2(G902), .A3(new_n816), .A4(new_n842), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n946), .B1(new_n954), .B2(new_n955), .ZN(G54));
  INV_X1    g770(.A(new_n946), .ZN(new_n957));
  NAND2_X1  g771(.A1(KEYINPUT58), .A2(G475), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n300), .B(new_n958), .C1(new_n922), .C2(new_n933), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n669), .A2(new_n670), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n962));
  INV_X1    g776(.A(new_n960), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT120), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n946), .B1(new_n962), .B2(new_n963), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT120), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n959), .A2(new_n960), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n965), .A2(new_n969), .ZN(G60));
  NOR2_X1   g784(.A1(new_n663), .A2(new_n664), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n666), .B(KEYINPUT59), .Z(new_n972));
  OAI211_X1 g786(.A(new_n971), .B(new_n972), .C1(new_n949), .C2(new_n951), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n957), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n971), .B1(new_n935), .B2(new_n972), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(G63));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT60), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n922), .B2(new_n933), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n979), .A2(new_n489), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n946), .B1(new_n979), .B2(new_n692), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT121), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n979), .B2(new_n692), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n984), .A2(KEYINPUT61), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n980), .B(new_n981), .C1(new_n984), .C2(KEYINPUT61), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(G66));
  INV_X1    g802(.A(new_n649), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n360), .B1(new_n989), .B2(G224), .ZN(new_n990));
  INV_X1    g804(.A(new_n901), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n990), .B1(new_n991), .B2(new_n360), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n941), .B1(G898), .B2(new_n360), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT122), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n992), .B(new_n994), .ZN(G69));
  XOR2_X1   g809(.A(new_n381), .B(new_n583), .Z(new_n996));
  INV_X1    g810(.A(KEYINPUT124), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n705), .A2(new_n741), .A3(new_n777), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n763), .A2(new_n790), .A3(new_n724), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n844), .A2(new_n315), .A3(new_n999), .A4(new_n730), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n801), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n998), .A2(new_n1001), .A3(new_n832), .A4(new_n848), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n997), .B1(new_n1003), .B2(new_n799), .ZN(new_n1004));
  INV_X1    g818(.A(new_n793), .ZN(new_n1005));
  AND4_X1   g819(.A1(new_n495), .A2(new_n783), .A3(new_n740), .A4(new_n787), .ZN(new_n1006));
  AOI21_X1  g820(.A(KEYINPUT42), .B1(new_n1006), .B2(KEYINPUT107), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1005), .B1(new_n1007), .B2(new_n796), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n1008), .A2(new_n1002), .A3(KEYINPUT124), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n360), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n360), .A2(G900), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(KEYINPUT125), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(KEYINPUT124), .B1(new_n1008), .B2(new_n1002), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n1001), .A2(new_n832), .A3(new_n848), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1015), .A2(new_n799), .A3(new_n997), .A4(new_n998), .ZN(new_n1016));
  AOI21_X1  g830(.A(G953), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT125), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n1017), .A2(new_n1018), .A3(new_n1011), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n996), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n998), .ZN(new_n1021));
  OAI21_X1  g835(.A(KEYINPUT62), .B1(new_n736), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT62), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n998), .B(new_n1023), .C1(new_n735), .C2(new_n734), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n803), .B1(KEYINPUT123), .B2(new_n895), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n895), .A2(KEYINPUT123), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n1025), .A2(new_n1026), .A3(new_n495), .A4(new_n732), .ZN(new_n1027));
  AND3_X1   g841(.A1(new_n832), .A2(new_n848), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1022), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(new_n996), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1029), .A2(new_n360), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1011), .B1(new_n261), .B2(G953), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(KEYINPUT126), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1020), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1033), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1010), .A2(KEYINPUT125), .A3(new_n1012), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1018), .B1(new_n1017), .B2(new_n1011), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1030), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1031), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1035), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1034), .A2(new_n1040), .ZN(G72));
  NOR3_X1   g855(.A1(new_n1004), .A2(new_n1009), .A3(new_n991), .ZN(new_n1042));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT63), .Z(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n385), .B(new_n382), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1046));
  AND2_X1   g860(.A1(new_n402), .A2(new_n406), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1045), .B1(new_n1047), .B2(new_n709), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n946), .B1(new_n930), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1044), .B1(new_n1029), .B2(new_n991), .ZN(new_n1050));
  OAI211_X1 g864(.A(new_n1050), .B(new_n371), .C1(new_n378), .C2(new_n405), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1046), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1052), .A2(KEYINPUT127), .ZN(new_n1053));
  INV_X1    g867(.A(KEYINPUT127), .ZN(new_n1054));
  NAND4_X1  g868(.A1(new_n1046), .A2(new_n1049), .A3(new_n1054), .A4(new_n1051), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1053), .A2(new_n1055), .ZN(G57));
endmodule


