//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1251, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  AND2_X1   g0026(.A1(KEYINPUT65), .A2(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(KEYINPUT65), .A2(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n202), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n212), .B(new_n226), .C1(new_n231), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n214), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n245), .B(new_n251), .ZN(G351));
  AOI21_X1  g0052(.A(new_n206), .B1(new_n201), .B2(new_n246), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n229), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n255), .A2(new_n257), .B1(G150), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n253), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(new_n260), .B2(new_n259), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n230), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n264), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n246), .B1(new_n205), .B2(G20), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n268), .A2(new_n269), .B1(new_n246), .B2(new_n267), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT9), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n277), .A3(G274), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G226), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XOR2_X1   g0082(.A(new_n282), .B(KEYINPUT66), .Z(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(G222), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n286), .B1(new_n220), .B2(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  AND2_X1   g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(new_n230), .ZN(new_n292));
  INV_X1    g0092(.A(new_n230), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(KEYINPUT67), .A3(new_n276), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n283), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(G200), .B2(new_n298), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n272), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n283), .A2(new_n306), .A3(new_n297), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n271), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n254), .A2(new_n220), .B1(new_n206), .B2(G68), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n310), .A2(KEYINPUT73), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n258), .A2(G50), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n310), .B2(KEYINPUT73), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n264), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT11), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT70), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n266), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n205), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n214), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT12), .ZN(new_n322));
  INV_X1    g0122(.A(G13), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(G1), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT12), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(G20), .A4(new_n214), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n264), .B1(new_n318), .B2(new_n319), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n214), .B1(new_n205), .B2(G20), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n322), .A2(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n314), .B2(new_n315), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n316), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n278), .B1(new_n280), .B2(new_n215), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT71), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n333), .B(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n284), .A2(G232), .A3(G1698), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n284), .A2(G226), .A3(new_n285), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n296), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT13), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT13), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n335), .A2(new_n343), .A3(new_n340), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n346), .A3(G169), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n306), .B2(new_n345), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n346), .B1(new_n345), .B2(G169), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n332), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n331), .B1(new_n299), .B2(new_n345), .ZN(new_n351));
  INV_X1    g0151(.A(G200), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n342), .B2(new_n344), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT72), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n353), .A2(KEYINPUT72), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OR2_X1    g0157(.A1(KEYINPUT65), .A2(G20), .ZN(new_n358));
  NAND2_X1  g0158(.A1(KEYINPUT65), .A2(G20), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n257), .A2(new_n258), .B1(new_n360), .B2(G77), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT15), .B(G87), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(new_n362), .B2(new_n254), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(new_n264), .B1(new_n220), .B2(new_n320), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n205), .A2(G20), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n327), .A2(G77), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n287), .A2(new_n215), .B1(new_n222), .B2(new_n284), .ZN(new_n368));
  INV_X1    g0168(.A(G33), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT3), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT3), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G33), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G232), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n373), .A2(new_n374), .A3(G1698), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n296), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n278), .B1(new_n280), .B2(new_n221), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n377), .A2(KEYINPUT69), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(KEYINPUT69), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n367), .B1(G200), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n299), .B2(new_n380), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n304), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n383), .B(new_n367), .C1(G179), .C2(new_n380), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n309), .A2(new_n350), .A3(new_n357), .A4(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n278), .B1(new_n280), .B2(new_n374), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT74), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n371), .ZN(new_n389));
  NAND2_X1  g0189(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(G33), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n370), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n281), .A2(G1698), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(G223), .B2(G1698), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n392), .A2(new_n394), .B1(new_n369), .B2(new_n216), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n387), .B1(new_n395), .B2(new_n296), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G179), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n304), .B2(new_n396), .ZN(new_n398));
  INV_X1    g0198(.A(G58), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n399), .A2(new_n214), .ZN(new_n400));
  OAI21_X1  g0200(.A(G20), .B1(new_n400), .B2(new_n201), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n258), .A2(G159), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n370), .ZN(new_n404));
  AND2_X1   g0204(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n405));
  NOR2_X1   g0205(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n404), .B1(new_n407), .B2(G33), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT7), .B1(new_n408), .B2(G20), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n360), .A2(KEYINPUT7), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n214), .B1(new_n410), .B2(new_n392), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n403), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT16), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n264), .ZN(new_n414));
  INV_X1    g0214(.A(new_n403), .ZN(new_n415));
  AOI21_X1  g0215(.A(G20), .B1(new_n370), .B2(new_n372), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT75), .B1(new_n416), .B2(KEYINPUT7), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT75), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT7), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n418), .B(new_n419), .C1(new_n284), .C2(G20), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n372), .B1(new_n407), .B2(G33), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n360), .A2(new_n419), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n417), .A2(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n415), .B1(new_n423), .B2(new_n214), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT16), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT76), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n424), .A2(KEYINPUT76), .A3(new_n425), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n414), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n268), .A2(new_n257), .A3(new_n365), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n266), .B2(new_n257), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT77), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n398), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  XOR2_X1   g0235(.A(new_n435), .B(KEYINPUT18), .Z(new_n436));
  INV_X1    g0236(.A(new_n429), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT76), .B1(new_n424), .B2(new_n425), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n264), .B(new_n413), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n396), .A2(new_n352), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(G190), .B2(new_n396), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n441), .A3(new_n433), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n442), .B(KEYINPUT17), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n436), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n386), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n417), .A2(new_n420), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n421), .A2(new_n422), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n222), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n258), .A2(G77), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n450), .B(KEYINPUT78), .ZN(new_n451));
  XNOR2_X1  g0251(.A(G97), .B(G107), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(KEYINPUT79), .B2(KEYINPUT6), .ZN(new_n453));
  NOR2_X1   g0253(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n454));
  INV_X1    g0254(.A(G97), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(KEYINPUT6), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n453), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n451), .B1(new_n457), .B2(new_n229), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n264), .B1(new_n449), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n266), .A2(G97), .ZN(new_n460));
  AOI211_X1 g0260(.A(new_n264), .B(new_n267), .C1(new_n205), .C2(G33), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(G97), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n391), .A2(G244), .A3(new_n285), .A4(new_n370), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT4), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(KEYINPUT4), .A2(G244), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n370), .A2(new_n372), .A3(new_n466), .A4(new_n285), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n370), .A2(new_n372), .A3(G250), .A4(G1698), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n295), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n205), .A2(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G274), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n293), .B2(new_n276), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g0279(.A(KEYINPUT5), .B(G41), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n274), .A2(G1), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n480), .A2(new_n481), .B1(new_n293), .B2(new_n276), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G257), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(G200), .B1(new_n471), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n277), .A2(G274), .ZN(new_n487));
  INV_X1    g0287(.A(new_n475), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n481), .B1(new_n488), .B2(new_n473), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(G257), .B2(new_n482), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n464), .B2(new_n463), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n491), .B(G190), .C1(new_n493), .C2(new_n295), .ZN(new_n494));
  AND4_X1   g0294(.A1(new_n459), .A2(new_n462), .A3(new_n486), .A4(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(G169), .B1(new_n471), .B2(new_n485), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n491), .B(G179), .C1(new_n493), .C2(new_n295), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n459), .A2(new_n462), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n391), .A2(new_n229), .A3(G68), .A4(new_n370), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n216), .A2(new_n455), .A3(new_n222), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT19), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n338), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n500), .B1(new_n360), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n358), .A2(G33), .A3(G97), .A4(new_n359), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n501), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n499), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n264), .ZN(new_n507));
  INV_X1    g0307(.A(new_n362), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n461), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n320), .A2(new_n362), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G238), .A2(G1698), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n221), .B2(G1698), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(new_n391), .A3(new_n370), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G116), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n295), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n481), .A2(new_n217), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n277), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n472), .B2(new_n487), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n304), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n478), .A2(new_n481), .B1(new_n517), .B2(new_n277), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n514), .A2(new_n515), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n306), .B(new_n521), .C1(new_n522), .C2(new_n295), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n511), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(G190), .B(new_n521), .C1(new_n522), .C2(new_n295), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n506), .A2(new_n264), .B1(new_n320), .B2(new_n362), .ZN(new_n526));
  OAI21_X1  g0326(.A(G200), .B1(new_n516), .B2(new_n519), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n461), .A2(G87), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n525), .A2(new_n526), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n495), .A2(new_n498), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n531), .B(KEYINPUT80), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n391), .A2(new_n229), .A3(G87), .A4(new_n370), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT22), .ZN(new_n534));
  XNOR2_X1  g0334(.A(KEYINPUT83), .B(KEYINPUT22), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n229), .A2(new_n284), .A3(new_n535), .A4(G87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT84), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT23), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n360), .A2(new_n542), .A3(new_n222), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n515), .A2(G20), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(KEYINPUT85), .B2(KEYINPUT24), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n539), .A2(new_n540), .ZN(new_n546));
  AND4_X1   g0346(.A1(new_n541), .A2(new_n543), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n537), .A2(new_n538), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n538), .B1(new_n537), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n264), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n267), .A2(new_n222), .ZN(new_n551));
  NOR2_X1   g0351(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n552));
  OR2_X1    g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g0353(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n551), .B2(new_n552), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n461), .A2(G107), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n484), .A2(new_n285), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n391), .A2(new_n370), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT87), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT87), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n391), .A2(new_n561), .A3(new_n370), .A4(new_n558), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G294), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n391), .A2(G250), .A3(new_n285), .A4(new_n370), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n560), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n296), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT88), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(KEYINPUT88), .A3(new_n296), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n483), .A2(new_n223), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n490), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n568), .A2(new_n299), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n566), .A2(new_n571), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n572), .A2(KEYINPUT89), .B1(new_n352), .B2(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n569), .A2(new_n571), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT89), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n299), .A4(new_n568), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n557), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n569), .A2(new_n571), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT88), .B1(new_n565), .B2(new_n296), .ZN(new_n580));
  OAI21_X1  g0380(.A(G169), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n566), .A2(G179), .A3(new_n571), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n581), .A2(new_n582), .B1(new_n550), .B2(new_n556), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(G116), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n585), .B1(new_n205), .B2(G33), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n585), .A2(new_n320), .B1(new_n327), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n369), .A2(G97), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n358), .A2(new_n588), .A3(new_n359), .A4(new_n469), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n263), .A2(new_n230), .B1(G20), .B2(new_n585), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT20), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(KEYINPUT20), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n304), .B1(new_n587), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n482), .A2(G270), .B1(new_n476), .B2(new_n478), .ZN(new_n597));
  INV_X1    g0397(.A(G303), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n284), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(G257), .A2(G1698), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n223), .B2(G1698), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n599), .B1(new_n408), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n597), .B(KEYINPUT81), .C1(new_n602), .C2(new_n295), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT81), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n601), .A2(new_n391), .A3(new_n370), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n373), .A2(G303), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n295), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n489), .A2(G270), .A3(new_n277), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n479), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n604), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n596), .A2(KEYINPUT21), .A3(new_n603), .A4(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n607), .A2(new_n609), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n320), .A2(new_n585), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n327), .A2(new_n586), .ZN(new_n614));
  INV_X1    g0414(.A(new_n594), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT20), .B1(new_n589), .B2(new_n590), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n612), .A2(new_n617), .A3(G179), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n603), .A2(new_n610), .A3(G169), .A4(new_n617), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT21), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT82), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(KEYINPUT82), .A3(new_n621), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n603), .A2(new_n610), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G200), .ZN(new_n628));
  INV_X1    g0428(.A(new_n617), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n628), .B(new_n629), .C1(new_n299), .C2(new_n627), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n532), .A2(new_n584), .A3(new_n626), .A4(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n446), .A2(new_n631), .ZN(G372));
  INV_X1    g0432(.A(new_n308), .ZN(new_n633));
  XOR2_X1   g0433(.A(new_n384), .B(KEYINPUT92), .Z(new_n634));
  NAND2_X1  g0434(.A1(new_n357), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n350), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT93), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(KEYINPUT93), .A3(new_n350), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n443), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n436), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n633), .B1(new_n641), .B2(new_n303), .ZN(new_n642));
  INV_X1    g0442(.A(new_n524), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n524), .A2(new_n529), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n498), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n643), .B1(new_n645), .B2(KEYINPUT26), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n496), .A2(new_n497), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT91), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n647), .A2(new_n648), .B1(new_n459), .B2(new_n462), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n496), .A2(KEYINPUT91), .A3(new_n497), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n649), .A2(new_n644), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT90), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n611), .A2(new_n618), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n620), .A2(KEYINPUT82), .A3(new_n621), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT82), .B1(new_n620), .B2(new_n621), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n531), .B1(new_n658), .B2(new_n583), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n654), .B1(new_n659), .B2(new_n578), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n581), .A2(new_n582), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n557), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n626), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n572), .A2(KEYINPUT89), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n573), .A2(new_n352), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n577), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n557), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n663), .A2(new_n668), .A3(KEYINPUT90), .A4(new_n531), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n653), .B1(new_n660), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n642), .B1(new_n446), .B2(new_n670), .ZN(G369));
  NAND2_X1  g0471(.A1(new_n229), .A2(new_n324), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n626), .B(new_n630), .C1(new_n629), .C2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n629), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n658), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n557), .A2(new_n678), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n584), .A2(new_n685), .B1(new_n583), .B2(new_n678), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n583), .A2(new_n679), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n626), .A2(new_n678), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n584), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT94), .ZN(G399));
  INV_X1    g0494(.A(new_n209), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n205), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n500), .A2(G116), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n697), .A2(new_n698), .B1(new_n233), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  NOR2_X1   g0500(.A1(new_n631), .A2(new_n678), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT96), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n516), .A2(new_n570), .A3(new_n519), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n704), .A2(new_n566), .A3(new_n612), .ZN(new_n705));
  INV_X1    g0505(.A(new_n497), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n703), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n705), .A2(KEYINPUT96), .A3(KEYINPUT30), .A4(new_n706), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n708), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n306), .B1(new_n516), .B2(new_n519), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n471), .A2(new_n485), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n573), .A3(new_n627), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n711), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n678), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g0520(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n702), .B(new_n720), .C1(new_n718), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n459), .A2(new_n462), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n647), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n486), .A2(new_n494), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n644), .B(new_n725), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n626), .B2(new_n662), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n668), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n524), .B1(new_n645), .B2(KEYINPUT26), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n649), .A2(new_n644), .A3(new_n651), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n730), .B1(new_n731), .B2(KEYINPUT26), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n678), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n670), .A2(new_n678), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(new_n734), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n723), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT97), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n700), .B1(new_n739), .B2(G1), .ZN(G364));
  XNOR2_X1  g0540(.A(new_n684), .B(KEYINPUT98), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n360), .A2(new_n323), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G45), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n697), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n741), .B(new_n744), .C1(G330), .C2(new_n683), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n352), .A2(G179), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(G20), .A3(G190), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n229), .B1(G190), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G294), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n373), .B1(new_n598), .B2(new_n747), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n229), .A2(new_n306), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G200), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n751), .B1(G322), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(new_n299), .A3(new_n352), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n229), .A2(G190), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n748), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n757), .A2(G311), .B1(new_n760), .B2(G329), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n306), .A2(new_n352), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT33), .B(G317), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n758), .A2(new_n746), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n764), .A2(new_n765), .B1(new_n767), .B2(G283), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n753), .A2(new_n352), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G326), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n755), .A2(new_n761), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n756), .A2(KEYINPUT101), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n756), .A2(KEYINPUT101), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n754), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n774), .A2(new_n220), .B1(new_n399), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(KEYINPUT102), .ZN(new_n777));
  INV_X1    g0577(.A(G159), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n759), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n763), .A2(new_n214), .B1(new_n749), .B2(new_n455), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n284), .B1(new_n216), .B2(new_n747), .C1(new_n766), .C2(new_n222), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n781), .B(new_n782), .C1(G50), .C2(new_n769), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n777), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n776), .A2(KEYINPUT102), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n771), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n230), .B1(G20), .B2(new_n304), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n695), .A2(new_n373), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT99), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n790), .A2(G355), .B1(new_n585), .B2(new_n695), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n251), .A2(new_n274), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n695), .A2(new_n408), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(G45), .B2(new_n232), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n791), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n787), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT100), .Z(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n744), .B1(new_n795), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n798), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n788), .B(new_n802), .C1(new_n683), .C2(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n745), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  INV_X1    g0606(.A(new_n787), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n769), .A2(G137), .B1(new_n764), .B2(G150), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT103), .B(G143), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n808), .B1(new_n775), .B2(new_n809), .C1(new_n774), .C2(new_n778), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT34), .Z(new_n811));
  OAI221_X1 g0611(.A(new_n408), .B1(new_n246), .B2(new_n747), .C1(new_n749), .C2(new_n399), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n214), .A2(new_n766), .B1(new_n759), .B2(new_n813), .ZN(new_n814));
  OR3_X1    g0614(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n774), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G116), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n769), .A2(G303), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n373), .B1(new_n222), .B2(new_n747), .C1(new_n749), .C2(new_n455), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G294), .B2(new_n754), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n216), .A2(new_n766), .B1(new_n763), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G311), .B2(new_n760), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n817), .A2(new_n818), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n807), .B1(new_n815), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n787), .A2(new_n796), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(new_n220), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n634), .A2(new_n367), .A3(new_n678), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n678), .A2(new_n367), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n385), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n827), .B1(new_n797), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n744), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n722), .A2(G330), .ZN(new_n835));
  INV_X1    g0635(.A(new_n653), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT90), .B1(new_n728), .B2(new_n668), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n659), .A2(new_n654), .A3(new_n578), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT104), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n385), .A2(new_n679), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT104), .B1(new_n670), .B2(new_n841), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n736), .B2(new_n831), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n835), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n744), .B1(new_n835), .B2(new_n846), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n834), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n849), .A2(KEYINPUT105), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(KEYINPUT105), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G384));
  INV_X1    g0653(.A(KEYINPUT35), .ZN(new_n854));
  OAI211_X1 g0654(.A(G116), .B(new_n231), .C1(new_n457), .C2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n854), .B2(new_n457), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT36), .ZN(new_n857));
  OR3_X1    g0657(.A1(new_n232), .A2(new_n220), .A3(new_n400), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n205), .B(G13), .C1(new_n858), .C2(new_n247), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n348), .A2(new_n349), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n332), .B(new_n678), .C1(new_n861), .C2(new_n356), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n332), .A2(new_n678), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n357), .A2(new_n350), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT106), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n384), .A2(new_n678), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n866), .B1(new_n845), .B2(new_n868), .ZN(new_n869));
  AOI211_X1 g0669(.A(KEYINPUT106), .B(new_n867), .C1(new_n843), .C2(new_n844), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT107), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n840), .B1(new_n839), .B2(new_n842), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n670), .A2(KEYINPUT104), .A3(new_n841), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n868), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT106), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n845), .A2(new_n866), .A3(new_n868), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(KEYINPUT107), .A3(new_n865), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n442), .A2(new_n435), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n430), .A2(new_n434), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n884), .A2(KEYINPUT109), .A3(new_n676), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT109), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n439), .A2(new_n433), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n887), .B2(new_n675), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n882), .B(new_n883), .C1(new_n885), .C2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT110), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n442), .A2(new_n435), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT109), .B1(new_n884), .B2(new_n676), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n887), .A2(new_n886), .A3(new_n675), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(KEYINPUT110), .A3(new_n883), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n412), .A2(KEYINPUT16), .ZN(new_n897));
  INV_X1    g0697(.A(new_n264), .ZN(new_n898));
  OR3_X1    g0698(.A1(new_n897), .A2(KEYINPUT108), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT108), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n413), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n433), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n675), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n398), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n904), .A3(new_n442), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n891), .A2(new_n896), .B1(KEYINPUT37), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n903), .B1(new_n436), .B2(new_n443), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n881), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n889), .A2(new_n890), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT110), .B1(new_n895), .B2(new_n883), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n907), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n873), .A2(new_n880), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n436), .A2(new_n675), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n908), .A2(new_n914), .A3(KEYINPUT39), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n885), .A2(new_n888), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n444), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n895), .A2(new_n883), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n891), .B2(new_n896), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n881), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT39), .B1(new_n924), .B2(new_n914), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n918), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n861), .A2(new_n332), .A3(new_n679), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n917), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n916), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n642), .B1(new_n446), .B2(new_n737), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(G330), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n862), .A2(new_n864), .B1(new_n828), .B2(new_n830), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n718), .A2(new_n721), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n934), .B(new_n935), .C1(new_n938), .C2(new_n701), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n908), .B2(new_n914), .ZN(new_n940));
  INV_X1    g0740(.A(new_n934), .ZN(new_n941));
  INV_X1    g0741(.A(new_n938), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n941), .B1(new_n942), .B2(new_n702), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n910), .A2(new_n911), .B1(new_n883), .B2(new_n895), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT38), .B1(new_n944), .B2(new_n920), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n906), .A2(new_n881), .A3(new_n907), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n940), .B1(new_n947), .B2(KEYINPUT40), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n446), .B1(new_n702), .B2(new_n942), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n933), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n950), .B2(new_n949), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n932), .A2(new_n952), .B1(new_n205), .B2(new_n742), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT111), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n932), .A2(new_n952), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n953), .A2(KEYINPUT111), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n860), .B1(new_n956), .B2(new_n957), .ZN(G367));
  INV_X1    g0758(.A(G150), .ZN(new_n959));
  INV_X1    g0759(.A(new_n769), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n959), .A2(new_n775), .B1(new_n960), .B2(new_n809), .ZN(new_n961));
  INV_X1    g0761(.A(G137), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n759), .A2(new_n962), .B1(new_n399), .B2(new_n747), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n763), .A2(new_n778), .B1(new_n749), .B2(new_n214), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT113), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n373), .B1(new_n767), .B2(G77), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n816), .A2(G50), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n965), .B(new_n968), .C1(new_n966), .C2(new_n967), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n775), .A2(new_n598), .ZN(new_n970));
  INV_X1    g0770(.A(new_n747), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(G116), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT46), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n222), .B2(new_n749), .C1(new_n750), .C2(new_n763), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n970), .B(new_n974), .C1(G311), .C2(new_n769), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n821), .B2(new_n774), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n766), .A2(new_n455), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n408), .B(new_n977), .C1(G317), .C2(new_n760), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT112), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n969), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT47), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n787), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n526), .A2(new_n528), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n678), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n644), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n643), .A2(new_n983), .A3(new_n678), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n985), .A2(new_n798), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n800), .B1(new_n695), .B2(new_n508), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n793), .A2(new_n241), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n744), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n982), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n743), .A2(G1), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n584), .A2(new_n690), .ZN(new_n993));
  INV_X1    g0793(.A(new_n690), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(new_n686), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(G330), .A3(new_n683), .ZN(new_n996));
  INV_X1    g0796(.A(new_n741), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n997), .B2(new_n995), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n724), .A2(new_n678), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n725), .B(new_n1000), .C1(new_n724), .C2(new_n726), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n649), .A2(new_n651), .A3(new_n678), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n691), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT45), .Z(new_n1005));
  NOR2_X1   g0805(.A1(new_n691), .A2(new_n1003), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT44), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(new_n687), .Z(new_n1009));
  NAND3_X1  g0809(.A1(new_n739), .A2(new_n999), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n739), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n696), .B(KEYINPUT41), .Z(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n992), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n993), .A2(new_n1003), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1015), .A2(KEYINPUT42), .B1(new_n498), .B2(new_n679), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1003), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(KEYINPUT42), .B2(new_n688), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n692), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n985), .A2(new_n986), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1016), .A2(new_n1019), .B1(KEYINPUT43), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(KEYINPUT43), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1021), .B(new_n1022), .Z(new_n1023));
  NOR3_X1   g0823(.A1(new_n684), .A2(new_n686), .A3(new_n1017), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n991), .B1(new_n1014), .B2(new_n1026), .ZN(G387));
  INV_X1    g0827(.A(new_n739), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(new_n998), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n696), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n739), .A2(new_n999), .ZN(new_n1031));
  OR3_X1    g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n793), .B1(new_n238), .B2(new_n274), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n790), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n1034), .B2(new_n698), .ZN(new_n1035));
  OR3_X1    g0835(.A1(new_n256), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1036));
  OAI21_X1  g0836(.A(KEYINPUT50), .B1(new_n256), .B2(G50), .ZN(new_n1037));
  AOI21_X1  g0837(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1036), .A2(new_n698), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1035), .A2(new_n1039), .B1(new_n222), .B2(new_n695), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n408), .B1(new_n220), .B2(new_n747), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1041), .B(new_n977), .C1(G50), .C2(new_n754), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n778), .B2(new_n960), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n749), .A2(new_n362), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G150), .B2(new_n760), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n214), .B2(new_n756), .C1(new_n256), .C2(new_n763), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n754), .A2(G317), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n769), .A2(G322), .B1(new_n764), .B2(G311), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n774), .C2(new_n598), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n749), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1054), .A2(G283), .B1(new_n971), .B2(G294), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT49), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n766), .A2(new_n585), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n408), .B(new_n1058), .C1(G326), .C2(new_n760), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1047), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n833), .B1(new_n800), .B2(new_n1040), .C1(new_n1060), .C2(new_n807), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT114), .Z(new_n1062));
  NAND2_X1  g0862(.A1(new_n686), .A2(new_n798), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1062), .A2(new_n1063), .B1(new_n999), .B2(new_n992), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1032), .A2(new_n1064), .ZN(G393));
  NAND2_X1  g0865(.A1(new_n1009), .A2(new_n992), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n801), .B1(new_n455), .B2(new_n209), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n245), .A2(new_n695), .A3(new_n408), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n833), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n408), .B1(new_n214), .B2(new_n747), .C1(new_n766), .C2(new_n216), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1054), .A2(G77), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n759), .B2(new_n809), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(G50), .C2(new_n764), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n256), .B2(new_n774), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G150), .A2(new_n769), .B1(new_n754), .B2(G159), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT51), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G311), .A2(new_n754), .B1(new_n769), .B2(G317), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT52), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n757), .A2(G294), .B1(new_n764), .B2(G303), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n373), .B1(new_n747), .B2(new_n821), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n767), .B2(G107), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n760), .A2(G322), .B1(new_n1054), .B2(G116), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n1074), .A2(new_n1076), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1069), .B1(new_n1084), .B2(new_n787), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n1003), .B2(new_n803), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1066), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1029), .A2(new_n1009), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1010), .A2(new_n696), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(G390));
  NAND3_X1  g0890(.A1(new_n835), .A2(new_n831), .A3(new_n865), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n945), .A2(new_n946), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n865), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n867), .B1(new_n733), .B2(new_n831), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n927), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n928), .B1(new_n879), .B2(new_n865), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1091), .B(new_n1096), .C1(new_n1097), .C2(new_n926), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n992), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n933), .B1(new_n942), .B2(new_n702), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n934), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n871), .A2(new_n927), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT39), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n945), .B2(new_n946), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n908), .A2(new_n914), .A3(KEYINPUT39), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1102), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1101), .B1(new_n1108), .B2(KEYINPUT115), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT115), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n871), .A2(new_n927), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n1102), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1099), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n926), .A2(new_n797), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n826), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT54), .B(G143), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n816), .A2(new_n1117), .B1(G137), .B2(new_n764), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1118), .A2(KEYINPUT116), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n747), .B2(new_n959), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1120), .A2(new_n747), .A3(new_n959), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1122), .A2(new_n373), .ZN(new_n1123));
  INV_X1    g0923(.A(G128), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1121), .B(new_n1123), .C1(new_n960), .C2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n760), .A2(G125), .B1(new_n767), .B2(G50), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n778), .B2(new_n749), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(G132), .C2(new_n754), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1118), .A2(KEYINPUT116), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1119), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n816), .A2(G97), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n769), .A2(G283), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n373), .B1(new_n216), .B2(new_n747), .C1(new_n766), .C2(new_n214), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G116), .B2(new_n754), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1071), .B1(new_n750), .B2(new_n759), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G107), .B2(new_n764), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1130), .A2(new_n1137), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n833), .B1(new_n257), .B2(new_n1115), .C1(new_n1138), .C2(new_n807), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1114), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(KEYINPUT118), .B1(new_n1113), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1101), .ZN(new_n1142));
  OAI211_X1 g0942(.A(KEYINPUT115), .B(new_n1096), .C1(new_n1097), .C2(new_n926), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1112), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n992), .A3(new_n1098), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT118), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1140), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1141), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n445), .A2(new_n1100), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1150), .B(new_n642), .C1(new_n446), .C2(new_n737), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1100), .A2(new_n831), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1091), .B(new_n1094), .C1(new_n865), .C2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n722), .A2(G330), .A3(new_n831), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1154), .A2(new_n1093), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n879), .B1(new_n1155), .B2(new_n1142), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1151), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1144), .A2(new_n1157), .A3(new_n1098), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1144), .B2(new_n1098), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n1030), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT119), .B1(new_n1149), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1159), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1144), .A2(new_n1157), .A3(new_n1098), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n696), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT119), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1164), .A2(new_n1165), .A3(new_n1148), .A4(new_n1141), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1161), .A2(new_n1166), .ZN(G378));
  INV_X1    g0967(.A(new_n1151), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n303), .A2(new_n308), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT123), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1170), .B(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n271), .A2(new_n675), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT122), .Z(new_n1175));
  XOR2_X1   g0975(.A(new_n1173), .B(new_n1175), .Z(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n948), .B2(new_n933), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1173), .B(new_n1175), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n924), .A2(new_n914), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n935), .B1(new_n1179), .B2(new_n943), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1178), .B(G330), .C1(new_n1180), .C2(new_n940), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n930), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1177), .A2(new_n916), .A3(new_n1181), .A4(new_n929), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1183), .A2(KEYINPUT57), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1169), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1186), .B(new_n696), .C1(new_n1188), .C2(KEYINPUT57), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1183), .A2(new_n992), .A3(new_n1184), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n833), .B1(G50), .B2(new_n1115), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n369), .A2(new_n273), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT120), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n246), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n273), .B2(new_n392), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n455), .A2(new_n763), .B1(new_n759), .B2(new_n821), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n508), .B2(new_n757), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1054), .A2(G68), .B1(new_n971), .B2(G77), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n766), .A2(new_n399), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1199), .A2(G41), .A3(new_n408), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G107), .A2(new_n754), .B1(new_n769), .B2(G116), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT58), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1195), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1193), .B1(new_n760), .B2(G124), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n757), .A2(G137), .B1(new_n971), .B2(new_n1117), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n813), .B2(new_n763), .C1(new_n1124), .C2(new_n775), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n769), .A2(G125), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n959), .B2(new_n749), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1209), .A2(KEYINPUT121), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(KEYINPUT121), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1207), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT59), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1205), .B1(new_n778), .B2(new_n766), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1204), .B1(new_n1203), .B2(new_n1202), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1191), .B1(new_n1216), .B2(new_n787), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1176), .B2(new_n797), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1190), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1189), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n992), .B(KEYINPUT124), .Z(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n833), .B1(G68), .B2(new_n1115), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n585), .A2(new_n763), .B1(new_n759), .B2(new_n598), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1044), .B(new_n1226), .C1(G97), .C2(new_n971), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G283), .A2(new_n754), .B1(new_n769), .B2(G294), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(new_n222), .C2(new_n774), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n373), .B1(new_n766), .B2(new_n220), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT125), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n392), .B(new_n1199), .C1(G159), .C2(new_n971), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n813), .B2(new_n960), .C1(new_n962), .C2(new_n775), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n757), .A2(G150), .B1(G50), .B2(new_n1054), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n1124), .B2(new_n759), .C1(new_n763), .C2(new_n1116), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n1229), .A2(new_n1231), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1225), .B1(new_n1236), .B2(new_n787), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n865), .B2(new_n797), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1224), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1221), .A2(new_n1168), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1153), .A2(new_n1156), .A3(new_n1151), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n1013), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(new_n1243), .ZN(G381));
  OR4_X1    g1044(.A1(G396), .A2(G393), .A3(G384), .A4(G390), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1245), .A2(G387), .A3(G381), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1149), .A2(new_n1160), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1246), .A2(new_n1247), .A3(new_n1189), .A4(new_n1219), .ZN(G407));
  NAND2_X1  g1048(.A1(new_n677), .A2(G213), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G407), .B(G213), .C1(G375), .C2(new_n1251), .ZN(G409));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1161), .A2(new_n1166), .A3(new_n1189), .A4(new_n1219), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1188), .A2(new_n1013), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1218), .B1(new_n1187), .B2(new_n1222), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1247), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1250), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1153), .A2(new_n1156), .A3(KEYINPUT60), .A4(new_n1151), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n696), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1241), .A2(KEYINPUT60), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1260), .B1(new_n1261), .B2(new_n1242), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1263), .A2(KEYINPUT126), .A3(new_n852), .A4(new_n1240), .ZN(new_n1264));
  OR2_X1    g1064(.A1(new_n852), .A2(KEYINPUT126), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n852), .A2(KEYINPUT126), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1265), .B(new_n1266), .C1(new_n1262), .C2(new_n1239), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1250), .A2(G2897), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1268), .B(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1253), .B1(new_n1258), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT63), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1249), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1268), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1273), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(G387), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(G390), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G387), .B(new_n1087), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(G393), .B(G396), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT127), .B1(new_n1278), .B2(G390), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT127), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1279), .A2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G387), .B(G390), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G393), .B(new_n805), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1284), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1268), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1272), .A2(new_n1277), .A3(new_n1290), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1258), .A2(new_n1293), .A3(new_n1268), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1293), .B1(new_n1258), .B2(new_n1268), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1294), .A2(new_n1271), .A3(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1292), .B1(new_n1296), .B2(new_n1290), .ZN(G405));
  NAND2_X1  g1097(.A1(G375), .A2(new_n1247), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1254), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1290), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1284), .A2(new_n1289), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(new_n1254), .A3(new_n1298), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1303), .B(new_n1276), .ZN(G402));
endmodule


