//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT64), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  AND3_X1   g038(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT65), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT65), .B1(new_n461), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n462), .ZN(new_n470));
  NAND3_X1  g045(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(G101), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(new_n475), .ZN(G160));
  AND3_X1   g051(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n472), .A2(KEYINPUT67), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n483), .A2(new_n459), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n459), .A2(G138), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n470), .B2(new_n471), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT69), .B1(new_n479), .B2(new_n493), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n462), .A2(G2104), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT65), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n492), .A2(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n493), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n496), .A2(new_n497), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n509));
  NAND2_X1  g084(.A1(G126), .A2(G2105), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n472), .B2(new_n511), .ZN(new_n512));
  AOI211_X1 g087(.A(KEYINPUT68), .B(new_n510), .C1(new_n470), .C2(new_n471), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n459), .A2(G114), .ZN(new_n514));
  OAI21_X1  g089(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n508), .A2(new_n516), .ZN(G164));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT71), .B1(new_n518), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G651), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G50), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n525), .A2(new_n529), .ZN(new_n533));
  INV_X1    g108(.A(G88), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n528), .A2(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n531), .A2(G51), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n542));
  INV_X1    g117(.A(G89), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n541), .B(new_n542), .C1(new_n533), .C2(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  AOI22_X1  g120(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n527), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n531), .A2(G52), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n533), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n527), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n531), .A2(G43), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n533), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  AOI22_X1  g137(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(new_n527), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n525), .A2(new_n529), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n531), .A2(G53), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n566), .B(KEYINPUT9), .C1(new_n530), .C2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n565), .A2(G91), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n564), .A2(new_n571), .ZN(G299));
  OR2_X1    g147(.A1(new_n547), .A2(new_n550), .ZN(G301));
  NAND2_X1  g148(.A1(new_n531), .A2(G49), .ZN(new_n574));
  INV_X1    g149(.A(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n533), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n523), .A2(new_n524), .ZN(new_n577));
  INV_X1    g152(.A(G74), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n527), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n576), .A2(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n565), .A2(G86), .B1(G48), .B2(new_n531), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(KEYINPUT73), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n584), .A2(KEYINPUT73), .A3(G651), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n581), .B1(new_n586), .B2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n565), .A2(G85), .B1(G47), .B2(new_n531), .ZN(new_n589));
  AND2_X1   g164(.A1(G72), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n525), .B2(G60), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT74), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI211_X1 g168(.A(KEYINPUT74), .B(new_n590), .C1(new_n525), .C2(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n589), .B1(new_n593), .B2(new_n594), .ZN(G290));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(G301), .A2(new_n596), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n525), .A2(G92), .A3(new_n529), .ZN(new_n598));
  XOR2_X1   g173(.A(KEYINPUT75), .B(KEYINPUT10), .Z(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n531), .A2(G54), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n525), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n527), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n597), .B1(new_n606), .B2(new_n596), .ZN(G284));
  AOI21_X1  g182(.A(new_n597), .B1(new_n606), .B2(new_n596), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g193(.A1(new_n460), .A2(G2105), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n503), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n620), .B(new_n621), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n484), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n486), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n459), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n624), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XOR2_X1   g208(.A(G2443), .B(G2446), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT79), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT78), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n635), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT14), .ZN(new_n645));
  OAI21_X1  g220(.A(G14), .B1(new_n639), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n639), .ZN(G401));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT80), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT82), .Z(new_n650));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(KEYINPUT17), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n652), .B(new_n654), .C1(new_n650), .C2(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n650), .A2(new_n655), .A3(new_n653), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n649), .A2(new_n651), .A3(new_n654), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n656), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT83), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT20), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n665), .A2(new_n667), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n674), .A2(new_n670), .A3(new_n668), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n672), .B(new_n675), .C1(new_n670), .C2(new_n674), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G229));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G22), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G166), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1971), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n683), .A2(G6), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G305), .B2(G16), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT32), .B(G1981), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n689), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n683), .A2(G23), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n576), .A2(new_n579), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(new_n683), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT33), .B(G1976), .Z(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT88), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  NOR4_X1   g273(.A1(new_n686), .A2(new_n691), .A3(new_n692), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT89), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT34), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G25), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT84), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n484), .A2(G131), .ZN(new_n707));
  OR2_X1    g282(.A1(G95), .A2(G2105), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n708), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n486), .A2(G119), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT85), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT85), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n706), .B1(new_n714), .B2(new_n704), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT35), .B(G1991), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT86), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n715), .B(new_n717), .Z(new_n718));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n722));
  OR2_X1    g297(.A1(G16), .A2(G24), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G290), .B2(new_n683), .ZN(new_n724));
  INV_X1    g299(.A(G1986), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n725), .B2(new_n724), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n720), .A2(new_n721), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n702), .A2(new_n703), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n702), .A2(KEYINPUT36), .A3(new_n703), .A4(new_n728), .ZN(new_n732));
  NOR2_X1   g307(.A1(G171), .A2(new_n683), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G5), .B2(new_n683), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT97), .Z(new_n737));
  NOR2_X1   g312(.A1(G168), .A2(new_n683), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n683), .B2(G21), .ZN(new_n739));
  INV_X1    g314(.A(G1966), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT96), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n739), .A2(new_n740), .ZN(new_n743));
  INV_X1    g318(.A(G28), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(KEYINPUT30), .ZN(new_n745));
  AOI21_X1  g320(.A(G29), .B1(new_n744), .B2(KEYINPUT30), .ZN(new_n746));
  OR2_X1    g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  NAND2_X1  g322(.A1(KEYINPUT31), .A2(G11), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n745), .A2(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n629), .B2(new_n704), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n743), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n737), .A2(new_n742), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT98), .ZN(new_n753));
  NOR2_X1   g328(.A1(G4), .A2(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n606), .B2(G16), .ZN(new_n755));
  INV_X1    g330(.A(G1348), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n704), .A2(G26), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT93), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n486), .A2(G128), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n459), .A2(G116), .ZN(new_n762));
  OAI21_X1  g337(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n763));
  AND3_X1   g338(.A1(new_n484), .A2(KEYINPUT91), .A3(G140), .ZN(new_n764));
  AOI21_X1  g339(.A(KEYINPUT91), .B1(new_n484), .B2(G140), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n761), .B1(new_n762), .B2(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G29), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n767), .A2(KEYINPUT92), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(KEYINPUT92), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n760), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT94), .B(G2067), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n757), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G29), .A2(G33), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT25), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n503), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(new_n459), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n777), .B(new_n779), .C1(G139), .C2(new_n484), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n775), .B1(new_n780), .B2(G29), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n484), .A2(G141), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n486), .A2(G129), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT26), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n786), .A2(new_n787), .B1(G105), .B2(new_n619), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n782), .A2(new_n783), .A3(new_n788), .ZN(new_n789));
  MUX2_X1   g364(.A(G32), .B(new_n789), .S(G29), .Z(new_n790));
  XOR2_X1   g365(.A(KEYINPUT27), .B(G1996), .Z(new_n791));
  OAI22_X1  g366(.A1(new_n781), .A2(G2072), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n734), .A2(new_n735), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G19), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n557), .B2(G16), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n793), .B1(G1341), .B2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G2078), .ZN(new_n797));
  NOR2_X1   g372(.A1(G164), .A2(new_n704), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G27), .B2(new_n704), .ZN(new_n799));
  AOI211_X1 g374(.A(new_n792), .B(new_n796), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n683), .A2(G20), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT23), .Z(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G299), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1956), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n704), .A2(G35), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G162), .B2(new_n704), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT29), .Z(new_n809));
  INV_X1    g384(.A(G2090), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(KEYINPUT99), .ZN(new_n812));
  NAND2_X1  g387(.A1(G160), .A2(G29), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT24), .B(G34), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(new_n704), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT95), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(G2084), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G1341), .B2(new_n795), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n781), .A2(G2072), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n790), .A2(new_n791), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n821), .B(new_n822), .C1(new_n797), .C2(new_n799), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n810), .B2(new_n809), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n800), .A2(new_n812), .A3(new_n820), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n811), .A2(KEYINPUT99), .ZN(new_n826));
  NOR4_X1   g401(.A1(new_n753), .A2(new_n774), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n731), .A2(new_n732), .A3(new_n827), .ZN(G311));
  NAND3_X1  g403(.A1(new_n731), .A2(new_n732), .A3(new_n827), .ZN(G150));
  AOI22_X1  g404(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n527), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n531), .A2(G55), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n533), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G860), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n606), .A2(G559), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n557), .A2(new_n835), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n553), .A2(new_n556), .B1(new_n831), .B2(new_n834), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n841), .B(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n836), .B1(new_n845), .B2(KEYINPUT39), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n838), .B1(new_n846), .B2(new_n847), .ZN(G145));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n780), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n789), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n484), .A2(G142), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n486), .A2(G130), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n459), .A2(G118), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n852), .B(new_n853), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n622), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n850), .B(new_n789), .ZN(new_n859));
  INV_X1    g434(.A(new_n857), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n766), .B(G164), .Z(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(new_n714), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n714), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n858), .A2(new_n864), .A3(new_n865), .A4(new_n861), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n629), .B(G160), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n490), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  INV_X1    g448(.A(new_n871), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n867), .A2(new_n868), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT102), .ZN(new_n877));
  AOI21_X1  g452(.A(G37), .B1(new_n869), .B2(new_n871), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(new_n875), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n877), .A2(KEYINPUT40), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT40), .B1(new_n877), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(G395));
  NAND2_X1  g458(.A1(new_n604), .A2(new_n610), .ZN(new_n884));
  OAI21_X1  g459(.A(G299), .B1(new_n600), .B2(new_n603), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(KEYINPUT41), .A3(new_n885), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n615), .B(new_n844), .ZN(new_n891));
  MUX2_X1   g466(.A(new_n890), .B(new_n886), .S(new_n891), .Z(new_n892));
  XNOR2_X1  g467(.A(G290), .B(G288), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT103), .ZN(new_n894));
  XNOR2_X1  g469(.A(G305), .B(G303), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n893), .A2(KEYINPUT103), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n897), .A2(new_n895), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT42), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n892), .B(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(G868), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(G868), .B2(new_n835), .ZN(G295));
  OAI21_X1  g479(.A(new_n903), .B1(G868), .B2(new_n835), .ZN(G331));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n906));
  NAND2_X1  g481(.A1(G301), .A2(G286), .ZN(new_n907));
  NAND2_X1  g482(.A1(G171), .A2(G168), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(new_n844), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n907), .A2(new_n908), .B1(new_n842), .B2(new_n843), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n910), .A2(new_n886), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n890), .ZN(new_n913));
  INV_X1    g488(.A(new_n910), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n911), .A2(KEYINPUT104), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n909), .A2(KEYINPUT104), .A3(new_n844), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n912), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(G37), .B1(new_n918), .B2(new_n900), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n898), .B1(new_n895), .B2(new_n894), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n918), .B2(KEYINPUT105), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n910), .A2(new_n886), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n909), .A2(new_n844), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n911), .A2(KEYINPUT104), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n910), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n924), .B1(new_n928), .B2(new_n890), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n919), .B1(new_n921), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n910), .A2(new_n911), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT106), .B1(new_n890), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n922), .B1(new_n915), .B2(new_n916), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n890), .A2(KEYINPUT106), .A3(new_n935), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n920), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n919), .A3(KEYINPUT43), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n906), .B1(new_n934), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n919), .A3(new_n933), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT107), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n941), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n918), .A2(KEYINPUT105), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n929), .A2(new_n930), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n920), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT43), .B1(new_n950), .B2(new_n919), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT44), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n953));
  INV_X1    g528(.A(new_n944), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n933), .B1(new_n950), .B2(new_n919), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n952), .B(new_n953), .C1(new_n956), .C2(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n946), .A2(new_n957), .ZN(G397));
  OAI21_X1  g533(.A(new_n507), .B1(new_n464), .B2(new_n465), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n494), .A2(new_n495), .ZN(new_n960));
  INV_X1    g535(.A(G138), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(G2105), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n495), .B(new_n962), .C1(new_n477), .C2(new_n478), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT4), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n959), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n514), .A2(new_n515), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT68), .B1(new_n479), .B2(new_n510), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n472), .A2(new_n509), .A3(new_n511), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(KEYINPUT45), .ZN(new_n971));
  INV_X1    g546(.A(G40), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n468), .A2(new_n972), .A3(new_n475), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n766), .B(G2067), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n979), .A2(KEYINPUT109), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(KEYINPUT109), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n789), .B(G1996), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n980), .A2(new_n981), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n977), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n714), .B(new_n717), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(G290), .B(G1986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n977), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n973), .A2(new_n970), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(G8), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(G1976), .B2(new_n694), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(KEYINPUT111), .B(G1976), .Z(new_n994));
  OAI211_X1 g569(.A(new_n991), .B(new_n992), .C1(new_n694), .C2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n996));
  INV_X1    g571(.A(G1981), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n997), .B(new_n581), .C1(new_n586), .C2(new_n587), .ZN(new_n998));
  INV_X1    g573(.A(new_n581), .ZN(new_n999));
  OAI21_X1  g574(.A(G1981), .B1(new_n999), .B2(new_n585), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n996), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n990), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n993), .B(new_n995), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G303), .A2(G8), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT55), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n473), .A2(new_n474), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n459), .ZN(new_n1012));
  INV_X1    g587(.A(new_n467), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n503), .B2(G125), .ZN(new_n1014));
  OAI211_X1 g589(.A(G40), .B(new_n1012), .C1(new_n1014), .C2(new_n459), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(KEYINPUT45), .B2(new_n970), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n971), .A2(KEYINPUT110), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n970), .A2(new_n1018), .A3(KEYINPUT45), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1016), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1971), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n973), .B1(new_n970), .B2(new_n1023), .ZN(new_n1024));
  AOI211_X1 g599(.A(KEYINPUT50), .B(G1384), .C1(new_n965), .C2(new_n969), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n810), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1010), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1006), .B1(new_n1009), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n1031));
  INV_X1    g606(.A(G1384), .ZN(new_n1032));
  OAI211_X1 g607(.A(KEYINPUT45), .B(new_n1032), .C1(new_n508), .C2(new_n516), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n973), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1032), .B1(new_n508), .B2(new_n516), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n1018), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(KEYINPUT110), .A3(new_n1036), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1034), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1027), .B(new_n1031), .C1(new_n1040), .C2(G1971), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G8), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1031), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1030), .B(new_n1008), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1971), .B1(new_n1046), .B2(new_n1016), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1035), .A2(KEYINPUT50), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n970), .A2(new_n1023), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n973), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(G2090), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT114), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(G8), .A3(new_n1041), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1030), .B1(new_n1053), .B2(new_n1008), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1029), .B1(new_n1045), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT123), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT123), .B(new_n1029), .C1(new_n1045), .C2(new_n1054), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G286), .A2(G8), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1061), .A2(KEYINPUT119), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(KEYINPUT119), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1062), .A2(new_n1063), .A3(KEYINPUT51), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n740), .B1(new_n1034), .B2(new_n971), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1048), .A2(new_n1049), .A3(new_n818), .A4(new_n973), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1010), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g644(.A(KEYINPUT120), .B(new_n1010), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1060), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1024), .A2(G2084), .A3(new_n1025), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1966), .B1(new_n1016), .B2(new_n1037), .ZN(new_n1073));
  OAI21_X1  g648(.A(G8), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT120), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(KEYINPUT121), .A3(new_n1076), .A4(new_n1064), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT51), .B1(new_n1067), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1071), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1078), .B1(new_n1073), .B2(new_n1072), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1020), .B2(G2078), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1026), .A2(KEYINPUT117), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1050), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n735), .A3(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1016), .A2(KEYINPUT53), .A3(new_n797), .A4(new_n1037), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1085), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G171), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1083), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(KEYINPUT62), .ZN(new_n1097));
  AOI211_X1 g672(.A(KEYINPUT125), .B(new_n1081), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1094), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(G171), .B2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1085), .A2(G301), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1092), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1102), .B1(new_n1092), .B2(new_n1103), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1040), .A2(new_n1108), .ZN(new_n1109));
  XOR2_X1   g684(.A(G299), .B(KEYINPUT57), .Z(new_n1110));
  NAND2_X1  g685(.A1(new_n1050), .A2(new_n804), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1107), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1114), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(KEYINPUT61), .A3(new_n1112), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n989), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT58), .B(G1341), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1020), .A2(G1996), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n557), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1123), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(new_n557), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1086), .A2(new_n756), .A3(new_n1088), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n989), .A2(G2067), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1127), .A2(new_n606), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1124), .A2(new_n1126), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n606), .ZN(new_n1133));
  INV_X1    g708(.A(new_n606), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(new_n1129), .A3(new_n1127), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1128), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1118), .A2(new_n1131), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1113), .B1(new_n1133), .B2(new_n1116), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1096), .B(new_n1106), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1059), .B1(new_n1099), .B2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G288), .A2(G1976), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n990), .B1(new_n1142), .B2(new_n998), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1006), .B(KEYINPUT113), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1028), .A2(new_n1009), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1143), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1006), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1145), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1054), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(new_n1044), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1074), .A2(G286), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT63), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1008), .A2(KEYINPUT116), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1028), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(KEYINPUT63), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1028), .B2(new_n1154), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1144), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1147), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n988), .B1(new_n1140), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n766), .A2(G2067), .ZN(new_n1161));
  AOI211_X1 g736(.A(new_n717), .B(new_n710), .C1(new_n712), .C2(new_n713), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1161), .B1(new_n983), .B2(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n984), .A2(G1986), .A3(G290), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT48), .ZN(new_n1165));
  OAI22_X1  g740(.A1(new_n1163), .A2(new_n984), .B1(new_n986), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(G1996), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n977), .A2(KEYINPUT46), .A3(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT127), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT46), .B1(new_n977), .B2(new_n1167), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT126), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n978), .A2(new_n789), .ZN(new_n1172));
  AOI211_X1 g747(.A(new_n1169), .B(new_n1171), .C1(new_n977), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT47), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1166), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1160), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g753(.A(G319), .ZN(new_n1180));
  NOR4_X1   g754(.A1(G229), .A2(new_n1180), .A3(G401), .A4(G227), .ZN(new_n1181));
  INV_X1    g755(.A(new_n880), .ZN(new_n1182));
  AOI21_X1  g756(.A(new_n879), .B1(new_n878), .B2(new_n875), .ZN(new_n1183));
  OAI21_X1  g757(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g758(.A1(new_n1184), .A2(new_n956), .ZN(G308));
  OAI221_X1 g759(.A(new_n1181), .B1(new_n955), .B2(new_n954), .C1(new_n1182), .C2(new_n1183), .ZN(G225));
endmodule


