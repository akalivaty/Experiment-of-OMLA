//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206));
  NOR3_X1   g005(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n205), .B(new_n206), .C1(new_n207), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n211), .A2(new_n205), .A3(new_n206), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT79), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n208), .A2(KEYINPUT78), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT79), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G155gat), .B2(G162gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(G155gat), .A3(G162gat), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n215), .A2(new_n216), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n210), .B1(new_n212), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n202), .B1(new_n222), .B2(KEYINPUT3), .ZN(new_n223));
  AND2_X1   g022(.A1(G211gat), .A2(G218gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(G211gat), .A2(G218gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(G197gat), .A2(G204gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(G197gat), .A2(G204gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G211gat), .B(G218gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(G197gat), .B(G204gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n230), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n223), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT29), .B1(new_n231), .B2(new_n235), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n222), .B1(new_n238), .B2(KEYINPUT3), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G228gat), .A2(G233gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT81), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n241), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n237), .B(new_n239), .C1(new_n242), .C2(new_n241), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(G22gat), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT82), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n245), .ZN(new_n248));
  INV_X1    g047(.A(G22gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G78gat), .B(G106gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT31), .ZN(new_n252));
  INV_X1    g051(.A(G50gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  AND4_X1   g053(.A1(new_n246), .A2(new_n247), .A3(new_n250), .A4(new_n254), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n247), .A2(new_n254), .B1(new_n250), .B2(new_n246), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OR2_X1    g056(.A1(KEYINPUT70), .A2(G134gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(KEYINPUT70), .A2(G134gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(G127gat), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT71), .B(G127gat), .ZN(new_n261));
  INV_X1    g060(.A(G134gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n264));
  INV_X1    g063(.A(G113gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n265), .A2(G120gat), .ZN(new_n266));
  INV_X1    g065(.A(G120gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(G113gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n264), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n264), .B1(new_n262), .B2(G127gat), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n270), .B1(G127gat), .B2(new_n262), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(new_n265), .B2(G120gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n267), .A2(KEYINPUT72), .A3(G113gat), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n273), .B(new_n274), .C1(G113gat), .C2(new_n267), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n263), .A2(new_n269), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G169gat), .ZN(new_n277));
  INV_X1    g076(.A(G176gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT69), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT26), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT26), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n281), .A2(new_n277), .A3(new_n278), .A4(KEYINPUT69), .ZN(new_n282));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT27), .ZN(new_n288));
  INV_X1    g087(.A(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(KEYINPUT67), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G183gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n291), .B1(new_n295), .B2(KEYINPUT27), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n287), .B1(new_n296), .B2(G190gat), .ZN(new_n297));
  INV_X1    g096(.A(G190gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT68), .ZN(new_n299));
  NAND2_X1  g098(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n290), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n299), .B1(new_n290), .B2(new_n300), .ZN(new_n303));
  OAI211_X1 g102(.A(KEYINPUT28), .B(new_n298), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n286), .B1(new_n297), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT25), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT23), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(G169gat), .B2(G176gat), .ZN(new_n309));
  AND4_X1   g108(.A1(new_n306), .A2(new_n307), .A3(new_n309), .A4(new_n283), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT65), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n289), .A2(new_n298), .ZN(new_n314));
  NAND3_X1  g113(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n310), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n307), .A2(new_n309), .A3(new_n283), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT67), .B(G183gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n311), .B1(new_n319), .B2(new_n298), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(KEYINPUT66), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n322), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n318), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n317), .B1(new_n325), .B2(new_n306), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n276), .B1(new_n305), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT64), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n284), .A2(new_n285), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n290), .B1(new_n319), .B2(new_n288), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT28), .B1(new_n331), .B2(new_n298), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n298), .A2(KEYINPUT28), .ZN(new_n333));
  INV_X1    g132(.A(new_n303), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n333), .B1(new_n334), .B2(new_n301), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n330), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n292), .A2(new_n294), .A3(new_n298), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT24), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n285), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n337), .A2(new_n339), .A3(new_n321), .A4(new_n323), .ZN(new_n340));
  INV_X1    g139(.A(new_n318), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n339), .A2(new_n312), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n311), .A2(KEYINPUT65), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n315), .B(new_n314), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n342), .A2(KEYINPUT25), .B1(new_n345), .B2(new_n310), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n258), .A2(G127gat), .A3(new_n259), .ZN(new_n347));
  AND2_X1   g146(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n348), .A2(new_n349), .A3(new_n262), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n269), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n271), .A2(new_n275), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n346), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n327), .A2(new_n329), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT32), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT33), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G15gat), .B(G43gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n356), .B1(new_n362), .B2(KEYINPUT33), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n355), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n327), .A2(new_n354), .ZN(new_n366));
  INV_X1    g165(.A(new_n329), .ZN(new_n367));
  NOR2_X1   g166(.A1(KEYINPUT73), .A2(KEYINPUT34), .ZN(new_n368));
  AND2_X1   g167(.A1(KEYINPUT73), .A2(KEYINPUT34), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n305), .A2(new_n326), .A3(new_n276), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n353), .B1(new_n336), .B2(new_n346), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n367), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n368), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n363), .A2(new_n365), .A3(new_n370), .A4(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n355), .A2(new_n364), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n361), .B1(new_n355), .B2(new_n357), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n368), .B1(new_n366), .B2(new_n367), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n369), .A2(new_n368), .ZN(new_n380));
  AOI211_X1 g179(.A(new_n329), .B(new_n380), .C1(new_n327), .C2(new_n354), .ZN(new_n381));
  OAI22_X1  g180(.A1(new_n377), .A2(new_n378), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n257), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n222), .A2(KEYINPUT3), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n216), .A2(new_n220), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n211), .A2(new_n205), .A3(new_n206), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n218), .A4(new_n215), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n210), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n389), .A3(new_n353), .ZN(new_n390));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT4), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n353), .B2(new_n222), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n276), .A2(KEYINPUT4), .A3(new_n210), .A4(new_n387), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n390), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n391), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n353), .A2(new_n222), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n351), .A2(new_n352), .B1(new_n387), .B2(new_n210), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n399), .A3(KEYINPUT5), .ZN(new_n400));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT0), .ZN(new_n402));
  INV_X1    g201(.A(G57gat), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n403), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n404), .A2(new_n405), .A3(G85gat), .ZN(new_n406));
  AOI21_X1  g205(.A(G85gat), .B1(new_n404), .B2(new_n405), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n353), .B2(new_n222), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n396), .A2(KEYINPUT5), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n390), .A2(new_n410), .A3(new_n394), .A4(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n400), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT80), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n412), .ZN(new_n416));
  INV_X1    g215(.A(new_n408), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n400), .A2(new_n408), .A3(KEYINPUT80), .A4(new_n412), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n415), .A2(new_n418), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n408), .B1(new_n400), .B2(new_n412), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT6), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n426), .B1(new_n305), .B2(new_n326), .ZN(new_n427));
  INV_X1    g226(.A(new_n236), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT29), .B1(new_n336), .B2(new_n346), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n427), .B(new_n428), .C1(new_n429), .C2(new_n426), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n429), .A2(KEYINPUT76), .A3(new_n426), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT76), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n202), .B1(new_n305), .B2(new_n326), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(new_n425), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n427), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n431), .B1(new_n436), .B2(new_n236), .ZN(new_n437));
  XNOR2_X1  g236(.A(G64gat), .B(G92gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT77), .ZN(new_n439));
  XNOR2_X1  g238(.A(G8gat), .B(G36gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(KEYINPUT30), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n425), .B1(new_n336), .B2(new_n346), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT76), .B1(new_n429), .B2(new_n426), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n434), .A2(new_n433), .A3(new_n425), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n430), .B1(new_n446), .B2(new_n428), .ZN(new_n447));
  INV_X1    g246(.A(new_n441), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n430), .B(new_n441), .C1(new_n446), .C2(new_n428), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n424), .A2(new_n442), .A3(new_n449), .A4(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT35), .B1(new_n383), .B2(new_n453), .ZN(new_n454));
  AND4_X1   g253(.A1(new_n424), .A2(new_n442), .A3(new_n449), .A4(new_n452), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n376), .A2(new_n382), .A3(KEYINPUT74), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n379), .A2(new_n381), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT74), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n363), .A4(new_n365), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT35), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n455), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n454), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n376), .A2(new_n382), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT36), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n456), .A2(new_n465), .A3(new_n459), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT75), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n456), .A2(KEYINPUT75), .A3(new_n465), .A4(new_n459), .ZN(new_n470));
  INV_X1    g269(.A(new_n257), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n469), .A2(new_n470), .B1(new_n453), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n424), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT84), .B(KEYINPUT37), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n430), .B(new_n474), .C1(new_n446), .C2(new_n428), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n443), .B1(new_n425), .B2(new_n434), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n236), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n446), .B2(new_n236), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n475), .A2(new_n479), .A3(new_n480), .A4(new_n448), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n473), .A2(new_n450), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n448), .B(new_n475), .C1(new_n437), .C2(new_n476), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT38), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT85), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n486), .A3(KEYINPUT38), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n482), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n442), .A2(new_n449), .A3(new_n452), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n397), .A2(new_n398), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(new_n391), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n390), .A2(new_n410), .A3(new_n394), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n396), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n417), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n490), .A3(new_n396), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n495), .A2(KEYINPUT40), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT40), .B1(new_n495), .B2(new_n496), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n497), .A2(new_n498), .A3(new_n422), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n489), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n257), .ZN(new_n501));
  OAI22_X1  g300(.A1(new_n472), .A2(KEYINPUT83), .B1(new_n488), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n469), .A2(new_n470), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n453), .A2(new_n471), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n503), .A2(KEYINPUT83), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n463), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G229gat), .A2(G233gat), .ZN(new_n507));
  INV_X1    g306(.A(G29gat), .ZN(new_n508));
  INV_X1    g307(.A(G36gat), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT14), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT14), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n511), .A2(G29gat), .A3(G36gat), .ZN(new_n512));
  AOI211_X1 g311(.A(new_n510), .B(new_n512), .C1(G29gat), .C2(G36gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT15), .ZN(new_n514));
  XOR2_X1   g313(.A(G43gat), .B(G50gat), .Z(new_n515));
  NOR3_X1   g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(KEYINPUT86), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(new_n514), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT15), .B1(new_n515), .B2(KEYINPUT86), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT87), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT87), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n522), .B(new_n513), .C1(new_n518), .C2(new_n519), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n516), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(G1gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n527), .B(new_n528), .C1(G1gat), .C2(new_n525), .ZN(new_n529));
  NOR2_X1   g328(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n524), .A2(KEYINPUT17), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n531), .B1(new_n524), .B2(KEYINPUT17), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n507), .B(new_n532), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n524), .B(new_n531), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n507), .B(KEYINPUT89), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT13), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n536), .A2(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G113gat), .B(G141gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT11), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(new_n277), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(G197gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT12), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n538), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n547), .B1(new_n538), .B2(new_n542), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n506), .A2(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n524), .A2(KEYINPUT17), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT94), .B(G85gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G92gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G85gat), .A2(G92gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT7), .ZN(new_n559));
  INV_X1    g358(.A(G99gat), .ZN(new_n560));
  INV_X1    g359(.A(G106gat), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT8), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n557), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT95), .ZN(new_n564));
  XOR2_X1   g363(.A(G99gat), .B(G106gat), .Z(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n565), .ZN(new_n567));
  INV_X1    g366(.A(new_n565), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n557), .A2(new_n568), .A3(new_n559), .A4(new_n562), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(KEYINPUT95), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n553), .A2(new_n533), .A3(new_n566), .A4(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n524), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n566), .ZN(new_n573));
  AND2_X1   g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n572), .A2(new_n573), .B1(KEYINPUT41), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n576), .B(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n574), .A2(KEYINPUT41), .ZN(new_n580));
  XNOR2_X1  g379(.A(G190gat), .B(G218gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n579), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT9), .ZN(new_n585));
  INV_X1    g384(.A(G64gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(G57gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n403), .A2(G64gat), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT90), .ZN(new_n590));
  OR2_X1    g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OR3_X1    g392(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n590), .B1(new_n589), .B2(new_n593), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n587), .A2(KEYINPUT91), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n587), .A2(KEYINPUT91), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n597), .A3(new_n588), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n592), .B1(new_n591), .B2(new_n585), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n594), .A2(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT20), .ZN(new_n606));
  INV_X1    g405(.A(G211gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n531), .B1(new_n601), .B2(new_n602), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G183gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT93), .ZN(new_n612));
  XNOR2_X1  g411(.A(G127gat), .B(G155gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n610), .B(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n608), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n584), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT96), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n600), .B1(new_n570), .B2(new_n566), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n567), .A2(new_n569), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n624), .A2(new_n600), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n622), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n573), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n621), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n621), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n623), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G176gat), .ZN(new_n633));
  INV_X1    g432(.A(G204gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n619), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n552), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n473), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n489), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT16), .B(G8gat), .ZN(new_n646));
  OR3_X1    g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT97), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n644), .A2(new_n646), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n649), .A2(new_n645), .B1(G8gat), .B2(new_n644), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1325gat));
  INV_X1    g452(.A(new_n641), .ZN(new_n654));
  OAI21_X1  g453(.A(G15gat), .B1(new_n654), .B2(new_n503), .ZN(new_n655));
  INV_X1    g454(.A(new_n460), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(G15gat), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n655), .B1(new_n654), .B2(new_n657), .ZN(G1326gat));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n471), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT43), .B(G22gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  NOR3_X1   g460(.A1(new_n584), .A2(new_n618), .A3(new_n639), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n552), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(new_n508), .A3(new_n473), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT45), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n584), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n506), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT35), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n464), .A2(new_n255), .A3(new_n256), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n671), .B1(new_n455), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n461), .A2(new_n460), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n453), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n670), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n454), .A2(new_n462), .A3(KEYINPUT99), .ZN(new_n677));
  AND4_X1   g476(.A1(new_n421), .A2(new_n481), .A3(new_n423), .A4(new_n450), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n483), .A2(new_n486), .A3(KEYINPUT38), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n486), .B1(new_n483), .B2(KEYINPUT38), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n471), .B1(new_n489), .B2(new_n499), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n676), .A2(new_n677), .B1(new_n683), .B2(new_n472), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n667), .B1(new_n684), .B2(new_n584), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n618), .A2(new_n550), .A3(new_n639), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n669), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT100), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n669), .A2(new_n685), .A3(new_n689), .A4(new_n686), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G29gat), .B1(new_n691), .B2(new_n424), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n666), .A2(new_n692), .ZN(G1328gat));
  INV_X1    g492(.A(new_n489), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n663), .A2(G36gat), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT46), .ZN(new_n696));
  OAI21_X1  g495(.A(G36gat), .B1(new_n691), .B2(new_n694), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1329gat));
  NOR3_X1   g497(.A1(new_n663), .A2(G43gat), .A3(new_n656), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G43gat), .B1(new_n687), .B2(new_n503), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(KEYINPUT47), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n503), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n703), .A3(new_n690), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G43gat), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n699), .B1(new_n705), .B2(KEYINPUT101), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n704), .A2(new_n707), .A3(G43gat), .ZN(new_n708));
  AOI211_X1 g507(.A(KEYINPUT102), .B(KEYINPUT47), .C1(new_n706), .C2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT102), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n705), .A2(KEYINPUT101), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n708), .A3(new_n700), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n702), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT103), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n717), .B(new_n702), .C1(new_n709), .C2(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(G1330gat));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n471), .A2(new_n253), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT104), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n664), .A2(KEYINPUT105), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G50gat), .B1(new_n687), .B2(new_n257), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n720), .B(G50gat), .C1(new_n691), .C2(new_n257), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n664), .A2(new_n722), .B1(KEYINPUT105), .B2(KEYINPUT48), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(G1331gat));
  INV_X1    g527(.A(new_n684), .ZN(new_n729));
  INV_X1    g528(.A(new_n639), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n619), .A2(new_n551), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n424), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(new_n403), .ZN(G1332gat));
  NOR2_X1   g533(.A1(new_n732), .A2(new_n694), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  AND2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n735), .B2(new_n736), .ZN(G1333gat));
  INV_X1    g538(.A(new_n732), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n460), .B(KEYINPUT106), .Z(new_n741));
  AOI21_X1  g540(.A(G71gat), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n703), .A2(G71gat), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT107), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g545(.A1(new_n740), .A2(new_n471), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g547(.A1(new_n618), .A2(new_n551), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n729), .A2(new_n583), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n730), .B1(new_n750), .B2(KEYINPUT51), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(KEYINPUT51), .B2(new_n750), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(new_n473), .A3(new_n555), .ZN(new_n754));
  AND4_X1   g553(.A1(new_n639), .A2(new_n669), .A3(new_n685), .A4(new_n749), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n755), .A2(new_n473), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n555), .B2(new_n756), .ZN(G1336gat));
  NAND3_X1  g556(.A1(new_n753), .A2(new_n556), .A3(new_n489), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n489), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G92gat), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n758), .A2(new_n759), .B1(new_n761), .B2(KEYINPUT108), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n761), .A2(KEYINPUT108), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT52), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(KEYINPUT109), .A2(KEYINPUT52), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n758), .B(new_n765), .C1(new_n761), .C2(KEYINPUT52), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1337gat));
  AOI21_X1  g566(.A(G99gat), .B1(new_n753), .B2(new_n460), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n503), .A2(new_n560), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n768), .B1(new_n755), .B2(new_n769), .ZN(G1338gat));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n561), .A3(new_n471), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n755), .A2(new_n471), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n561), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g573(.A1(new_n619), .A2(new_n551), .A3(new_n639), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n635), .B1(new_n628), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n626), .A2(new_n627), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n629), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n626), .A2(new_n621), .A3(new_n627), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(KEYINPUT54), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n628), .A2(new_n778), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(KEYINPUT111), .A3(new_n783), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n780), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  OAI22_X1  g588(.A1(new_n789), .A2(KEYINPUT55), .B1(new_n548), .B2(new_n549), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n784), .A2(new_n785), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT111), .B1(new_n787), .B2(new_n783), .ZN(new_n792));
  OAI211_X1 g591(.A(KEYINPUT55), .B(new_n779), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n637), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n538), .A2(new_n542), .A3(new_n547), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n553), .A2(new_n531), .A3(new_n533), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n507), .B1(new_n796), .B2(new_n532), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n539), .A2(new_n541), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n546), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n790), .A2(new_n794), .B1(new_n730), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n584), .ZN(new_n802));
  INV_X1    g601(.A(new_n794), .ZN(new_n803));
  INV_X1    g602(.A(new_n800), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n789), .A2(KEYINPUT55), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n803), .A2(new_n583), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n618), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n777), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n473), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n810), .A2(new_n489), .A3(new_n383), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(new_n265), .A3(new_n551), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n808), .A2(new_n471), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n489), .A2(new_n424), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n460), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G113gat), .B1(new_n815), .B2(new_n550), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n812), .B1(new_n818), .B2(new_n819), .ZN(G1340gat));
  NOR3_X1   g619(.A1(new_n815), .A2(new_n267), .A3(new_n730), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n811), .A2(new_n639), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n822), .B2(new_n267), .ZN(G1341gat));
  INV_X1    g622(.A(new_n261), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n811), .A2(new_n824), .A3(new_n618), .ZN(new_n825));
  INV_X1    g624(.A(new_n618), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n261), .B1(new_n815), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT113), .Z(G1342gat));
  NAND4_X1  g628(.A1(new_n811), .A2(new_n258), .A3(new_n259), .A4(new_n583), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n830), .A2(KEYINPUT56), .ZN(new_n831));
  OAI21_X1  g630(.A(G134gat), .B1(new_n815), .B2(new_n584), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(KEYINPUT56), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(G1343gat));
  NAND2_X1  g633(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n835));
  OR3_X1    g634(.A1(new_n808), .A2(KEYINPUT115), .A3(new_n424), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n703), .A2(new_n489), .A3(new_n257), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n551), .A2(new_n203), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840));
  OAI22_X1  g639(.A1(new_n838), .A2(new_n839), .B1(KEYINPUT116), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n814), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n808), .B2(new_n257), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n257), .A2(new_n843), .ZN(new_n845));
  INV_X1    g644(.A(new_n806), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n583), .B1(new_n801), .B2(KEYINPUT114), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n848));
  OAI221_X1 g647(.A(new_n848), .B1(new_n730), .B2(new_n800), .C1(new_n790), .C2(new_n794), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n846), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n618), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n845), .B1(new_n777), .B2(new_n851), .ZN(new_n852));
  AOI211_X1 g651(.A(new_n703), .B(new_n842), .C1(new_n844), .C2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n203), .B1(new_n853), .B2(new_n551), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n840), .A2(KEYINPUT116), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT117), .Z(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  OR3_X1    g656(.A1(new_n841), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n841), .B2(new_n854), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1344gat));
  NAND2_X1  g659(.A1(new_n639), .A2(new_n204), .ZN(new_n861));
  OR3_X1    g660(.A1(new_n838), .A2(KEYINPUT118), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT118), .B1(new_n838), .B2(new_n861), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n703), .A2(new_n842), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n809), .A2(new_n845), .ZN(new_n867));
  INV_X1    g666(.A(new_n775), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n826), .B1(new_n850), .B2(KEYINPUT119), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n870));
  AOI211_X1 g669(.A(new_n870), .B(new_n846), .C1(new_n847), .C2(new_n849), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n868), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT57), .B1(new_n872), .B2(new_n471), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n867), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI211_X1 g674(.A(KEYINPUT120), .B(KEYINPUT57), .C1(new_n872), .C2(new_n471), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n639), .B(new_n866), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n204), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n873), .A2(new_n874), .ZN(new_n880));
  INV_X1    g679(.A(new_n876), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n881), .A3(new_n867), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n882), .A2(KEYINPUT121), .A3(new_n639), .A4(new_n866), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n865), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  AOI211_X1 g683(.A(KEYINPUT59), .B(new_n204), .C1(new_n853), .C2(new_n639), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n864), .B1(new_n884), .B2(new_n885), .ZN(G1345gat));
  INV_X1    g685(.A(new_n838), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n213), .A3(new_n618), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n853), .A2(new_n618), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n213), .ZN(G1346gat));
  NAND3_X1  g689(.A1(new_n887), .A2(new_n214), .A3(new_n583), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n853), .A2(new_n583), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n214), .ZN(G1347gat));
  NOR4_X1   g692(.A1(new_n808), .A2(new_n473), .A3(new_n694), .A4(new_n383), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n277), .A3(new_n551), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT122), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n694), .A2(new_n473), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n741), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT123), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n813), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n550), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n901), .ZN(G1348gat));
  OAI21_X1  g701(.A(G176gat), .B1(new_n900), .B2(new_n730), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n894), .A2(new_n278), .A3(new_n639), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1349gat));
  OAI211_X1 g704(.A(new_n894), .B(new_n618), .C1(new_n303), .C2(new_n302), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n295), .B1(new_n900), .B2(new_n826), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT60), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n909), .A2(KEYINPUT124), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n912), .B1(new_n908), .B2(KEYINPUT60), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT125), .B1(new_n909), .B2(new_n910), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n908), .A2(new_n915), .A3(KEYINPUT60), .ZN(new_n916));
  OAI22_X1  g715(.A1(new_n911), .A2(new_n913), .B1(new_n914), .B2(new_n916), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n894), .A2(new_n298), .A3(new_n583), .ZN(new_n918));
  OAI21_X1  g717(.A(G190gat), .B1(new_n900), .B2(new_n584), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1351gat));
  NAND3_X1  g721(.A1(new_n503), .A2(new_n489), .A3(new_n471), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n808), .A2(new_n473), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(KEYINPUT126), .B(G197gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n551), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n503), .A2(new_n897), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n882), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(new_n551), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n926), .B1(new_n930), .B2(new_n925), .ZN(G1352gat));
  NAND3_X1  g730(.A1(new_n924), .A2(new_n634), .A3(new_n639), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT62), .Z(new_n933));
  AND3_X1   g732(.A1(new_n882), .A2(new_n639), .A3(new_n928), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(new_n634), .ZN(G1353gat));
  NAND3_X1  g734(.A1(new_n882), .A2(new_n618), .A3(new_n928), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n607), .B1(KEYINPUT127), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT63), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n936), .B(new_n938), .C1(KEYINPUT127), .C2(new_n937), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n607), .A3(new_n618), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G1354gat));
  AOI21_X1  g743(.A(G218gat), .B1(new_n924), .B2(new_n583), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n583), .A2(G218gat), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n929), .B2(new_n946), .ZN(G1355gat));
endmodule


