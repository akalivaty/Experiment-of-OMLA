

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U322 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n416) );
  XNOR2_X1 U323 ( .A(n354), .B(n353), .ZN(n357) );
  XNOR2_X1 U324 ( .A(n352), .B(KEYINPUT94), .ZN(n353) );
  XOR2_X1 U325 ( .A(n572), .B(n458), .Z(n544) );
  XNOR2_X1 U326 ( .A(n449), .B(KEYINPUT38), .ZN(n497) );
  XOR2_X1 U327 ( .A(n473), .B(KEYINPUT28), .Z(n528) );
  XNOR2_X1 U328 ( .A(n362), .B(n422), .ZN(n515) );
  XOR2_X1 U329 ( .A(n350), .B(n349), .Z(n512) );
  XOR2_X1 U330 ( .A(G29GAT), .B(G43GAT), .Z(n290) );
  XNOR2_X1 U331 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n291) );
  XOR2_X1 U332 ( .A(G92GAT), .B(G64GAT), .Z(n292) );
  NOR2_X1 U333 ( .A1(n572), .A2(n455), .ZN(n456) );
  INV_X1 U334 ( .A(n515), .ZN(n469) );
  INV_X1 U335 ( .A(G197GAT), .ZN(n321) );
  OR2_X1 U336 ( .A1(n525), .A2(n469), .ZN(n471) );
  XNOR2_X1 U337 ( .A(n322), .B(n321), .ZN(n324) );
  XNOR2_X1 U338 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U339 ( .A(n324), .B(n323), .ZN(n351) );
  XNOR2_X1 U340 ( .A(n394), .B(n393), .ZN(n461) );
  XNOR2_X1 U341 ( .A(n468), .B(n291), .ZN(n525) );
  NAND2_X1 U342 ( .A1(n376), .A2(n375), .ZN(n480) );
  XNOR2_X1 U343 ( .A(n432), .B(n431), .ZN(n572) );
  XNOR2_X1 U344 ( .A(n417), .B(n416), .ZN(n511) );
  XNOR2_X1 U345 ( .A(G176GAT), .B(n361), .ZN(n422) );
  XOR2_X1 U346 ( .A(KEYINPUT124), .B(n568), .Z(n579) );
  NOR2_X1 U347 ( .A1(n476), .A2(n475), .ZN(n561) );
  XOR2_X1 U348 ( .A(n310), .B(n309), .Z(n526) );
  XNOR2_X1 U349 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n477) );
  XNOR2_X1 U350 ( .A(n450), .B(G43GAT), .ZN(n451) );
  XNOR2_X1 U351 ( .A(n478), .B(n477), .ZN(G1351GAT) );
  XNOR2_X1 U352 ( .A(n452), .B(n451), .ZN(G1330GAT) );
  XOR2_X1 U353 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n294) );
  XNOR2_X1 U354 ( .A(G99GAT), .B(KEYINPUT82), .ZN(n293) );
  XNOR2_X1 U355 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U356 ( .A(n295), .B(G190GAT), .Z(n297) );
  XOR2_X1 U357 ( .A(G15GAT), .B(G127GAT), .Z(n404) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(n404), .ZN(n296) );
  XNOR2_X1 U359 ( .A(n297), .B(n296), .ZN(n302) );
  XNOR2_X1 U360 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n298) );
  XOR2_X1 U361 ( .A(n298), .B(KEYINPUT81), .Z(n348) );
  XOR2_X1 U362 ( .A(G120GAT), .B(G71GAT), .Z(n428) );
  XNOR2_X1 U363 ( .A(n348), .B(n428), .ZN(n300) );
  NAND2_X1 U364 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U365 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U366 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U367 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n304) );
  XNOR2_X1 U368 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n303) );
  XNOR2_X1 U369 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U370 ( .A(KEYINPUT19), .B(n305), .Z(n359) );
  XOR2_X1 U371 ( .A(G176GAT), .B(KEYINPUT65), .Z(n307) );
  XNOR2_X1 U372 ( .A(G169GAT), .B(G113GAT), .ZN(n306) );
  XNOR2_X1 U373 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U374 ( .A(n359), .B(n308), .ZN(n309) );
  INV_X1 U375 ( .A(n526), .ZN(n476) );
  XOR2_X1 U376 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n312) );
  XNOR2_X1 U377 ( .A(KEYINPUT87), .B(KEYINPUT24), .ZN(n311) );
  XNOR2_X1 U378 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U379 ( .A(G204GAT), .B(KEYINPUT23), .Z(n314) );
  XOR2_X1 U380 ( .A(G141GAT), .B(G22GAT), .Z(n435) );
  XOR2_X1 U381 ( .A(G50GAT), .B(G162GAT), .Z(n384) );
  XNOR2_X1 U382 ( .A(n435), .B(n384), .ZN(n313) );
  XNOR2_X1 U383 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U384 ( .A(n316), .B(n315), .Z(n318) );
  NAND2_X1 U385 ( .A1(G228GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U386 ( .A(n318), .B(n317), .ZN(n320) );
  XNOR2_X1 U387 ( .A(G106GAT), .B(G78GAT), .ZN(n319) );
  XNOR2_X1 U388 ( .A(n319), .B(G148GAT), .ZN(n427) );
  XOR2_X1 U389 ( .A(n320), .B(n427), .Z(n328) );
  XNOR2_X1 U390 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n322) );
  XOR2_X1 U391 ( .A(KEYINPUT85), .B(G218GAT), .Z(n323) );
  XOR2_X1 U392 ( .A(G155GAT), .B(KEYINPUT86), .Z(n326) );
  XNOR2_X1 U393 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n325) );
  XNOR2_X1 U394 ( .A(n326), .B(n325), .ZN(n347) );
  XNOR2_X1 U395 ( .A(n351), .B(n347), .ZN(n327) );
  XNOR2_X1 U396 ( .A(n328), .B(n327), .ZN(n473) );
  XOR2_X1 U397 ( .A(G57GAT), .B(G127GAT), .Z(n330) );
  XNOR2_X1 U398 ( .A(G141GAT), .B(G120GAT), .ZN(n329) );
  XNOR2_X1 U399 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U400 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n332) );
  XNOR2_X1 U401 ( .A(KEYINPUT4), .B(KEYINPUT92), .ZN(n331) );
  XNOR2_X1 U402 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U403 ( .A(n334), .B(n333), .Z(n345) );
  XOR2_X1 U404 ( .A(KEYINPUT5), .B(KEYINPUT89), .Z(n336) );
  XNOR2_X1 U405 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n335) );
  XNOR2_X1 U406 ( .A(n336), .B(n335), .ZN(n343) );
  XOR2_X1 U407 ( .A(G113GAT), .B(G1GAT), .Z(n443) );
  XOR2_X1 U408 ( .A(G85GAT), .B(G162GAT), .Z(n338) );
  XNOR2_X1 U409 ( .A(G29GAT), .B(G148GAT), .ZN(n337) );
  XNOR2_X1 U410 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U411 ( .A(n443), .B(n339), .Z(n341) );
  NAND2_X1 U412 ( .A1(G225GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U413 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U414 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U415 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U416 ( .A(n347), .B(n346), .ZN(n350) );
  INV_X1 U417 ( .A(n348), .ZN(n349) );
  XOR2_X1 U418 ( .A(G169GAT), .B(G8GAT), .Z(n444) );
  XOR2_X1 U419 ( .A(n351), .B(n444), .Z(n354) );
  NAND2_X1 U420 ( .A1(G226GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U421 ( .A(G36GAT), .B(G190GAT), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n355), .B(KEYINPUT74), .ZN(n378) );
  XOR2_X1 U423 ( .A(n378), .B(KEYINPUT93), .Z(n356) );
  XNOR2_X1 U424 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U425 ( .A(n359), .B(n358), .ZN(n362) );
  XNOR2_X1 U426 ( .A(G204GAT), .B(KEYINPUT68), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n292), .B(n360), .ZN(n361) );
  XNOR2_X1 U428 ( .A(KEYINPUT27), .B(n515), .ZN(n368) );
  NAND2_X1 U429 ( .A1(n512), .A2(n368), .ZN(n363) );
  XOR2_X1 U430 ( .A(KEYINPUT95), .B(n363), .Z(n524) );
  NOR2_X1 U431 ( .A1(n528), .A2(n524), .ZN(n364) );
  NAND2_X1 U432 ( .A1(n476), .A2(n364), .ZN(n376) );
  NOR2_X1 U433 ( .A1(n473), .A2(n526), .ZN(n366) );
  XNOR2_X1 U434 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U436 ( .A(KEYINPUT96), .B(n367), .Z(n566) );
  NAND2_X1 U437 ( .A1(n368), .A2(n566), .ZN(n372) );
  NAND2_X1 U438 ( .A1(n526), .A2(n515), .ZN(n369) );
  NAND2_X1 U439 ( .A1(n473), .A2(n369), .ZN(n370) );
  XOR2_X1 U440 ( .A(KEYINPUT25), .B(n370), .Z(n371) );
  NAND2_X1 U441 ( .A1(n372), .A2(n371), .ZN(n374) );
  INV_X1 U442 ( .A(n512), .ZN(n373) );
  NAND2_X1 U443 ( .A1(n374), .A2(n373), .ZN(n375) );
  XNOR2_X1 U444 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n290), .B(n377), .ZN(n436) );
  XNOR2_X1 U446 ( .A(n436), .B(n378), .ZN(n383) );
  XOR2_X1 U447 ( .A(KEYINPUT75), .B(KEYINPUT71), .Z(n380) );
  NAND2_X1 U448 ( .A1(G232GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U449 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U450 ( .A(n381), .B(KEYINPUT10), .Z(n382) );
  XNOR2_X1 U451 ( .A(n383), .B(n382), .ZN(n388) );
  XOR2_X1 U452 ( .A(G99GAT), .B(G85GAT), .Z(n425) );
  XOR2_X1 U453 ( .A(n425), .B(G92GAT), .Z(n386) );
  XNOR2_X1 U454 ( .A(G106GAT), .B(n384), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U456 ( .A(n388), .B(n387), .Z(n394) );
  XOR2_X1 U457 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n390) );
  XNOR2_X1 U458 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n392) );
  XNOR2_X1 U460 ( .A(G134GAT), .B(G218GAT), .ZN(n391) );
  XOR2_X1 U461 ( .A(KEYINPUT36), .B(n461), .Z(n578) );
  NAND2_X1 U462 ( .A1(n480), .A2(n578), .ZN(n415) );
  XOR2_X1 U463 ( .A(G78GAT), .B(G155GAT), .Z(n396) );
  XNOR2_X1 U464 ( .A(G22GAT), .B(G211GAT), .ZN(n395) );
  XNOR2_X1 U465 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U466 ( .A(G64GAT), .B(G71GAT), .Z(n398) );
  XNOR2_X1 U467 ( .A(G8GAT), .B(G183GAT), .ZN(n397) );
  XNOR2_X1 U468 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U469 ( .A(n400), .B(n399), .Z(n406) );
  XOR2_X1 U470 ( .A(KEYINPUT13), .B(G57GAT), .Z(n421) );
  XOR2_X1 U471 ( .A(n421), .B(KEYINPUT80), .Z(n402) );
  NAND2_X1 U472 ( .A1(G231GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U473 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U474 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n414) );
  XOR2_X1 U476 ( .A(KEYINPUT79), .B(KEYINPUT77), .Z(n408) );
  XNOR2_X1 U477 ( .A(KEYINPUT12), .B(KEYINPUT78), .ZN(n407) );
  XNOR2_X1 U478 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U479 ( .A(KEYINPUT76), .B(KEYINPUT14), .Z(n410) );
  XNOR2_X1 U480 ( .A(G1GAT), .B(KEYINPUT15), .ZN(n409) );
  XNOR2_X1 U481 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U482 ( .A(n412), .B(n411), .Z(n413) );
  XOR2_X1 U483 ( .A(n414), .B(n413), .Z(n549) );
  INV_X1 U484 ( .A(n549), .ZN(n576) );
  NOR2_X1 U485 ( .A1(n415), .A2(n576), .ZN(n417) );
  XOR2_X1 U486 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n419) );
  NAND2_X1 U487 ( .A1(G230GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U488 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U489 ( .A(KEYINPUT32), .B(n420), .Z(n432) );
  XNOR2_X1 U490 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U491 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n423) );
  XNOR2_X1 U492 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U493 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U494 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U495 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U496 ( .A(G15GAT), .B(G197GAT), .Z(n434) );
  XNOR2_X1 U497 ( .A(G36GAT), .B(G50GAT), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n448) );
  XOR2_X1 U499 ( .A(n436), .B(n435), .Z(n438) );
  NAND2_X1 U500 ( .A1(G229GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U502 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n440) );
  XNOR2_X1 U503 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U505 ( .A(n442), .B(n441), .Z(n446) );
  XNOR2_X1 U506 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U507 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n569) );
  INV_X1 U509 ( .A(n569), .ZN(n542) );
  OR2_X1 U510 ( .A1(n572), .A2(n542), .ZN(n482) );
  NOR2_X1 U511 ( .A1(n511), .A2(n482), .ZN(n449) );
  NAND2_X1 U512 ( .A1(n497), .A2(n526), .ZN(n452) );
  XOR2_X1 U513 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n450) );
  NAND2_X1 U514 ( .A1(n576), .A2(n578), .ZN(n453) );
  XNOR2_X1 U515 ( .A(n453), .B(KEYINPUT113), .ZN(n454) );
  XOR2_X1 U516 ( .A(KEYINPUT45), .B(n454), .Z(n455) );
  XNOR2_X1 U517 ( .A(KEYINPUT114), .B(n456), .ZN(n457) );
  NAND2_X1 U518 ( .A1(n457), .A2(n542), .ZN(n467) );
  XOR2_X1 U519 ( .A(KEYINPUT64), .B(KEYINPUT41), .Z(n458) );
  NOR2_X1 U520 ( .A1(n542), .A2(n544), .ZN(n460) );
  INV_X1 U521 ( .A(KEYINPUT46), .ZN(n459) );
  XNOR2_X1 U522 ( .A(n460), .B(n459), .ZN(n463) );
  INV_X1 U523 ( .A(n461), .ZN(n536) );
  NOR2_X1 U524 ( .A1(n536), .A2(n576), .ZN(n462) );
  NAND2_X1 U525 ( .A1(n463), .A2(n462), .ZN(n465) );
  XOR2_X1 U526 ( .A(KEYINPUT47), .B(KEYINPUT112), .Z(n464) );
  XNOR2_X1 U527 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U528 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U529 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n470) );
  XNOR2_X1 U530 ( .A(n471), .B(n470), .ZN(n472) );
  NOR2_X1 U531 ( .A1(n472), .A2(n512), .ZN(n567) );
  NAND2_X1 U532 ( .A1(n473), .A2(n567), .ZN(n474) );
  XOR2_X1 U533 ( .A(KEYINPUT55), .B(n474), .Z(n475) );
  NAND2_X1 U534 ( .A1(n561), .A2(n536), .ZN(n478) );
  XOR2_X1 U535 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n485) );
  NOR2_X1 U536 ( .A1(n536), .A2(n549), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n479), .B(KEYINPUT16), .ZN(n481) );
  NAND2_X1 U538 ( .A1(n481), .A2(n480), .ZN(n500) );
  NOR2_X1 U539 ( .A1(n482), .A2(n500), .ZN(n483) );
  XNOR2_X1 U540 ( .A(KEYINPUT98), .B(n483), .ZN(n492) );
  NAND2_X1 U541 ( .A1(n492), .A2(n512), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U544 ( .A1(n492), .A2(n515), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n489) );
  NAND2_X1 U547 ( .A1(n492), .A2(n526), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(n491) );
  XOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT100), .Z(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  NAND2_X1 U551 ( .A1(n492), .A2(n528), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n493), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .Z(n495) );
  NAND2_X1 U554 ( .A1(n497), .A2(n512), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NAND2_X1 U556 ( .A1(n497), .A2(n515), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U558 ( .A1(n497), .A2(n528), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n498), .B(KEYINPUT104), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n502) );
  XNOR2_X1 U562 ( .A(KEYINPUT105), .B(n544), .ZN(n558) );
  NAND2_X1 U563 ( .A1(n542), .A2(n558), .ZN(n510) );
  NOR2_X1 U564 ( .A1(n500), .A2(n510), .ZN(n507) );
  NAND2_X1 U565 ( .A1(n507), .A2(n512), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n503), .Z(G1332GAT) );
  NAND2_X1 U568 ( .A1(n515), .A2(n507), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U570 ( .A(G71GAT), .B(KEYINPUT107), .Z(n506) );
  NAND2_X1 U571 ( .A1(n507), .A2(n526), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U574 ( .A1(n507), .A2(n528), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n514) );
  NOR2_X1 U577 ( .A1(n511), .A2(n510), .ZN(n519) );
  NAND2_X1 U578 ( .A1(n519), .A2(n512), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n515), .A2(n519), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U582 ( .A(G99GAT), .B(KEYINPUT109), .Z(n518) );
  NAND2_X1 U583 ( .A1(n519), .A2(n526), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(G1338GAT) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n523) );
  XOR2_X1 U586 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n521) );
  NAND2_X1 U587 ( .A1(n519), .A2(n528), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n541) );
  NAND2_X1 U591 ( .A1(n541), .A2(n526), .ZN(n527) );
  NOR2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n537), .A2(n569), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U596 ( .A1(n537), .A2(n558), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n535) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n533) );
  NAND2_X1 U600 ( .A1(n537), .A2(n576), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n539) );
  NAND2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n566), .A2(n541), .ZN(n551) );
  NOR2_X1 U608 ( .A1(n542), .A2(n551), .ZN(n543) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n543), .Z(G1344GAT) );
  NOR2_X1 U610 ( .A1(n551), .A2(n544), .ZN(n548) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n549), .A2(n551), .ZN(n550) );
  XOR2_X1 U616 ( .A(G155GAT), .B(n550), .Z(G1346GAT) );
  NOR2_X1 U617 ( .A1(n461), .A2(n551), .ZN(n552) );
  XOR2_X1 U618 ( .A(KEYINPUT120), .B(n552), .Z(n553) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(n553), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n561), .A2(n569), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(n554), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U625 ( .A(KEYINPUT122), .B(n557), .Z(n560) );
  NAND2_X1 U626 ( .A1(n558), .A2(n561), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U628 ( .A1(n576), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n564) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(n565), .Z(n571) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U635 ( .A1(n579), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n579), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U640 ( .A(n575), .B(G204GAT), .Z(G1353GAT) );
  NAND2_X1 U641 ( .A1(n579), .A2(n576), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n580), .B(KEYINPUT62), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

