//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT68), .Z(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(new_n453), .B2(G2106), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT69), .ZN(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT70), .Z(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT71), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(KEYINPUT71), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n469), .A2(new_n471), .A3(new_n465), .A4(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n466), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n475), .B1(new_n479), .B2(G2105), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n482));
  INV_X1    g057(.A(G136), .ZN(new_n483));
  INV_X1    g058(.A(G124), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n469), .A2(new_n471), .A3(G2105), .A4(new_n472), .ZN(new_n485));
  OAI221_X1 g060(.A(new_n482), .B1(new_n473), .B2(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XOR2_X1   g061(.A(KEYINPUT72), .B(KEYINPUT73), .Z(new_n487));
  OR2_X1    g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n487), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n465), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  OAI22_X1  g069(.A1(new_n485), .A2(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n473), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n476), .A2(new_n465), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT74), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n506), .A2(KEYINPUT75), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT75), .B1(new_n506), .B2(new_n507), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G88), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  OR3_X1    g088(.A1(new_n512), .A2(KEYINPUT76), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n507), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT76), .B1(new_n512), .B2(new_n513), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n511), .A2(new_n514), .A3(new_n517), .A4(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT77), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n515), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n510), .A2(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n521), .B1(new_n523), .B2(new_n515), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT77), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  AND3_X1   g107(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(G543), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n507), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n506), .A2(KEYINPUT75), .A3(new_n507), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT78), .B(G52), .Z(new_n543));
  OAI22_X1  g118(.A1(new_n542), .A2(new_n513), .B1(new_n515), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(G171));
  AOI22_X1  g120(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n513), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n548), .B2(new_n515), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(G81), .B2(new_n510), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT79), .ZN(G188));
  NAND3_X1  g131(.A1(new_n507), .A2(G53), .A3(G543), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT80), .ZN(new_n560));
  INV_X1    g135(.A(new_n506), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  INV_X1    g139(.A(G91), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n558), .B(new_n564), .C1(new_n565), .C2(new_n539), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  OR2_X1    g142(.A1(new_n506), .A2(G74), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n568), .A2(G651), .B1(new_n516), .B2(G49), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT81), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n539), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n510), .A2(KEYINPUT81), .A3(G87), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n510), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n561), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G48), .B2(new_n516), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n516), .A2(G47), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  OAI221_X1 g160(.A(new_n583), .B1(new_n513), .B2(new_n584), .C1(new_n539), .C2(new_n585), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(KEYINPUT82), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(KEYINPUT82), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(new_n516), .A2(G54), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT83), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(G66), .B2(new_n506), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n590), .B1(new_n594), .B2(new_n513), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(KEYINPUT10), .B1(new_n510), .B2(G92), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n537), .A2(KEYINPUT10), .A3(G92), .A4(new_n538), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n596), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n601), .B2(G171), .ZN(G284));
  OAI21_X1  g178(.A(new_n602), .B1(new_n601), .B2(G171), .ZN(G321));
  NAND2_X1  g179(.A1(G299), .A2(new_n601), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G168), .B2(new_n601), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(G168), .B2(new_n601), .ZN(G280));
  NAND3_X1  g182(.A1(new_n537), .A2(G92), .A3(new_n538), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n595), .B1(new_n610), .B2(new_n598), .ZN(new_n611));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G860), .ZN(G148));
  OAI21_X1  g188(.A(KEYINPUT84), .B1(new_n550), .B2(G868), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n600), .A2(G559), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n615), .A2(new_n601), .ZN(new_n616));
  MUX2_X1   g191(.A(new_n614), .B(KEYINPUT84), .S(new_n616), .Z(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n620));
  INV_X1    g195(.A(G123), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n485), .B2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n473), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G135), .ZN(new_n624));
  INV_X1    g199(.A(G2096), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT85), .B(G2100), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XOR2_X1   g205(.A(new_n628), .B(new_n630), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n624), .A2(new_n625), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n626), .A2(new_n631), .A3(new_n632), .ZN(G156));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n636), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n639), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(new_n647), .A3(G14), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT86), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n625), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1981), .B(G1986), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT87), .ZN(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n670), .A2(KEYINPUT88), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n670), .B2(KEYINPUT88), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT20), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n671), .A2(new_n677), .A3(new_n674), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n670), .A2(new_n673), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n668), .A2(new_n669), .ZN(new_n682));
  MUX2_X1   g257(.A(new_n673), .B(new_n681), .S(new_n682), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n679), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n680), .B1(new_n679), .B2(new_n683), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n666), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n686), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n688), .A2(new_n684), .A3(new_n665), .ZN(new_n689));
  XOR2_X1   g264(.A(G1991), .B(G1996), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n687), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n691), .B1(new_n687), .B2(new_n689), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n664), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n687), .A2(new_n689), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(new_n690), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n697), .A2(new_n663), .A3(new_n692), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  NAND2_X1  g275(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT94), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G6), .ZN(new_n705));
  INV_X1    g280(.A(G305), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n704), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT32), .B(G1981), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT92), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n704), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n704), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(G1971), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(G1971), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n710), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n704), .A2(G23), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n575), .B2(new_n704), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT33), .B(G1976), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT34), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n704), .A2(G24), .ZN(new_n722));
  INV_X1    g297(.A(G290), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n704), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT91), .ZN(new_n725));
  INV_X1    g300(.A(G1986), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G25), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT90), .Z(new_n730));
  AND2_X1   g305(.A1(new_n623), .A2(G131), .ZN(new_n731));
  INV_X1    g306(.A(G119), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n465), .A2(G107), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n485), .A2(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n730), .B1(new_n736), .B2(new_n728), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT35), .B(G1991), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  OR4_X1    g314(.A1(new_n703), .A2(new_n721), .A3(new_n727), .A4(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT25), .Z(new_n742));
  AOI22_X1  g317(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(new_n465), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G139), .B2(new_n623), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT96), .Z(new_n746));
  MUX2_X1   g321(.A(G33), .B(new_n746), .S(G29), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n728), .A2(G27), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n748), .A2(KEYINPUT100), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(KEYINPUT100), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n749), .B(new_n750), .C1(G164), .C2(new_n728), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n747), .A2(G2072), .B1(G2078), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G2072), .B2(new_n747), .ZN(new_n753));
  NOR2_X1   g328(.A1(G171), .A2(new_n704), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G5), .B2(new_n704), .ZN(new_n755));
  INV_X1    g330(.A(G1961), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT24), .ZN(new_n759));
  INV_X1    g334(.A(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G160), .B2(new_n728), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G2084), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n704), .A2(G20), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT23), .ZN(new_n766));
  INV_X1    g341(.A(G299), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(new_n704), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT101), .B(G1956), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n757), .A2(new_n758), .A3(new_n764), .A4(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(G11), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(G11), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n775), .A2(G28), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n728), .B1(new_n775), .B2(G28), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n773), .B(new_n774), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n624), .B2(G29), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n779), .B1(G2078), .B2(new_n751), .C1(new_n768), .C2(new_n769), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n753), .A2(new_n771), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n550), .A2(G16), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G16), .B2(G19), .ZN(new_n783));
  INV_X1    g358(.A(G1341), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n783), .A2(new_n784), .B1(G2084), .B2(new_n763), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n784), .B2(new_n783), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n704), .A2(G4), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n611), .B2(new_n704), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n786), .B1(G1348), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G1348), .B2(new_n788), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n728), .A2(G26), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT28), .Z(new_n792));
  OR2_X1    g367(.A1(G104), .A2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n794));
  INV_X1    g369(.A(G140), .ZN(new_n795));
  INV_X1    g370(.A(G128), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n794), .B1(new_n473), .B2(new_n795), .C1(new_n796), .C2(new_n485), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n792), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2067), .ZN(new_n803));
  OAI21_X1  g378(.A(KEYINPUT99), .B1(G16), .B2(G21), .ZN(new_n804));
  NOR2_X1   g379(.A1(G286), .A2(new_n704), .ZN(new_n805));
  MUX2_X1   g380(.A(new_n804), .B(KEYINPUT99), .S(new_n805), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1966), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n781), .A2(new_n790), .A3(new_n803), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n728), .A2(G35), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G162), .B2(new_n728), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT29), .B(G2090), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n728), .A2(G32), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n623), .A2(G141), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT97), .ZN(new_n815));
  NAND3_X1  g390(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT26), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT98), .ZN(new_n819));
  INV_X1    g394(.A(new_n485), .ZN(new_n820));
  AOI211_X1 g395(.A(new_n817), .B(new_n819), .C1(G129), .C2(new_n820), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n813), .B1(new_n822), .B2(new_n728), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT27), .ZN(new_n824));
  INV_X1    g399(.A(G1996), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n808), .A2(new_n812), .A3(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n727), .A2(new_n739), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n703), .B1(new_n828), .B2(new_n721), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n740), .A2(new_n827), .A3(new_n829), .ZN(G311));
  NAND3_X1  g405(.A1(new_n740), .A2(new_n827), .A3(new_n829), .ZN(G150));
  AOI22_X1  g406(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(new_n513), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n537), .A2(G93), .A3(new_n538), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT102), .B(G55), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n516), .A2(new_n835), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n834), .A2(KEYINPUT103), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(KEYINPUT103), .B1(new_n834), .B2(new_n836), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT104), .ZN(new_n840));
  INV_X1    g415(.A(new_n550), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT104), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n842), .B(new_n833), .C1(new_n837), .C2(new_n838), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n839), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n845), .A2(new_n842), .A3(new_n550), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n611), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n851));
  AOI21_X1  g426(.A(G860), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n839), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(G145));
  INV_X1    g431(.A(G37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n623), .A2(G142), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n820), .A2(G130), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n465), .A2(G118), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n858), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n630), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n736), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT107), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n801), .B(G164), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(new_n746), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n746), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n822), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n822), .B1(new_n867), .B2(new_n868), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n865), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n869), .A3(new_n864), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n490), .B(new_n624), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G160), .ZN(new_n876));
  XNOR2_X1  g451(.A(KEYINPUT105), .B(KEYINPUT106), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n872), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n865), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n869), .A3(new_n873), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(new_n872), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n857), .B(new_n879), .C1(new_n882), .C2(new_n878), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n885), .A2(KEYINPUT111), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n847), .B(new_n615), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT109), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n600), .B2(new_n767), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n611), .A2(KEYINPUT108), .A3(G299), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n600), .A2(new_n890), .A3(new_n767), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT108), .B1(new_n611), .B2(G299), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT109), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n611), .A2(G299), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n891), .A2(new_n892), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n897), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n900), .A2(new_n901), .B1(KEYINPUT41), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n898), .A2(KEYINPUT110), .A3(new_n899), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n888), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n887), .A2(new_n904), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n886), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n886), .ZN(new_n910));
  INV_X1    g485(.A(new_n908), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n905), .A2(new_n906), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n910), .B(new_n911), .C1(new_n912), .C2(new_n888), .ZN(new_n913));
  AOI21_X1  g488(.A(G305), .B1(new_n587), .B2(new_n588), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(G288), .A2(G166), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n575), .A2(G303), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n587), .A2(G305), .A3(new_n588), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n915), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n919), .ZN(new_n921));
  OAI22_X1  g496(.A1(new_n921), .A2(new_n914), .B1(new_n917), .B2(new_n916), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(KEYINPUT111), .B2(new_n885), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n909), .A2(new_n913), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n909), .B2(new_n913), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n839), .A2(new_n601), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(G295));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n928), .ZN(G331));
  NAND2_X1  g505(.A1(new_n900), .A2(new_n901), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n904), .A2(KEYINPUT41), .ZN(new_n932));
  XNOR2_X1  g507(.A(G286), .B(G171), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n847), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n844), .A2(new_n846), .A3(new_n933), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n931), .A2(new_n906), .A3(new_n932), .A4(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n904), .A3(new_n936), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n923), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n940), .A2(new_n857), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n923), .B1(new_n938), .B2(new_n939), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT43), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n844), .A2(new_n846), .A3(new_n933), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n933), .B1(new_n844), .B2(new_n846), .ZN(new_n946));
  OAI211_X1 g521(.A(KEYINPUT41), .B(new_n898), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n899), .B1(new_n935), .B2(new_n936), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n947), .B(new_n923), .C1(new_n948), .C2(new_n903), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT112), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT41), .B1(new_n945), .B2(new_n946), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n904), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n923), .A4(new_n947), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(new_n857), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n955), .A2(new_n956), .A3(new_n942), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT44), .B1(new_n944), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n956), .B1(new_n941), .B2(new_n943), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n955), .A2(KEYINPUT43), .A3(new_n942), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(G397));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(G164), .B2(G1384), .ZN(new_n965));
  NAND2_X1  g540(.A1(G160), .A2(G40), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n822), .B(G1996), .ZN(new_n969));
  INV_X1    g544(.A(G2067), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n801), .B(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n968), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT114), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n736), .B(new_n738), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n723), .A2(new_n726), .A3(new_n967), .ZN(new_n976));
  NAND3_X1  g551(.A1(G290), .A2(G1986), .A3(new_n967), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT113), .Z(new_n979));
  NOR2_X1   g554(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(G303), .A2(G8), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT55), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(G164), .B2(G1384), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n497), .A2(new_n499), .ZN(new_n986));
  INV_X1    g561(.A(new_n495), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(KEYINPUT115), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n983), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n966), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n988), .A2(new_n983), .A3(new_n989), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G2090), .ZN(new_n996));
  NOR2_X1   g571(.A1(G164), .A2(G1384), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n966), .B1(new_n997), .B2(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n965), .ZN(new_n999));
  INV_X1    g574(.A(G1971), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n995), .A2(new_n996), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n982), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n992), .A2(new_n985), .A3(new_n990), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n573), .A2(new_n574), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(G1976), .A3(new_n569), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1004), .A2(new_n1006), .A3(G8), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT52), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(KEYINPUT118), .A3(KEYINPUT52), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n575), .B2(G1976), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1004), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(new_n1002), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1016), .A2(new_n1018), .A3(new_n1006), .A4(new_n1019), .ZN(new_n1020));
  OR2_X1    g595(.A1(G305), .A2(G1981), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G305), .A2(G1981), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1021), .A2(KEYINPUT49), .A3(new_n1022), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1018), .A3(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1003), .A2(new_n1012), .A3(new_n1020), .A4(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n985), .A2(new_n990), .A3(new_n983), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n966), .A2(G2090), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1032), .A2(KEYINPUT116), .B1(new_n999), .B2(new_n1000), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1029), .A2(new_n1034), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1002), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n982), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT117), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1040), .A3(new_n1037), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1028), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1029), .A2(new_n1030), .A3(new_n992), .ZN(new_n1043));
  INV_X1    g618(.A(G2078), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n998), .A2(new_n1044), .A3(new_n965), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1043), .A2(new_n756), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT45), .B1(new_n985), .B2(new_n990), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n988), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n992), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1044), .A2(KEYINPUT53), .ZN(new_n1051));
  OR3_X1    g626(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(G301), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1966), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G2084), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1029), .A2(new_n1058), .A3(new_n1030), .A4(new_n992), .ZN(new_n1059));
  OAI211_X1 g634(.A(KEYINPUT120), .B(new_n1054), .C1(new_n1048), .C2(new_n1050), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1057), .A2(G168), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(G8), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1057), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1059), .ZN(new_n1066));
  OAI21_X1  g641(.A(G286), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(G8), .A3(new_n1061), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1064), .B1(KEYINPUT51), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT62), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1042), .B(new_n1053), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1061), .A2(G8), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1060), .A2(new_n1059), .ZN(new_n1073));
  AOI21_X1  g648(.A(G168), .B1(new_n1073), .B2(new_n1057), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT51), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1063), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(KEYINPUT62), .ZN(new_n1077));
  INV_X1    g652(.A(G1348), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1043), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1017), .A2(new_n970), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT121), .B(G1956), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n991), .B2(new_n994), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n992), .A2(new_n965), .A3(new_n1049), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT56), .B(G2072), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  XOR2_X1   g662(.A(G299), .B(KEYINPUT57), .Z(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1081), .A2(new_n1089), .A3(new_n611), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1088), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n611), .B1(new_n1081), .B2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1043), .A2(new_n1078), .B1(new_n1017), .B2(new_n970), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(KEYINPUT60), .A3(new_n600), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1096), .A2(new_n1098), .B1(new_n1095), .B2(new_n1081), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT58), .B(G1341), .Z(new_n1100));
  AOI22_X1  g675(.A1(new_n1085), .A2(new_n825), .B1(new_n1004), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n550), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT59), .B1(new_n1101), .B2(new_n841), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1084), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1088), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1093), .A2(KEYINPUT61), .A3(new_n1089), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1106), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1099), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1106), .A2(new_n1110), .A3(new_n1111), .A4(KEYINPUT122), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1094), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1043), .A2(new_n756), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1044), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n465), .B1(new_n479), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n477), .A2(KEYINPUT124), .A3(new_n478), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n475), .B(new_n1120), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(new_n965), .A3(new_n1049), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1118), .A2(new_n1119), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1126), .A2(G171), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1117), .B1(new_n1127), .B2(new_n1053), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1117), .B1(new_n1126), .B2(G171), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1052), .A2(new_n1118), .A3(new_n1119), .A4(G301), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1047), .A2(KEYINPUT125), .A3(G301), .A4(new_n1052), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1128), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1135), .A2(new_n1042), .A3(new_n1076), .ZN(new_n1136));
  OAI22_X1  g711(.A1(new_n1071), .A2(new_n1077), .B1(new_n1116), .B2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1012), .A2(new_n1020), .A3(new_n1027), .ZN(new_n1139));
  INV_X1    g714(.A(G1976), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1027), .A2(new_n1140), .A3(new_n575), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1021), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1138), .A2(new_n1139), .B1(new_n1018), .B2(new_n1142), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1002), .B(G286), .C1(new_n1073), .C2(new_n1057), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT63), .B1(new_n1042), .B2(new_n1144), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1139), .A2(new_n1146), .A3(KEYINPUT63), .A4(new_n1144), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1138), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1143), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n980), .B1(new_n1137), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n968), .B1(new_n971), .B2(new_n822), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n967), .A2(KEYINPUT46), .A3(new_n825), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT46), .B1(new_n967), .B2(new_n825), .ZN(new_n1153));
  OR3_X1    g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT47), .ZN(new_n1155));
  XOR2_X1   g730(.A(new_n976), .B(KEYINPUT48), .Z(new_n1156));
  OAI21_X1  g731(.A(new_n1155), .B1(new_n975), .B2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n731), .A2(new_n738), .A3(new_n735), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n973), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n799), .A2(new_n970), .A3(new_n800), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n968), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1150), .A2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g738(.A1(new_n960), .A2(new_n961), .ZN(new_n1165));
  NOR2_X1   g739(.A1(G227), .A2(new_n463), .ZN(new_n1166));
  NAND2_X1  g740(.A1(new_n648), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n1168));
  XNOR2_X1  g742(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  INV_X1    g743(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g744(.A(KEYINPUT127), .B1(new_n699), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n1172));
  AOI211_X1 g746(.A(new_n1172), .B(new_n1169), .C1(new_n695), .C2(new_n698), .ZN(new_n1173));
  OAI21_X1  g747(.A(new_n883), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g748(.A1(new_n1165), .A2(new_n1174), .ZN(G308));
  OAI221_X1 g749(.A(new_n883), .B1(new_n1171), .B2(new_n1173), .C1(new_n960), .C2(new_n961), .ZN(G225));
endmodule


