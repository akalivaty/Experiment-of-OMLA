

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797;

  INV_X1 U377 ( .A(G902), .ZN(n418) );
  XNOR2_X1 U378 ( .A(G113), .B(G104), .ZN(n516) );
  INV_X2 U379 ( .A(G953), .ZN(n772) );
  INV_X1 U380 ( .A(n551), .ZN(n658) );
  NOR2_X1 U381 ( .A1(n772), .A2(G952), .ZN(n706) );
  AND2_X2 U382 ( .A1(n438), .A2(n443), .ZN(n442) );
  AND2_X2 U383 ( .A1(n422), .A2(n421), .ZN(n420) );
  OR2_X2 U384 ( .A1(n428), .A2(n432), .ZN(n402) );
  AND2_X2 U385 ( .A1(n581), .A2(n580), .ZN(n594) );
  NAND2_X1 U386 ( .A1(n366), .A2(n762), .ZN(n378) );
  XNOR2_X2 U387 ( .A(n368), .B(KEYINPUT84), .ZN(n367) );
  INV_X1 U388 ( .A(n706), .ZN(n356) );
  NOR2_X1 U389 ( .A1(n590), .A2(n582), .ZN(n558) );
  AND2_X1 U390 ( .A1(n582), .A2(n590), .ZN(n583) );
  XNOR2_X1 U391 ( .A(n557), .B(KEYINPUT32), .ZN(n684) );
  INV_X1 U392 ( .A(n356), .ZN(n381) );
  INV_X1 U393 ( .A(n706), .ZN(n357) );
  INV_X1 U394 ( .A(KEYINPUT56), .ZN(n387) );
  INV_X1 U395 ( .A(KEYINPUT60), .ZN(n385) );
  XNOR2_X2 U396 ( .A(G107), .B(G104), .ZN(n450) );
  AND2_X1 U397 ( .A1(n377), .A2(n375), .ZN(n374) );
  NAND2_X1 U398 ( .A1(n379), .A2(n385), .ZN(n377) );
  AND2_X1 U399 ( .A1(n383), .A2(n371), .ZN(n370) );
  AND2_X1 U400 ( .A1(n762), .A2(G210), .ZN(n362) );
  AND2_X1 U401 ( .A1(n762), .A2(n384), .ZN(n359) );
  AND2_X1 U402 ( .A1(n762), .A2(G472), .ZN(n361) );
  AND2_X1 U403 ( .A1(n762), .A2(G217), .ZN(n358) );
  AND2_X1 U404 ( .A1(n762), .A2(G478), .ZN(n360) );
  XNOR2_X1 U405 ( .A(n614), .B(KEYINPUT40), .ZN(n796) );
  NOR2_X1 U406 ( .A1(n659), .A2(n662), .ZN(n632) );
  AND2_X1 U407 ( .A1(n380), .A2(n373), .ZN(n371) );
  NOR2_X1 U408 ( .A1(n382), .A2(n381), .ZN(n380) );
  AND2_X1 U409 ( .A1(n695), .A2(n385), .ZN(n376) );
  AND2_X1 U410 ( .A1(n386), .A2(G475), .ZN(n384) );
  NOR2_X1 U411 ( .A1(n386), .A2(G475), .ZN(n382) );
  INV_X1 U412 ( .A(n695), .ZN(n386) );
  XOR2_X1 U413 ( .A(KEYINPUT59), .B(n694), .Z(n695) );
  INV_X1 U414 ( .A(n385), .ZN(n373) );
  XNOR2_X1 U415 ( .A(KEYINPUT69), .B(G131), .ZN(n521) );
  XNOR2_X1 U416 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n458) );
  XNOR2_X1 U417 ( .A(G110), .B(G137), .ZN(n411) );
  XNOR2_X1 U418 ( .A(G119), .B(G128), .ZN(n460) );
  XNOR2_X1 U419 ( .A(KEYINPUT89), .B(KEYINPUT15), .ZN(n466) );
  XNOR2_X1 U420 ( .A(KEYINPUT71), .B(KEYINPUT16), .ZN(n481) );
  NAND2_X2 U421 ( .A1(n367), .A2(n666), .ZN(n366) );
  NAND2_X1 U422 ( .A1(n366), .A2(n358), .ZN(n365) );
  INV_X1 U423 ( .A(n378), .ZN(n363) );
  NAND2_X1 U424 ( .A1(n366), .A2(n359), .ZN(n383) );
  NAND2_X1 U425 ( .A1(n366), .A2(n360), .ZN(n677) );
  NAND2_X1 U426 ( .A1(n366), .A2(n361), .ZN(n680) );
  NAND2_X1 U427 ( .A1(n366), .A2(n362), .ZN(n705) );
  NAND2_X1 U428 ( .A1(n363), .A2(G469), .ZN(n700) );
  AND2_X1 U429 ( .A1(n364), .A2(n356), .ZN(G66) );
  XNOR2_X1 U430 ( .A(n365), .B(n674), .ZN(n364) );
  NAND2_X1 U431 ( .A1(n445), .A2(n444), .ZN(n368) );
  NAND2_X1 U432 ( .A1(n383), .A2(n380), .ZN(n379) );
  NAND2_X1 U433 ( .A1(n370), .A2(n369), .ZN(n372) );
  NAND2_X1 U434 ( .A1(n378), .A2(n695), .ZN(n369) );
  NAND2_X1 U435 ( .A1(n374), .A2(n372), .ZN(G60) );
  NAND2_X1 U436 ( .A1(n378), .A2(n376), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n388), .B(n387), .ZN(G51) );
  NAND2_X1 U438 ( .A1(n391), .A2(n356), .ZN(n388) );
  XNOR2_X1 U439 ( .A(n389), .B(KEYINPUT123), .ZN(G63) );
  NAND2_X1 U440 ( .A1(n395), .A2(n357), .ZN(n389) );
  XNOR2_X1 U441 ( .A(n390), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U442 ( .A1(n393), .A2(n357), .ZN(n390) );
  XNOR2_X1 U443 ( .A(n705), .B(n392), .ZN(n391) );
  INV_X1 U444 ( .A(n704), .ZN(n392) );
  XNOR2_X1 U445 ( .A(n680), .B(n394), .ZN(n393) );
  INV_X1 U446 ( .A(n679), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n677), .B(n396), .ZN(n395) );
  INV_X1 U448 ( .A(n676), .ZN(n396) );
  OR2_X2 U449 ( .A1(n548), .A2(n625), .ZN(n738) );
  NOR2_X1 U450 ( .A1(G902), .A2(G237), .ZN(n496) );
  INV_X1 U451 ( .A(G469), .ZN(n419) );
  NAND2_X1 U452 ( .A1(G902), .A2(G469), .ZN(n421) );
  NAND2_X1 U453 ( .A1(n738), .A2(KEYINPUT109), .ZN(n433) );
  INV_X1 U454 ( .A(KEYINPUT109), .ZN(n430) );
  XNOR2_X1 U455 ( .A(G116), .B(KEYINPUT7), .ZN(n528) );
  AND2_X1 U456 ( .A1(n573), .A2(n570), .ZN(n725) );
  XOR2_X1 U457 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n463) );
  AND2_X1 U458 ( .A1(n717), .A2(n629), .ZN(n631) );
  NAND2_X1 U459 ( .A1(n436), .A2(n435), .ZN(n748) );
  XOR2_X1 U460 ( .A(KEYINPUT105), .B(KEYINPUT9), .Z(n530) );
  XNOR2_X1 U461 ( .A(G107), .B(G122), .ZN(n529) );
  NAND2_X1 U462 ( .A1(n598), .A2(KEYINPUT85), .ZN(n443) );
  NAND2_X1 U463 ( .A1(n419), .A2(n418), .ZN(n417) );
  NOR2_X1 U464 ( .A1(G953), .A2(G237), .ZN(n513) );
  XNOR2_X1 U465 ( .A(G101), .B(KEYINPUT90), .ZN(n451) );
  AND2_X1 U466 ( .A1(n424), .A2(n683), .ZN(n667) );
  XNOR2_X1 U467 ( .A(n426), .B(n425), .ZN(n424) );
  INV_X1 U468 ( .A(KEYINPUT48), .ZN(n425) );
  NAND2_X1 U469 ( .A1(G234), .A2(G237), .ZN(n505) );
  XNOR2_X1 U470 ( .A(n501), .B(n500), .ZN(n611) );
  XNOR2_X1 U471 ( .A(n741), .B(n471), .ZN(n548) );
  XNOR2_X1 U472 ( .A(n460), .B(n458), .ZN(n409) );
  BUF_X1 U473 ( .A(n527), .Z(n537) );
  XNOR2_X1 U474 ( .A(G122), .B(G143), .ZN(n520) );
  XOR2_X1 U475 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n515) );
  XOR2_X1 U476 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n492) );
  NAND2_X1 U477 ( .A1(n667), .A2(n724), .ZN(n786) );
  INV_X1 U478 ( .A(KEYINPUT74), .ZN(n609) );
  XNOR2_X1 U479 ( .A(n468), .B(KEYINPUT25), .ZN(n406) );
  XNOR2_X1 U480 ( .A(n525), .B(n401), .ZN(n573) );
  XNOR2_X1 U481 ( .A(n524), .B(n526), .ZN(n401) );
  XOR2_X1 U482 ( .A(KEYINPUT122), .B(n675), .Z(n676) );
  INV_X2 U483 ( .A(n744), .ZN(n605) );
  XOR2_X1 U484 ( .A(KEYINPUT101), .B(G472), .Z(n397) );
  INV_X1 U485 ( .A(n605), .ZN(n435) );
  OR2_X1 U486 ( .A1(n604), .A2(n510), .ZN(n398) );
  AND2_X1 U487 ( .A1(n654), .A2(n653), .ZN(n399) );
  BUF_X1 U488 ( .A(n735), .Z(n765) );
  XNOR2_X1 U489 ( .A(n400), .B(n519), .ZN(n523) );
  XNOR2_X1 U490 ( .A(n518), .B(n522), .ZN(n400) );
  NAND2_X1 U491 ( .A1(n725), .A2(n549), .ZN(n404) );
  NAND2_X1 U492 ( .A1(n402), .A2(n630), .ZN(n480) );
  AND2_X1 U493 ( .A1(n584), .A2(KEYINPUT66), .ZN(n588) );
  NAND2_X2 U494 ( .A1(n420), .A2(n416), .ZN(n565) );
  XNOR2_X2 U495 ( .A(n403), .B(KEYINPUT22), .ZN(n412) );
  NOR2_X2 U496 ( .A1(n569), .A2(n404), .ZN(n403) );
  XNOR2_X2 U497 ( .A(n405), .B(KEYINPUT0), .ZN(n569) );
  NAND2_X1 U498 ( .A1(n511), .A2(n398), .ZN(n405) );
  XNOR2_X2 U499 ( .A(G146), .B(G125), .ZN(n486) );
  INV_X1 U500 ( .A(n738), .ZN(n431) );
  XNOR2_X2 U501 ( .A(n407), .B(n406), .ZN(n625) );
  NAND2_X1 U502 ( .A1(n674), .A2(n418), .ZN(n407) );
  XNOR2_X1 U503 ( .A(n470), .B(KEYINPUT21), .ZN(n741) );
  XNOR2_X1 U504 ( .A(n462), .B(n408), .ZN(n465) );
  XNOR2_X1 U505 ( .A(n410), .B(n409), .ZN(n408) );
  XNOR2_X1 U506 ( .A(n459), .B(n411), .ZN(n410) );
  NAND2_X1 U507 ( .A1(n412), .A2(n552), .ZN(n553) );
  NAND2_X1 U508 ( .A1(n412), .A2(n556), .ZN(n557) );
  NAND2_X1 U509 ( .A1(n576), .A2(n412), .ZN(n681) );
  XNOR2_X2 U510 ( .A(n413), .B(KEYINPUT19), .ZN(n511) );
  NAND2_X1 U511 ( .A1(n611), .A2(n726), .ZN(n413) );
  XNOR2_X2 U512 ( .A(n415), .B(n414), .ZN(n483) );
  XNOR2_X2 U513 ( .A(KEYINPUT3), .B(G119), .ZN(n414) );
  XNOR2_X2 U514 ( .A(G116), .B(G113), .ZN(n415) );
  XNOR2_X2 U515 ( .A(n565), .B(n457), .ZN(n550) );
  OR2_X1 U516 ( .A1(n696), .A2(n417), .ZN(n416) );
  NAND2_X1 U517 ( .A1(n696), .A2(G469), .ZN(n422) );
  XNOR2_X2 U518 ( .A(n477), .B(n456), .ZN(n696) );
  INV_X1 U519 ( .A(n786), .ZN(n444) );
  NAND2_X1 U520 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U521 ( .A1(n657), .A2(n656), .ZN(n426) );
  XNOR2_X2 U522 ( .A(n571), .B(KEYINPUT107), .ZN(n717) );
  XNOR2_X2 U523 ( .A(n605), .B(KEYINPUT6), .ZN(n630) );
  NAND2_X1 U524 ( .A1(n423), .A2(n727), .ZN(n613) );
  NAND2_X1 U525 ( .A1(n423), .A2(n640), .ZN(n682) );
  XNOR2_X1 U526 ( .A(n610), .B(n609), .ZN(n423) );
  XNOR2_X1 U527 ( .A(n427), .B(KEYINPUT30), .ZN(n606) );
  NAND2_X1 U528 ( .A1(n744), .A2(n726), .ZN(n427) );
  XNOR2_X2 U529 ( .A(n478), .B(n397), .ZN(n744) );
  OR2_X1 U530 ( .A1(n551), .A2(n738), .ZN(n437) );
  NOR2_X1 U531 ( .A1(n550), .A2(n429), .ZN(n428) );
  NAND2_X1 U532 ( .A1(n431), .A2(n430), .ZN(n429) );
  NAND2_X1 U533 ( .A1(n434), .A2(n433), .ZN(n432) );
  NAND2_X1 U534 ( .A1(n550), .A2(KEYINPUT109), .ZN(n434) );
  INV_X1 U535 ( .A(n437), .ZN(n436) );
  NAND2_X1 U536 ( .A1(n671), .A2(KEYINPUT85), .ZN(n438) );
  NAND2_X1 U537 ( .A1(n442), .A2(n439), .ZN(n445) );
  NAND2_X1 U538 ( .A1(n441), .A2(n440), .ZN(n439) );
  NOR2_X1 U539 ( .A1(n598), .A2(KEYINPUT85), .ZN(n440) );
  INV_X1 U540 ( .A(n671), .ZN(n441) );
  XOR2_X1 U541 ( .A(n639), .B(n540), .Z(n446) );
  AND2_X1 U542 ( .A1(n655), .A2(n399), .ZN(n656) );
  BUF_X1 U543 ( .A(n783), .Z(n785) );
  BUF_X1 U544 ( .A(n777), .Z(n778) );
  BUF_X1 U545 ( .A(n692), .Z(n693) );
  XNOR2_X2 U546 ( .A(G128), .B(KEYINPUT78), .ZN(n447) );
  XNOR2_X2 U547 ( .A(n447), .B(G143), .ZN(n488) );
  XNOR2_X2 U548 ( .A(n488), .B(G134), .ZN(n527) );
  XNOR2_X2 U549 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n487), .B(G137), .ZN(n448) );
  XNOR2_X1 U551 ( .A(n448), .B(n521), .ZN(n449) );
  XNOR2_X2 U552 ( .A(n527), .B(n449), .ZN(n783) );
  XNOR2_X2 U553 ( .A(n783), .B(G146), .ZN(n477) );
  XNOR2_X1 U554 ( .A(n450), .B(G110), .ZN(n452) );
  XNOR2_X1 U555 ( .A(n452), .B(n451), .ZN(n484) );
  XNOR2_X1 U556 ( .A(G140), .B(KEYINPUT97), .ZN(n454) );
  NAND2_X1 U557 ( .A1(n772), .A2(G227), .ZN(n453) );
  XNOR2_X1 U558 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U559 ( .A(n484), .B(n455), .ZN(n456) );
  INV_X1 U560 ( .A(KEYINPUT1), .ZN(n457) );
  XOR2_X1 U561 ( .A(KEYINPUT98), .B(KEYINPUT75), .Z(n459) );
  NAND2_X1 U562 ( .A1(G234), .A2(n772), .ZN(n461) );
  XOR2_X1 U563 ( .A(KEYINPUT8), .B(n461), .Z(n533) );
  NAND2_X1 U564 ( .A1(G221), .A2(n533), .ZN(n462) );
  XNOR2_X1 U565 ( .A(n486), .B(G140), .ZN(n464) );
  XNOR2_X1 U566 ( .A(n464), .B(n463), .ZN(n784) );
  XNOR2_X1 U567 ( .A(n465), .B(n784), .ZN(n674) );
  XNOR2_X1 U568 ( .A(n466), .B(n418), .ZN(n598) );
  NAND2_X1 U569 ( .A1(n598), .A2(G234), .ZN(n467) );
  XNOR2_X1 U570 ( .A(n467), .B(KEYINPUT20), .ZN(n469) );
  NAND2_X1 U571 ( .A1(G217), .A2(n469), .ZN(n468) );
  NAND2_X1 U572 ( .A1(n469), .A2(G221), .ZN(n470) );
  INV_X1 U573 ( .A(KEYINPUT99), .ZN(n471) );
  NAND2_X1 U574 ( .A1(n513), .A2(G210), .ZN(n472) );
  XNOR2_X1 U575 ( .A(n472), .B(KEYINPUT5), .ZN(n474) );
  XNOR2_X1 U576 ( .A(G101), .B(KEYINPUT100), .ZN(n473) );
  XNOR2_X1 U577 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U578 ( .A(n475), .B(n483), .ZN(n476) );
  XNOR2_X1 U579 ( .A(n477), .B(n476), .ZN(n678) );
  OR2_X2 U580 ( .A1(n678), .A2(G902), .ZN(n478) );
  INV_X1 U581 ( .A(KEYINPUT33), .ZN(n479) );
  XNOR2_X1 U582 ( .A(n480), .B(n479), .ZN(n735) );
  XNOR2_X1 U583 ( .A(n481), .B(G122), .ZN(n482) );
  XNOR2_X1 U584 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X1 U585 ( .A(n485), .B(n484), .ZN(n777) );
  XNOR2_X1 U586 ( .A(n487), .B(n486), .ZN(n489) );
  XNOR2_X1 U587 ( .A(n488), .B(n489), .ZN(n494) );
  NAND2_X1 U588 ( .A1(G224), .A2(n772), .ZN(n490) );
  XNOR2_X1 U589 ( .A(n490), .B(KEYINPUT91), .ZN(n491) );
  XNOR2_X1 U590 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U591 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U592 ( .A(n777), .B(n495), .ZN(n703) );
  INV_X1 U593 ( .A(n598), .ZN(n665) );
  NOR2_X1 U594 ( .A1(n703), .A2(n665), .ZN(n501) );
  XNOR2_X1 U595 ( .A(n496), .B(KEYINPUT73), .ZN(n502) );
  NAND2_X1 U596 ( .A1(n502), .A2(G210), .ZN(n499) );
  INV_X1 U597 ( .A(KEYINPUT79), .ZN(n497) );
  XNOR2_X1 U598 ( .A(n497), .B(KEYINPUT92), .ZN(n498) );
  XNOR2_X1 U599 ( .A(n499), .B(n498), .ZN(n500) );
  NAND2_X1 U600 ( .A1(n502), .A2(G214), .ZN(n504) );
  INV_X1 U601 ( .A(KEYINPUT93), .ZN(n503) );
  XNOR2_X1 U602 ( .A(n504), .B(n503), .ZN(n726) );
  XNOR2_X1 U603 ( .A(n505), .B(KEYINPUT94), .ZN(n506) );
  XNOR2_X1 U604 ( .A(KEYINPUT14), .B(n506), .ZN(n508) );
  NAND2_X1 U605 ( .A1(n508), .A2(G952), .ZN(n507) );
  XOR2_X1 U606 ( .A(KEYINPUT95), .B(n507), .Z(n758) );
  NOR2_X1 U607 ( .A1(n758), .A2(G953), .ZN(n604) );
  NAND2_X1 U608 ( .A1(G902), .A2(n508), .ZN(n600) );
  NOR2_X1 U609 ( .A1(G898), .A2(n772), .ZN(n509) );
  XOR2_X1 U610 ( .A(KEYINPUT96), .B(n509), .Z(n779) );
  NOR2_X1 U611 ( .A1(n600), .A2(n779), .ZN(n510) );
  NOR2_X2 U612 ( .A1(n735), .A2(n569), .ZN(n512) );
  XNOR2_X1 U613 ( .A(n512), .B(KEYINPUT34), .ZN(n541) );
  NAND2_X1 U614 ( .A1(G214), .A2(n513), .ZN(n514) );
  XNOR2_X1 U615 ( .A(n515), .B(n514), .ZN(n519) );
  XOR2_X1 U616 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n517) );
  XNOR2_X1 U617 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U618 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U619 ( .A(n523), .B(n784), .ZN(n694) );
  NOR2_X1 U620 ( .A1(G902), .A2(n694), .ZN(n525) );
  XNOR2_X1 U621 ( .A(KEYINPUT13), .B(KEYINPUT104), .ZN(n524) );
  INV_X1 U622 ( .A(G475), .ZN(n526) );
  XNOR2_X1 U623 ( .A(n528), .B(KEYINPUT106), .ZN(n532) );
  XNOR2_X1 U624 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U625 ( .A(n532), .B(n531), .Z(n535) );
  NAND2_X1 U626 ( .A1(G217), .A2(n533), .ZN(n534) );
  XNOR2_X1 U627 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U628 ( .A(n537), .B(n536), .ZN(n675) );
  NAND2_X1 U629 ( .A1(n675), .A2(n418), .ZN(n539) );
  INV_X1 U630 ( .A(G478), .ZN(n538) );
  XNOR2_X1 U631 ( .A(n539), .B(n538), .ZN(n570) );
  OR2_X1 U632 ( .A1(n573), .A2(n570), .ZN(n639) );
  INV_X1 U633 ( .A(KEYINPUT77), .ZN(n540) );
  NAND2_X1 U634 ( .A1(n541), .A2(n446), .ZN(n544) );
  INV_X1 U635 ( .A(KEYINPUT76), .ZN(n542) );
  XNOR2_X1 U636 ( .A(n542), .B(KEYINPUT35), .ZN(n543) );
  XNOR2_X2 U637 ( .A(n544), .B(n543), .ZN(n692) );
  INV_X1 U638 ( .A(n692), .ZN(n546) );
  INV_X1 U639 ( .A(KEYINPUT87), .ZN(n545) );
  NAND2_X1 U640 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U641 ( .A1(n547), .A2(KEYINPUT44), .ZN(n563) );
  INV_X1 U642 ( .A(n548), .ZN(n549) );
  BUF_X1 U643 ( .A(n550), .Z(n551) );
  AND2_X1 U644 ( .A1(n551), .A2(n605), .ZN(n552) );
  XNOR2_X1 U645 ( .A(n553), .B(KEYINPUT67), .ZN(n554) );
  NAND2_X1 U646 ( .A1(n554), .A2(n625), .ZN(n685) );
  XNOR2_X1 U647 ( .A(n625), .B(KEYINPUT108), .ZN(n740) );
  NAND2_X1 U648 ( .A1(n658), .A2(n740), .ZN(n555) );
  NOR2_X1 U649 ( .A1(n555), .A2(n630), .ZN(n556) );
  NAND2_X2 U650 ( .A1(n685), .A2(n684), .ZN(n590) );
  INV_X1 U651 ( .A(KEYINPUT88), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n692), .A2(n558), .ZN(n561) );
  NOR2_X1 U653 ( .A1(KEYINPUT44), .A2(KEYINPUT87), .ZN(n559) );
  AND2_X1 U654 ( .A1(n559), .A2(KEYINPUT66), .ZN(n560) );
  NAND2_X1 U655 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U656 ( .A1(n563), .A2(n562), .ZN(n581) );
  NAND2_X1 U657 ( .A1(n692), .A2(KEYINPUT87), .ZN(n579) );
  NOR2_X1 U658 ( .A1(n748), .A2(n569), .ZN(n564) );
  XNOR2_X1 U659 ( .A(n564), .B(KEYINPUT31), .ZN(n721) );
  INV_X1 U660 ( .A(n738), .ZN(n567) );
  BUF_X1 U661 ( .A(n565), .Z(n566) );
  AND2_X1 U662 ( .A1(n567), .A2(n566), .ZN(n599) );
  NAND2_X1 U663 ( .A1(n599), .A2(n605), .ZN(n568) );
  OR2_X1 U664 ( .A1(n569), .A2(n568), .ZN(n707) );
  NAND2_X1 U665 ( .A1(n721), .A2(n707), .ZN(n574) );
  INV_X1 U666 ( .A(n570), .ZN(n572) );
  OR2_X1 U667 ( .A1(n573), .A2(n572), .ZN(n571) );
  INV_X1 U668 ( .A(n717), .ZN(n720) );
  NAND2_X1 U669 ( .A1(n573), .A2(n572), .ZN(n686) );
  NAND2_X1 U670 ( .A1(n720), .A2(n686), .ZN(n730) );
  NAND2_X1 U671 ( .A1(n574), .A2(n730), .ZN(n577) );
  OR2_X1 U672 ( .A1(n658), .A2(n740), .ZN(n575) );
  NOR2_X1 U673 ( .A1(n575), .A2(n630), .ZN(n576) );
  AND2_X1 U674 ( .A1(n577), .A2(n681), .ZN(n578) );
  AND2_X1 U675 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U676 ( .A1(n692), .A2(n583), .ZN(n584) );
  INV_X1 U677 ( .A(n590), .ZN(n586) );
  INV_X1 U678 ( .A(KEYINPUT44), .ZN(n585) );
  OR2_X1 U679 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U680 ( .A1(n588), .A2(n587), .ZN(n592) );
  INV_X1 U681 ( .A(KEYINPUT66), .ZN(n589) );
  NAND2_X1 U682 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U683 ( .A1(n592), .A2(n591), .ZN(n593) );
  INV_X1 U684 ( .A(KEYINPUT64), .ZN(n595) );
  XNOR2_X1 U685 ( .A(n595), .B(KEYINPUT45), .ZN(n596) );
  XNOR2_X2 U686 ( .A(n597), .B(n596), .ZN(n671) );
  XNOR2_X1 U687 ( .A(n599), .B(KEYINPUT112), .ZN(n608) );
  NOR2_X1 U688 ( .A1(G900), .A2(n600), .ZN(n601) );
  NAND2_X1 U689 ( .A1(G953), .A2(n601), .ZN(n602) );
  XOR2_X1 U690 ( .A(KEYINPUT110), .B(n602), .Z(n603) );
  NOR2_X1 U691 ( .A1(n604), .A2(n603), .ZN(n616) );
  NOR2_X1 U692 ( .A1(n616), .A2(n606), .ZN(n607) );
  NAND2_X1 U693 ( .A1(n608), .A2(n607), .ZN(n610) );
  INV_X1 U694 ( .A(n611), .ZN(n662) );
  XNOR2_X1 U695 ( .A(KEYINPUT72), .B(KEYINPUT38), .ZN(n612) );
  XNOR2_X1 U696 ( .A(n662), .B(n612), .ZN(n727) );
  XNOR2_X1 U697 ( .A(n613), .B(KEYINPUT39), .ZN(n664) );
  NAND2_X1 U698 ( .A1(n664), .A2(n717), .ZN(n614) );
  AND2_X1 U699 ( .A1(n726), .A2(n727), .ZN(n731) );
  NAND2_X1 U700 ( .A1(n725), .A2(n731), .ZN(n615) );
  XOR2_X1 U701 ( .A(KEYINPUT41), .B(n615), .Z(n766) );
  INV_X1 U702 ( .A(n766), .ZN(n751) );
  NOR2_X1 U703 ( .A1(n741), .A2(n616), .ZN(n617) );
  XNOR2_X1 U704 ( .A(KEYINPUT70), .B(n617), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n618) );
  OR2_X1 U706 ( .A1(n605), .A2(n618), .ZN(n620) );
  INV_X1 U707 ( .A(KEYINPUT28), .ZN(n619) );
  XNOR2_X1 U708 ( .A(n620), .B(n619), .ZN(n621) );
  AND2_X1 U709 ( .A1(n621), .A2(n566), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n751), .A2(n636), .ZN(n622) );
  XNOR2_X1 U711 ( .A(n622), .B(KEYINPUT42), .ZN(n795) );
  NAND2_X1 U712 ( .A1(n796), .A2(n795), .ZN(n624) );
  XOR2_X1 U713 ( .A(KEYINPUT46), .B(KEYINPUT86), .Z(n623) );
  XNOR2_X1 U714 ( .A(n624), .B(n623), .ZN(n657) );
  INV_X1 U715 ( .A(n625), .ZN(n628) );
  NAND2_X1 U716 ( .A1(n626), .A2(n726), .ZN(n627) );
  NOR2_X1 U717 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U718 ( .A1(n631), .A2(n630), .ZN(n659) );
  XNOR2_X1 U719 ( .A(n632), .B(KEYINPUT36), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n633), .A2(n658), .ZN(n690) );
  INV_X1 U721 ( .A(n690), .ZN(n635) );
  INV_X1 U722 ( .A(n730), .ZN(n647) );
  NOR2_X1 U723 ( .A1(n647), .A2(KEYINPUT82), .ZN(n634) );
  NOR2_X1 U724 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U725 ( .A1(n636), .A2(n511), .ZN(n649) );
  INV_X1 U726 ( .A(n649), .ZN(n718) );
  NAND2_X1 U727 ( .A1(n718), .A2(KEYINPUT81), .ZN(n637) );
  NAND2_X1 U728 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U729 ( .A1(n639), .A2(n662), .ZN(n640) );
  XNOR2_X1 U730 ( .A(n682), .B(KEYINPUT83), .ZN(n641) );
  NOR2_X1 U731 ( .A1(n642), .A2(n641), .ZN(n655) );
  INV_X1 U732 ( .A(KEYINPUT47), .ZN(n646) );
  NOR2_X1 U733 ( .A1(n647), .A2(n649), .ZN(n643) );
  NOR2_X1 U734 ( .A1(KEYINPUT81), .A2(n643), .ZN(n644) );
  NAND2_X1 U735 ( .A1(n644), .A2(KEYINPUT82), .ZN(n645) );
  NAND2_X1 U736 ( .A1(n646), .A2(n645), .ZN(n654) );
  NAND2_X1 U737 ( .A1(KEYINPUT82), .A2(n647), .ZN(n651) );
  INV_X1 U738 ( .A(KEYINPUT81), .ZN(n648) );
  NAND2_X1 U739 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U740 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U741 ( .A1(n652), .A2(KEYINPUT47), .ZN(n653) );
  NOR2_X1 U742 ( .A1(n659), .A2(n658), .ZN(n661) );
  XNOR2_X1 U743 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n660) );
  XNOR2_X1 U744 ( .A(n661), .B(n660), .ZN(n663) );
  NAND2_X1 U745 ( .A1(n663), .A2(n662), .ZN(n683) );
  INV_X1 U746 ( .A(n686), .ZN(n714) );
  NAND2_X1 U747 ( .A1(n664), .A2(n714), .ZN(n724) );
  NAND2_X1 U748 ( .A1(n665), .A2(KEYINPUT2), .ZN(n666) );
  INV_X1 U749 ( .A(n667), .ZN(n670) );
  NAND2_X1 U750 ( .A1(n724), .A2(KEYINPUT2), .ZN(n668) );
  XNOR2_X1 U751 ( .A(n668), .B(KEYINPUT80), .ZN(n669) );
  NOR2_X1 U752 ( .A1(n670), .A2(n669), .ZN(n673) );
  BUF_X1 U753 ( .A(n671), .Z(n672) );
  NAND2_X1 U754 ( .A1(n673), .A2(n441), .ZN(n762) );
  XNOR2_X1 U755 ( .A(n678), .B(KEYINPUT62), .ZN(n679) );
  XNOR2_X1 U756 ( .A(n681), .B(G101), .ZN(G3) );
  XNOR2_X1 U757 ( .A(n682), .B(G143), .ZN(G45) );
  XNOR2_X1 U758 ( .A(n683), .B(G140), .ZN(G42) );
  XNOR2_X1 U759 ( .A(n684), .B(G119), .ZN(G21) );
  XNOR2_X1 U760 ( .A(n685), .B(G110), .ZN(G12) );
  NOR2_X1 U761 ( .A1(n721), .A2(n686), .ZN(n687) );
  XOR2_X1 U762 ( .A(G116), .B(n687), .Z(G18) );
  XOR2_X1 U763 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n689) );
  XNOR2_X1 U764 ( .A(G125), .B(KEYINPUT37), .ZN(n688) );
  XNOR2_X1 U765 ( .A(n689), .B(n688), .ZN(n691) );
  XOR2_X1 U766 ( .A(n691), .B(n690), .Z(G27) );
  XNOR2_X1 U767 ( .A(n693), .B(G122), .ZN(G24) );
  BUF_X1 U768 ( .A(n696), .Z(n698) );
  XOR2_X1 U769 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n697) );
  XNOR2_X1 U770 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U771 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U772 ( .A1(n701), .A2(n706), .ZN(G54) );
  XOR2_X1 U773 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n702) );
  XNOR2_X1 U774 ( .A(n703), .B(n702), .ZN(n704) );
  INV_X1 U775 ( .A(n707), .ZN(n709) );
  NAND2_X1 U776 ( .A1(n709), .A2(n717), .ZN(n708) );
  XNOR2_X1 U777 ( .A(n708), .B(G104), .ZN(G6) );
  XOR2_X1 U778 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n711) );
  NAND2_X1 U779 ( .A1(n709), .A2(n714), .ZN(n710) );
  XNOR2_X1 U780 ( .A(n711), .B(n710), .ZN(n713) );
  XOR2_X1 U781 ( .A(G107), .B(KEYINPUT27), .Z(n712) );
  XNOR2_X1 U782 ( .A(n713), .B(n712), .ZN(G9) );
  XOR2_X1 U783 ( .A(G128), .B(KEYINPUT29), .Z(n716) );
  NAND2_X1 U784 ( .A1(n718), .A2(n714), .ZN(n715) );
  XNOR2_X1 U785 ( .A(n716), .B(n715), .ZN(G30) );
  NAND2_X1 U786 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U787 ( .A(n719), .B(G146), .ZN(G48) );
  NOR2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U789 ( .A(KEYINPUT114), .B(n722), .Z(n723) );
  XNOR2_X1 U790 ( .A(G113), .B(n723), .ZN(G15) );
  XNOR2_X1 U791 ( .A(G134), .B(n724), .ZN(G36) );
  XNOR2_X1 U792 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n757) );
  INV_X1 U793 ( .A(n725), .ZN(n729) );
  NOR2_X1 U794 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U795 ( .A1(n729), .A2(n728), .ZN(n734) );
  NAND2_X1 U796 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U797 ( .A(KEYINPUT118), .B(n732), .Z(n733) );
  NOR2_X1 U798 ( .A1(n734), .A2(n733), .ZN(n736) );
  NOR2_X1 U799 ( .A1(n736), .A2(n765), .ZN(n737) );
  XNOR2_X1 U800 ( .A(n737), .B(KEYINPUT119), .ZN(n754) );
  NAND2_X1 U801 ( .A1(n551), .A2(n738), .ZN(n739) );
  XNOR2_X1 U802 ( .A(n739), .B(KEYINPUT50), .ZN(n747) );
  XOR2_X1 U803 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n743) );
  NAND2_X1 U804 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U805 ( .A(n743), .B(n742), .ZN(n745) );
  NOR2_X1 U806 ( .A1(n745), .A2(n435), .ZN(n746) );
  NAND2_X1 U807 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U808 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U809 ( .A(KEYINPUT51), .B(n750), .Z(n752) );
  NAND2_X1 U810 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U811 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U812 ( .A(n755), .B(KEYINPUT52), .ZN(n756) );
  XNOR2_X1 U813 ( .A(n757), .B(n756), .ZN(n759) );
  NOR2_X1 U814 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U815 ( .A1(G953), .A2(n760), .ZN(n770) );
  NOR2_X1 U816 ( .A1(n786), .A2(n672), .ZN(n761) );
  NOR2_X1 U817 ( .A1(n761), .A2(KEYINPUT2), .ZN(n764) );
  INV_X1 U818 ( .A(n762), .ZN(n763) );
  NOR2_X1 U819 ( .A1(n764), .A2(n763), .ZN(n768) );
  NOR2_X1 U820 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U821 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U822 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U823 ( .A(KEYINPUT53), .B(n771), .Z(G75) );
  NAND2_X1 U824 ( .A1(n441), .A2(n772), .ZN(n776) );
  NAND2_X1 U825 ( .A1(G953), .A2(G224), .ZN(n773) );
  XNOR2_X1 U826 ( .A(KEYINPUT61), .B(n773), .ZN(n774) );
  NAND2_X1 U827 ( .A1(n774), .A2(G898), .ZN(n775) );
  NAND2_X1 U828 ( .A1(n776), .A2(n775), .ZN(n782) );
  XNOR2_X1 U829 ( .A(n778), .B(KEYINPUT124), .ZN(n780) );
  NAND2_X1 U830 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U831 ( .A(n782), .B(n781), .Z(G69) );
  XOR2_X1 U832 ( .A(n785), .B(n784), .Z(n789) );
  XNOR2_X1 U833 ( .A(n786), .B(n789), .ZN(n787) );
  NOR2_X1 U834 ( .A1(G953), .A2(n787), .ZN(n788) );
  XNOR2_X1 U835 ( .A(n788), .B(KEYINPUT125), .ZN(n794) );
  XOR2_X1 U836 ( .A(G227), .B(n789), .Z(n790) );
  NAND2_X1 U837 ( .A1(n790), .A2(G900), .ZN(n791) );
  XNOR2_X1 U838 ( .A(KEYINPUT126), .B(n791), .ZN(n792) );
  NAND2_X1 U839 ( .A1(n792), .A2(G953), .ZN(n793) );
  NAND2_X1 U840 ( .A1(n794), .A2(n793), .ZN(G72) );
  XNOR2_X1 U841 ( .A(G137), .B(n795), .ZN(G39) );
  XOR2_X1 U842 ( .A(n796), .B(G131), .Z(n797) );
  XNOR2_X1 U843 ( .A(KEYINPUT127), .B(n797), .ZN(G33) );
endmodule

