//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  XNOR2_X1  g0002(.A(KEYINPUT65), .B(G77), .ZN(new_n203));
  AOI22_X1  g0003(.A1(new_n203), .A2(G244), .B1(G50), .B2(G226), .ZN(new_n204));
  INV_X1    g0004(.A(G68), .ZN(new_n205));
  XNOR2_X1  g0005(.A(KEYINPUT64), .B(G238), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI221_X1 g0008(.A(new_n204), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  OR2_X1    g0009(.A1(new_n209), .A2(KEYINPUT66), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G107), .A2(G264), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n209), .A2(KEYINPUT66), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT67), .Z(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G58), .B2(G232), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G20), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n217), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n219), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  INV_X1    g0034(.A(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n208), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G97), .B(G107), .ZN(new_n244));
  INV_X1    g0044(.A(G87), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n207), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G45), .ZN(new_n250));
  AOI21_X1  g0050(.A(G1), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(new_n249), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n252), .B1(new_n257), .B2(new_n222), .ZN(new_n258));
  INV_X1    g0058(.A(G238), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n255), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n257), .A2(new_n222), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n267));
  OAI21_X1  g0067(.A(G226), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n232), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n265), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G97), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n256), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n261), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT74), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(KEYINPUT74), .B(new_n261), .C1(new_n272), .C2(new_n274), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n260), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n279), .A2(KEYINPUT76), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT13), .B1(new_n279), .B2(KEYINPUT76), .ZN(new_n284));
  OAI211_X1 g0084(.A(G190), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n260), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT68), .B(G1698), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n270), .B1(new_n287), .B2(G226), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n288), .A2(new_n265), .B1(new_n256), .B2(new_n273), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT74), .B1(new_n289), .B2(new_n261), .ZN(new_n290));
  INV_X1    g0090(.A(new_n278), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n280), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n282), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G200), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n223), .A2(new_n256), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n223), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(G50), .A2(new_n297), .B1(new_n299), .B2(G77), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n223), .B2(G68), .ZN(new_n301));
  NAND3_X1  g0101(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n222), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(KEYINPUT11), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n303), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G1), .B2(new_n223), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n304), .B1(new_n205), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G1), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(G13), .A3(G20), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G68), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT12), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT11), .B1(new_n301), .B2(new_n303), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n307), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n285), .A2(new_n295), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT77), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n314), .B(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G87), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n262), .A2(new_n264), .A3(G226), .A4(G1698), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n262), .B(new_n264), .C1(new_n266), .C2(new_n267), .ZN(new_n319));
  INV_X1    g0119(.A(G223), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n317), .B(new_n318), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT81), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT3), .B(G33), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(new_n287), .A3(G223), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n325), .A2(KEYINPUT81), .A3(new_n317), .A4(new_n318), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(new_n261), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n258), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n254), .B1(new_n328), .B2(G232), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G200), .ZN(new_n331));
  INV_X1    g0131(.A(G58), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(new_n205), .ZN(new_n333));
  NOR2_X1   g0133(.A1(G58), .A2(G68), .ZN(new_n334));
  OAI21_X1  g0134(.A(G20), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G159), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n296), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n324), .B2(G20), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n337), .B1(new_n341), .B2(G68), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n305), .B1(new_n342), .B2(KEYINPUT16), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT80), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT80), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(new_n263), .A3(G33), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n348), .A3(new_n262), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n205), .B1(new_n350), .B2(new_n339), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n345), .B1(new_n351), .B2(new_n337), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT70), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT69), .B1(new_n354), .B2(new_n332), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT8), .ZN(new_n356));
  NAND2_X1  g0156(.A1(KEYINPUT8), .A2(G58), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n357), .A2(KEYINPUT69), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n306), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n309), .B2(new_n359), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n327), .A2(G190), .A3(new_n329), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n331), .A2(new_n353), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  OR2_X1    g0165(.A1(KEYINPUT82), .A2(KEYINPUT17), .ZN(new_n366));
  NAND2_X1  g0166(.A1(KEYINPUT82), .A2(KEYINPUT17), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n367), .B1(new_n365), .B2(new_n366), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT18), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n327), .A2(G179), .A3(new_n329), .ZN(new_n372));
  INV_X1    g0172(.A(G169), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n327), .B2(new_n329), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n362), .B1(new_n343), .B2(new_n352), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n371), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n330), .A2(G169), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n327), .A2(G179), .A3(new_n329), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n353), .A2(new_n363), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT18), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n265), .B1(G222), .B2(new_n287), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n320), .B2(new_n269), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n385), .B(new_n261), .C1(new_n203), .C2(new_n324), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n386), .B(new_n255), .C1(new_n235), .C2(new_n258), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n373), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n309), .A2(G50), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G50), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n306), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G150), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n296), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n223), .B1(new_n334), .B2(new_n391), .ZN(new_n396));
  AOI211_X1 g0196(.A(new_n395), .B(new_n396), .C1(new_n359), .C2(new_n299), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n390), .B(new_n393), .C1(new_n397), .C2(new_n305), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n388), .B(new_n398), .C1(G179), .C2(new_n387), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n370), .A2(new_n383), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n203), .A2(new_n309), .ZN(new_n401));
  INV_X1    g0201(.A(G77), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n306), .A2(new_n402), .ZN(new_n403));
  XOR2_X1   g0203(.A(KEYINPUT8), .B(G58), .Z(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n297), .ZN(new_n405));
  INV_X1    g0205(.A(new_n203), .ZN(new_n406));
  XOR2_X1   g0206(.A(KEYINPUT15), .B(G87), .Z(new_n407));
  INV_X1    g0207(.A(KEYINPUT72), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT15), .B(G87), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT72), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n405), .B1(new_n223), .B2(new_n406), .C1(new_n412), .C2(new_n298), .ZN(new_n413));
  AOI211_X1 g0213(.A(new_n401), .B(new_n403), .C1(new_n413), .C2(new_n303), .ZN(new_n414));
  INV_X1    g0214(.A(G107), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT71), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT71), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G107), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n265), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n324), .A2(G1698), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n420), .B1(new_n319), .B2(new_n232), .C1(new_n421), .C2(new_n206), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n261), .ZN(new_n423));
  INV_X1    g0223(.A(G244), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n423), .B(new_n255), .C1(new_n424), .C2(new_n258), .ZN(new_n425));
  OR3_X1    g0225(.A1(new_n425), .A2(KEYINPUT73), .A3(G179), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT73), .B1(new_n425), .B2(G179), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n414), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n373), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n425), .A2(G200), .ZN(new_n432));
  INV_X1    g0232(.A(G190), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n414), .C1(new_n433), .C2(new_n425), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n400), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(G179), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT14), .B1(new_n294), .B2(G169), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT14), .ZN(new_n439));
  AOI211_X1 g0239(.A(new_n439), .B(new_n373), .C1(new_n293), .C2(new_n282), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n437), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT78), .ZN(new_n442));
  INV_X1    g0242(.A(new_n313), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT78), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n437), .C1(new_n438), .C2(new_n440), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n398), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n447), .A2(KEYINPUT9), .B1(G200), .B2(new_n387), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT10), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n387), .A2(new_n433), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT9), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n398), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n396), .B1(new_n359), .B2(new_n299), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n394), .B2(new_n296), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n303), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(KEYINPUT9), .A3(new_n390), .A4(new_n393), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n387), .A2(G200), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n457), .A2(new_n452), .A3(new_n450), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT10), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  AND4_X1   g0261(.A1(new_n316), .A2(new_n436), .A3(new_n446), .A4(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(G257), .B1(new_n266), .B2(new_n267), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G264), .A2(G1698), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n324), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G303), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n265), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT88), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n466), .A2(KEYINPUT88), .A3(new_n468), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n261), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n308), .A2(G45), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT84), .B1(new_n475), .B2(G41), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT84), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(new_n249), .A3(KEYINPUT5), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n261), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI211_X1 g0282(.A(new_n474), .B(new_n480), .C1(new_n476), .C2(new_n478), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n482), .A2(G270), .B1(new_n483), .B2(G274), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n473), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n309), .A2(G116), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT89), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n488), .B(new_n223), .C1(G33), .C2(new_n273), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n305), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n207), .A2(G20), .ZN(new_n491));
  AOI21_X1  g0291(.A(G20), .B1(new_n256), .B2(G97), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(KEYINPUT89), .A3(new_n488), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n490), .A2(KEYINPUT20), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(new_n487), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n495), .A2(new_n493), .A3(new_n303), .A4(new_n491), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT20), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n486), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n308), .A2(G33), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n305), .A2(new_n309), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n207), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n485), .A2(new_n504), .A3(KEYINPUT90), .A4(G179), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT90), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n473), .A2(G179), .A3(new_n484), .ZN(new_n507));
  AOI211_X1 g0307(.A(new_n486), .B(new_n502), .C1(new_n494), .C2(new_n498), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n473), .A2(new_n484), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n504), .A2(new_n510), .A3(KEYINPUT21), .A4(G169), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n505), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT24), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n262), .A2(new_n264), .A3(G87), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n514), .A2(new_n515), .B1(G20), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT22), .A4(G87), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n520));
  AOI21_X1  g0320(.A(G20), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n419), .A2(KEYINPUT23), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n513), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n521), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(new_n523), .A3(new_n517), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(KEYINPUT24), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n303), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n501), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G107), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n309), .A2(G107), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n531), .B(KEYINPUT25), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n528), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n262), .A2(new_n264), .A3(G257), .A4(G1698), .ZN(new_n534));
  INV_X1    g0334(.A(G250), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n534), .B1(new_n319), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(G294), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n256), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n261), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n482), .A2(G264), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n483), .A2(G274), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n373), .ZN(new_n543));
  OR2_X1    g0343(.A1(new_n542), .A2(G179), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n533), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT21), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n510), .A2(G169), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n508), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n512), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT86), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT4), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n319), .B2(new_n424), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n324), .A2(G250), .A3(G1698), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n324), .A2(new_n287), .A3(KEYINPUT4), .A4(G244), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n553), .A2(new_n488), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n261), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n482), .A2(G257), .B1(new_n483), .B2(G274), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n557), .A2(KEYINPUT85), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT85), .B1(new_n557), .B2(new_n558), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n559), .A2(new_n560), .A3(G169), .ZN(new_n561));
  INV_X1    g0361(.A(G179), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n557), .A2(new_n562), .A3(new_n558), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n350), .A2(new_n339), .ZN(new_n564));
  XNOR2_X1  g0364(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n244), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n415), .A2(G97), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n564), .A2(new_n419), .B1(new_n568), .B2(G20), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n297), .A2(G77), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n305), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n309), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n273), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n501), .B2(new_n273), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n563), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n551), .B1(new_n561), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n557), .A2(new_n558), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT85), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n557), .A2(KEYINPUT85), .A3(new_n558), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n373), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n569), .A2(new_n570), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n303), .ZN(new_n583));
  INV_X1    g0383(.A(new_n574), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n581), .A2(new_n585), .A3(KEYINPUT86), .A4(new_n563), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n579), .A2(new_n580), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(G190), .B1(G200), .B2(new_n577), .ZN(new_n588));
  INV_X1    g0388(.A(new_n585), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n576), .A2(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(G87), .B1(new_n416), .B2(new_n418), .ZN(new_n591));
  NAND3_X1  g0391(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n591), .A2(new_n273), .B1(new_n223), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n298), .A2(new_n273), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n223), .A2(G68), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n594), .A2(KEYINPUT19), .B1(new_n265), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n303), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n412), .A2(new_n572), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n572), .A2(new_n303), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n409), .A2(new_n599), .A3(new_n411), .A4(new_n500), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(G33), .A2(G116), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n262), .A2(new_n264), .A3(G244), .A4(G1698), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n602), .B(new_n603), .C1(new_n319), .C2(new_n259), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n261), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n474), .A2(new_n253), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(G250), .B(new_n474), .C1(new_n257), .C2(new_n222), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n605), .A2(new_n562), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n608), .ZN(new_n610));
  AOI211_X1 g0410(.A(new_n606), .B(new_n610), .C1(new_n604), .C2(new_n261), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n601), .B(new_n609), .C1(new_n611), .C2(G169), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n605), .A2(G190), .A3(new_n607), .A4(new_n608), .ZN(new_n613));
  INV_X1    g0413(.A(G200), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT87), .B1(new_n529), .B2(G87), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT87), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n501), .A2(new_n617), .A3(new_n245), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n598), .B(new_n597), .C1(new_n616), .C2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n612), .B1(new_n615), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n542), .A2(new_n614), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n539), .A2(new_n540), .A3(new_n433), .A4(new_n541), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n528), .A2(new_n623), .A3(new_n530), .A4(new_n532), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT91), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n522), .A2(new_n513), .A3(new_n523), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n526), .A2(KEYINPUT24), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n628), .A2(new_n303), .B1(G107), .B2(new_n529), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT91), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n532), .A4(new_n623), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n620), .B1(new_n625), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n510), .A2(new_n433), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(G200), .B2(new_n510), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n508), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n550), .A2(new_n590), .A3(new_n632), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n463), .A2(new_n636), .ZN(G372));
  INV_X1    g0437(.A(KEYINPUT92), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n461), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n453), .A2(new_n460), .A3(KEYINPUT92), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n370), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n316), .A2(new_n431), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(new_n446), .ZN(new_n644));
  INV_X1    g0444(.A(new_n383), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n646), .A2(new_n399), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n590), .A2(new_n632), .A3(new_n549), .ZN(new_n648));
  NOR4_X1   g0448(.A1(new_n561), .A2(new_n620), .A3(new_n575), .A4(KEYINPUT26), .ZN(new_n649));
  INV_X1    g0449(.A(new_n620), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n576), .A2(new_n650), .A3(new_n586), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n649), .B1(new_n651), .B2(KEYINPUT26), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n648), .A2(new_n652), .A3(new_n612), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n647), .B1(new_n654), .B2(new_n463), .ZN(G369));
  INV_X1    g0455(.A(new_n635), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n512), .A2(new_n548), .ZN(new_n657));
  INV_X1    g0457(.A(G13), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(G20), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n308), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n508), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n657), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n657), .A2(new_n667), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n656), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g0470(.A(KEYINPUT93), .B(G330), .Z(new_n671));
  AND2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n625), .A2(new_n631), .B1(new_n533), .B2(new_n665), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n545), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n545), .A2(new_n665), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n673), .A2(new_n657), .A3(new_n545), .A4(new_n666), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n676), .A3(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n226), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G1), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n591), .A2(new_n273), .A3(new_n207), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n685), .A2(new_n686), .B1(new_n220), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n651), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT97), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n561), .A2(new_n575), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(KEYINPUT26), .A3(new_n650), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT97), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n651), .A2(new_n694), .A3(new_n689), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n648), .A2(new_n612), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .A3(new_n666), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n653), .A2(new_n666), .ZN(new_n700));
  XOR2_X1   g0500(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n507), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n611), .A2(new_n539), .A3(new_n540), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n703), .B(new_n704), .C1(new_n560), .C2(new_n559), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n587), .A2(KEYINPUT30), .A3(new_n703), .A4(new_n704), .ZN(new_n708));
  AOI21_X1  g0508(.A(G179), .B1(new_n473), .B2(new_n484), .ZN(new_n709));
  INV_X1    g0509(.A(new_n611), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(KEYINPUT94), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT94), .B1(new_n709), .B2(new_n710), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n577), .A2(new_n542), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n707), .B(new_n708), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT31), .B1(new_n716), .B2(new_n665), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT95), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n716), .A2(new_n665), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT95), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n590), .A2(new_n632), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(new_n550), .A3(new_n635), .A4(new_n666), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n719), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n699), .A2(new_n702), .B1(new_n728), .B2(new_n671), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n688), .B1(new_n729), .B2(G1), .ZN(G364));
  OR2_X1    g0530(.A1(new_n670), .A2(new_n671), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n670), .A2(new_n671), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n659), .A2(G45), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n733), .A2(KEYINPUT98), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(KEYINPUT98), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(G1), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n683), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n731), .A2(new_n732), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT99), .ZN(new_n740));
  NOR4_X1   g0540(.A1(new_n223), .A2(new_n433), .A3(new_n614), .A4(G179), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n433), .A2(G20), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT102), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n562), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n614), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n324), .B1(new_n245), .B2(new_n742), .C1(new_n747), .C2(new_n415), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT103), .Z(new_n749));
  NOR2_X1   g0549(.A1(new_n223), .A2(new_n562), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n433), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G190), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n752), .A2(G50), .B1(new_n755), .B2(new_n203), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n751), .A2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n433), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n223), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n756), .B1(new_n205), .B2(new_n758), .C1(new_n273), .C2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT32), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n745), .A2(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n762), .B1(new_n764), .B2(new_n336), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n763), .A2(KEYINPUT32), .A3(G159), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n761), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n750), .A2(G190), .A3(new_n614), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n749), .B(new_n767), .C1(new_n332), .C2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT104), .ZN(new_n770));
  INV_X1    g0570(.A(G283), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n747), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G317), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n758), .B1(KEYINPUT33), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(KEYINPUT33), .B2(new_n773), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n775), .B(new_n265), .C1(new_n467), .C2(new_n742), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n772), .B(new_n776), .C1(G329), .C2(new_n763), .ZN(new_n777));
  INV_X1    g0577(.A(new_n768), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G322), .ZN(new_n779));
  INV_X1    g0579(.A(new_n760), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT105), .B(G326), .Z(new_n781));
  AOI22_X1  g0581(.A1(G294), .A2(new_n780), .B1(new_n752), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(new_n754), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT106), .Z(new_n785));
  NAND3_X1  g0585(.A1(new_n777), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n770), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n222), .B1(G20), .B2(new_n373), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n738), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n243), .A2(G45), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n790), .A2(KEYINPUT100), .B1(new_n250), .B2(new_n221), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n682), .A2(new_n324), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n791), .B(new_n792), .C1(KEYINPUT100), .C2(new_n790), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n682), .A2(new_n265), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G355), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n793), .B(new_n795), .C1(G116), .C2(new_n226), .ZN(new_n796));
  OR3_X1    g0596(.A1(KEYINPUT101), .A2(G13), .A3(G33), .ZN(new_n797));
  OAI21_X1  g0597(.A(KEYINPUT101), .B1(G13), .B2(G33), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n788), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n796), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n801), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n789), .B(new_n803), .C1(new_n670), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n740), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  AND2_X1   g0608(.A1(new_n728), .A2(new_n671), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n430), .A2(new_n665), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n414), .A2(new_n666), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n428), .A2(new_n429), .B1(new_n434), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n700), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT108), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(KEYINPUT108), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n809), .A2(new_n814), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n816), .A2(new_n738), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n752), .A2(G137), .B1(new_n755), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G143), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n821), .B2(new_n768), .C1(new_n394), .C2(new_n758), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT34), .Z(new_n823));
  NOR2_X1   g0623(.A1(new_n747), .A2(new_n205), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n760), .A2(new_n332), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n324), .B1(new_n391), .B2(new_n742), .C1(new_n764), .C2(new_n826), .ZN(new_n827));
  NOR4_X1   g0627(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n245), .A2(new_n747), .B1(new_n764), .B2(new_n783), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n324), .B1(new_n778), .B2(G294), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n830), .B1(new_n415), .B2(new_n742), .C1(new_n207), .C2(new_n754), .ZN(new_n831));
  INV_X1    g0631(.A(new_n752), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(new_n467), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n758), .A2(new_n771), .B1(new_n273), .B2(new_n760), .ZN(new_n834));
  NOR4_X1   g0634(.A1(new_n829), .A2(new_n831), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n788), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n799), .A2(new_n788), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n836), .B1(G77), .B2(new_n838), .C1(new_n813), .C2(new_n800), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n738), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT107), .Z(new_n841));
  NAND2_X1  g0641(.A1(new_n819), .A2(new_n841), .ZN(G384));
  INV_X1    g0642(.A(KEYINPUT40), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n722), .B(new_n724), .C1(new_n636), .C2(new_n665), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n443), .A2(new_n665), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n446), .A2(new_n316), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(new_n446), .B2(new_n316), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n813), .B(new_n844), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT111), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n331), .A2(new_n353), .A3(new_n363), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n851), .A2(KEYINPUT82), .A3(KEYINPUT17), .A4(new_n364), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n383), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n342), .A2(new_n344), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n362), .B1(new_n854), .B2(new_n343), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n663), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n663), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n372), .A2(new_n374), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n365), .B1(new_n859), .B2(new_n855), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n861));
  XOR2_X1   g0661(.A(KEYINPUT110), .B(KEYINPUT37), .Z(new_n862));
  NAND2_X1  g0662(.A1(new_n380), .A2(new_n381), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n381), .A2(new_n858), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(new_n365), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n861), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n857), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n857), .B2(new_n866), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n849), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  INV_X1    g0670(.A(new_n856), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n370), .B2(new_n383), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n863), .A2(new_n864), .A3(new_n365), .ZN(new_n873));
  INV_X1    g0673(.A(new_n862), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n873), .A2(new_n874), .B1(KEYINPUT37), .B2(new_n860), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n870), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n857), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT111), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n869), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n843), .B1(new_n848), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n445), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n279), .A2(new_n281), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n280), .B(new_n260), .C1(new_n277), .C2(new_n278), .ZN(new_n883));
  OAI21_X1  g0683(.A(G169), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n439), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n294), .A2(KEYINPUT14), .A3(G169), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n444), .B1(new_n887), .B2(new_n437), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n314), .B(KEYINPUT77), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n443), .B(new_n665), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n446), .A2(new_n316), .A3(new_n845), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n864), .B1(new_n370), .B2(new_n383), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT112), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n874), .B1(new_n864), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n873), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n376), .A2(new_n663), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n862), .B1(new_n898), .B2(KEYINPUT112), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n865), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n870), .B1(new_n894), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n843), .B1(new_n902), .B2(new_n877), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n893), .A2(new_n813), .A3(new_n844), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n880), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n462), .A2(new_n844), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n905), .B(new_n906), .Z(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n671), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n699), .A2(new_n462), .A3(new_n702), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n647), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n653), .A2(new_n666), .A3(new_n813), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT109), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n810), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n893), .A2(new_n914), .A3(new_n869), .A4(new_n878), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n645), .A2(new_n663), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n446), .A2(new_n665), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n902), .A2(new_n877), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(new_n876), .B2(new_n877), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n915), .A2(new_n916), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n910), .B(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n908), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n308), .B2(new_n659), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n207), .B1(new_n568), .B2(KEYINPUT35), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(new_n224), .C1(KEYINPUT35), .C2(new_n568), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT36), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n203), .B1(new_n332), .B2(new_n205), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n929), .A2(new_n220), .B1(G50), .B2(new_n205), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(G1), .A3(new_n658), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n925), .A2(new_n928), .A3(new_n931), .ZN(G367));
  OAI221_X1 g0732(.A(new_n324), .B1(new_n754), .B2(new_n391), .C1(new_n394), .C2(new_n768), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n780), .A2(G68), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n758), .B2(new_n336), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n933), .B(new_n935), .C1(G58), .C2(new_n741), .ZN(new_n936));
  AOI22_X1  g0736(.A1(G137), .A2(new_n763), .B1(new_n746), .B2(new_n203), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n936), .B(new_n937), .C1(new_n821), .C2(new_n832), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT46), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n742), .B2(new_n207), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n940), .B1(new_n832), .B2(new_n783), .C1(new_n537), .C2(new_n758), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(G97), .B2(new_n746), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n741), .A2(KEYINPUT46), .A3(G116), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT115), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(KEYINPUT115), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n324), .B1(new_n755), .B2(G283), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G303), .B2(new_n778), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n942), .B(new_n948), .C1(new_n773), .C2(new_n764), .ZN(new_n949));
  INV_X1    g0749(.A(new_n419), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(new_n760), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n938), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(KEYINPUT116), .B(KEYINPUT47), .Z(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n738), .B1(new_n954), .B2(new_n788), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n619), .A2(new_n665), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n650), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n612), .B2(new_n956), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(new_n804), .ZN(new_n959));
  INV_X1    g0759(.A(new_n792), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n802), .B1(new_n226), .B2(new_n412), .C1(new_n239), .C2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n955), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n736), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n732), .A2(new_n677), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n680), .A2(new_n676), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n585), .A2(new_n665), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n590), .A2(new_n967), .B1(new_n692), .B2(new_n665), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n966), .A2(KEYINPUT44), .A3(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT44), .B1(new_n966), .B2(new_n968), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n966), .B2(new_n968), .ZN(new_n975));
  INV_X1    g0775(.A(new_n968), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n976), .A2(new_n676), .A3(new_n680), .A4(new_n973), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n965), .B1(new_n972), .B2(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n975), .A2(new_n977), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n966), .A2(new_n968), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n969), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n984), .A3(new_n679), .ZN(new_n985));
  INV_X1    g0785(.A(new_n680), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n675), .A2(new_n676), .B1(new_n657), .B2(new_n666), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n672), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n987), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n989), .A2(new_n732), .A3(new_n680), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n979), .A2(new_n729), .A3(new_n985), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n729), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n683), .B(KEYINPUT41), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT114), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT114), .ZN(new_n996));
  INV_X1    g0796(.A(new_n994), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(new_n992), .C2(new_n729), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n964), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n965), .A2(new_n976), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n968), .A2(new_n680), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT42), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n968), .A2(new_n545), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n576), .A2(new_n586), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n666), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1002), .B(new_n1010), .Z(new_n1011));
  AOI21_X1  g0811(.A(new_n963), .B1(new_n999), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT117), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI211_X1 g0814(.A(KEYINPUT117), .B(new_n963), .C1(new_n999), .C2(new_n1011), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(G387));
  NAND2_X1  g0817(.A1(new_n729), .A2(new_n991), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n683), .B(KEYINPUT119), .Z(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT120), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n729), .A2(new_n991), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1018), .A2(KEYINPUT120), .A3(new_n1020), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n991), .A2(new_n736), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n752), .A2(G322), .B1(new_n755), .B2(G303), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n783), .B2(new_n758), .C1(new_n773), .C2(new_n768), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT48), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n771), .B2(new_n760), .C1(new_n537), .C2(new_n742), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT49), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n324), .B1(new_n763), .B2(new_n781), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n207), .C2(new_n747), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n780), .A2(new_n409), .A3(new_n411), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n391), .B2(new_n768), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT118), .Z(new_n1037));
  NAND2_X1  g0837(.A1(new_n741), .A2(new_n203), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n763), .A2(G150), .B1(new_n359), .B2(new_n757), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n832), .A2(new_n336), .B1(new_n754), .B2(new_n205), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G97), .B2(new_n746), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1034), .B1(new_n265), .B2(new_n1042), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n236), .A2(new_n250), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1044), .A2(new_n792), .B1(new_n686), .B2(new_n794), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n404), .A2(new_n391), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT50), .Z(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n205), .B2(new_n402), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1048), .A2(G45), .A3(new_n686), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1045), .A2(new_n1049), .B1(G107), .B2(new_n226), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1043), .A2(new_n788), .B1(new_n802), .B2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n737), .C1(new_n678), .C2(new_n804), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1026), .A2(new_n1027), .A3(new_n1052), .ZN(G393));
  INV_X1    g0853(.A(KEYINPUT121), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n985), .A2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(new_n979), .Z(new_n1056));
  INV_X1    g0856(.A(new_n1018), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n992), .B(new_n1020), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n755), .A2(new_n404), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n402), .B2(new_n760), .C1(new_n758), .C2(new_n391), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT122), .Z(new_n1061));
  OAI22_X1  g0861(.A1(new_n832), .A2(new_n394), .B1(new_n336), .B2(new_n768), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT51), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n265), .B1(new_n741), .B2(G68), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G87), .A2(new_n746), .B1(new_n763), .B2(G143), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n324), .B1(new_n755), .B2(G294), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n207), .B2(new_n760), .C1(new_n758), .C2(new_n467), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n747), .A2(new_n415), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(G322), .C2(new_n763), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G317), .A2(new_n752), .B1(new_n778), .B2(G311), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT123), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT52), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(KEYINPUT52), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1070), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n742), .A2(new_n771), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1066), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n738), .B1(new_n1077), .B2(new_n788), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n976), .B2(new_n804), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n247), .A2(new_n792), .B1(G97), .B2(new_n682), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n802), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1056), .B2(new_n736), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1058), .A2(new_n1082), .ZN(G390));
  NAND3_X1  g0883(.A1(new_n728), .A2(new_n671), .A3(new_n813), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n846), .A2(new_n847), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n893), .A2(G330), .A3(new_n813), .A4(new_n844), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n914), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n893), .A2(new_n728), .A3(new_n671), .A4(new_n813), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n844), .A2(G330), .A3(new_n813), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1085), .A2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n810), .B(KEYINPUT109), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n665), .B1(new_n696), .B2(new_n697), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n813), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1090), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1089), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n462), .A2(G330), .A3(new_n844), .ZN(new_n1098));
  AND4_X1   g0898(.A1(new_n399), .A2(new_n909), .A3(new_n646), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1087), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n917), .B1(new_n877), .B2(new_n902), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1095), .B2(new_n1085), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n919), .A2(new_n920), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n892), .A2(new_n891), .B1(new_n911), .B2(new_n913), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1103), .B1(new_n1104), .B2(new_n917), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1100), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1090), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1102), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1097), .B(new_n1099), .C1(new_n1106), .C2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1086), .A2(new_n1087), .B1(new_n911), .B2(new_n913), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1096), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1099), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1087), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1102), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1109), .A2(new_n1116), .A3(new_n1020), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n359), .A2(new_n838), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT53), .B1(new_n742), .B2(new_n394), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n336), .B2(new_n760), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n757), .A2(G137), .ZN(new_n1121));
  INV_X1    g0921(.A(G128), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1121), .B1(new_n832), .B2(new_n1122), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n742), .A2(KEYINPUT53), .A3(new_n394), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n324), .B1(new_n768), .B2(new_n826), .ZN(new_n1125));
  NOR4_X1   g0925(.A1(new_n1120), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G50), .A2(new_n746), .B1(new_n763), .B2(G125), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1126), .B(new_n1127), .C1(new_n754), .C2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT124), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n824), .B1(G294), .B2(new_n763), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n758), .A2(new_n950), .B1(new_n402), .B2(new_n760), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n265), .B1(new_n207), .B2(new_n768), .C1(new_n742), .C2(new_n245), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(G97), .C2(new_n755), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1131), .B(new_n1134), .C1(new_n771), .C2(new_n832), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n788), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n737), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1118), .B(new_n1138), .C1(new_n1103), .C2(new_n799), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n736), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1117), .A2(new_n1141), .ZN(G378));
  INV_X1    g0942(.A(KEYINPUT57), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n880), .A2(G330), .A3(new_n904), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n922), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n639), .A2(new_n399), .A3(new_n640), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n447), .A2(new_n663), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1147), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n639), .A2(new_n399), .A3(new_n640), .A4(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(KEYINPUT55), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT55), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1148), .A2(new_n1153), .A3(new_n1150), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1152), .A2(KEYINPUT56), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT56), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n915), .A2(new_n916), .A3(new_n921), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1158), .A2(G330), .A3(new_n880), .A4(new_n904), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1145), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1157), .B1(new_n1145), .B2(new_n1159), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n647), .A2(new_n909), .A3(new_n1098), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1140), .B2(new_n1097), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1143), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1108), .A2(new_n1106), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1099), .B1(new_n1166), .B2(new_n1112), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1167), .B(KEYINPUT57), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1020), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n736), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1157), .A2(new_n799), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n752), .A2(G125), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n758), .B2(new_n826), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n778), .A2(G128), .B1(new_n755), .B2(G137), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n742), .B2(new_n1128), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(G150), .C2(new_n780), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT59), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G41), .B1(new_n763), .B2(G124), .ZN(new_n1178));
  AOI21_X1  g0978(.A(G33), .B1(new_n746), .B2(G159), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n249), .B1(new_n415), .B2(new_n768), .C1(new_n412), .C2(new_n754), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n752), .A2(G116), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n757), .A2(G97), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n934), .A2(new_n1182), .A3(new_n1183), .A4(new_n1038), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1181), .A2(new_n1184), .A3(new_n324), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n332), .B2(new_n747), .C1(new_n771), .C2(new_n764), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT58), .ZN(new_n1187));
  AOI21_X1  g0987(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1180), .B(new_n1187), .C1(G50), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n738), .B1(new_n1189), .B2(new_n788), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1171), .B(new_n1190), .C1(G50), .C2(new_n838), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1170), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1169), .A2(new_n1193), .ZN(G375));
  NAND3_X1  g0994(.A1(new_n1089), .A2(new_n1163), .A3(new_n1096), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1195), .A2(new_n1112), .A3(new_n994), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT125), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n758), .A2(new_n1128), .B1(new_n391), .B2(new_n760), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n324), .B1(new_n394), .B2(new_n754), .C1(new_n742), .C2(new_n336), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(G137), .C2(new_n778), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G58), .A2(new_n746), .B1(new_n763), .B2(G128), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n826), .C2(new_n832), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G77), .A2(new_n746), .B1(new_n763), .B2(G303), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n757), .A2(G116), .B1(new_n752), .B2(G294), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n265), .B1(new_n742), .B2(new_n273), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n419), .B2(new_n755), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1203), .A2(new_n1035), .A3(new_n1204), .A4(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n768), .A2(new_n771), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1202), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n788), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(G68), .B2(new_n838), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n738), .B(new_n1211), .C1(new_n1085), .C2(new_n799), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1097), .B2(new_n736), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1197), .A2(new_n1213), .ZN(G381));
  INV_X1    g1014(.A(G384), .ZN(new_n1215));
  INV_X1    g1015(.A(G390), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1016), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AND4_X1   g1017(.A1(new_n1141), .A2(new_n1117), .A3(new_n1170), .A4(new_n1191), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1169), .A2(new_n1218), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1026), .A2(new_n807), .A3(new_n1027), .A4(new_n1052), .ZN(new_n1220));
  OR4_X1    g1020(.A1(G381), .A2(new_n1217), .A3(new_n1219), .A4(new_n1220), .ZN(G407));
  OAI211_X1 g1021(.A(G407), .B(G213), .C1(G343), .C2(new_n1219), .ZN(G409));
  AND2_X1   g1022(.A1(new_n664), .A2(G213), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1167), .B(new_n994), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1218), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1167), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1019), .B1(new_n1226), .B2(new_n1143), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1192), .B1(new_n1227), .B2(new_n1168), .ZN(new_n1228));
  INV_X1    g1028(.A(G378), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1225), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT60), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1195), .A2(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1089), .A2(new_n1163), .A3(KEYINPUT60), .A4(new_n1096), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1232), .A2(new_n1020), .A3(new_n1112), .A4(new_n1233), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1234), .A2(G384), .A3(new_n1213), .ZN(new_n1235));
  AOI21_X1  g1035(.A(G384), .B1(new_n1234), .B2(new_n1213), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G2897), .B(new_n1223), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(new_n1213), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1215), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1234), .A2(G384), .A3(new_n1213), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1223), .A2(G2897), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1237), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT61), .B1(new_n1230), .B2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1225), .B(new_n1245), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT62), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1229), .B1(new_n1169), .B2(new_n1193), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT62), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n1225), .A4(new_n1245), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1244), .A2(new_n1247), .A3(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1216), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G393), .A2(G396), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1012), .A2(G390), .B1(new_n1220), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n999), .A2(new_n1011), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n962), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1216), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1012), .A2(G390), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1254), .A2(KEYINPUT126), .A3(new_n1220), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT126), .B1(new_n1254), .B2(new_n1220), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1253), .A2(new_n1255), .B1(new_n1260), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1252), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(KEYINPUT61), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1249), .A2(KEYINPUT63), .A3(new_n1225), .A4(new_n1245), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1246), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT63), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1230), .B2(new_n1243), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1266), .B(new_n1267), .C1(new_n1268), .C2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1265), .A2(new_n1271), .ZN(G405));
  INV_X1    g1072(.A(new_n1245), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1117), .A2(new_n1170), .A3(new_n1141), .A4(new_n1191), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1227), .B2(new_n1168), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1248), .B2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1245), .B(new_n1219), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT127), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1278), .A2(new_n1279), .A3(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1279), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(G402));
endmodule


