//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n189), .B2(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n187), .A2(KEYINPUT23), .A3(G119), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n190), .A3(new_n196), .ZN(new_n197));
  OR2_X1    g011(.A1(new_n197), .A2(KEYINPUT73), .ZN(new_n198));
  INV_X1    g012(.A(G110), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n199), .B1(new_n197), .B2(KEYINPUT73), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n193), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT16), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT74), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT74), .A4(KEYINPUT16), .ZN(new_n209));
  INV_X1    g023(.A(new_n203), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AND4_X1   g026(.A1(G146), .A2(new_n208), .A3(new_n209), .A4(new_n212), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n206), .A2(new_n207), .B1(new_n211), .B2(new_n210), .ZN(new_n214));
  AOI21_X1  g028(.A(G146), .B1(new_n214), .B2(new_n209), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n201), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n203), .A2(new_n205), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G146), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n197), .A2(G110), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n191), .A2(new_n192), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n214), .A2(G146), .A3(new_n209), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT75), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT75), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n216), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G953), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(G221), .A3(G234), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n229), .B(KEYINPUT22), .ZN(new_n230));
  INV_X1    g044(.A(G137), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n230), .B(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n225), .A2(new_n227), .A3(new_n232), .ZN(new_n233));
  OR2_X1    g047(.A1(new_n224), .A2(new_n232), .ZN(new_n234));
  INV_X1    g048(.A(G217), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(G234), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G902), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n234), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT77), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n233), .A2(KEYINPUT77), .A3(new_n234), .A4(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n233), .A2(new_n236), .A3(new_n234), .A4(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n237), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n233), .A2(new_n236), .A3(new_n234), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(new_n244), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n243), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G475), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n213), .A2(new_n215), .ZN(new_n253));
  NOR2_X1   g067(.A1(G237), .A2(G953), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G214), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(G143), .A2(G214), .ZN(new_n258));
  AOI21_X1  g072(.A(G131), .B1(new_n258), .B2(new_n254), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G237), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n261), .A2(new_n228), .A3(G143), .A4(G214), .ZN(new_n262));
  INV_X1    g076(.A(G214), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n263), .A2(G237), .A3(G953), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n262), .B1(new_n264), .B2(G143), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n260), .A2(KEYINPUT89), .B1(new_n265), .B2(G131), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT17), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT89), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n257), .A2(new_n268), .A3(new_n259), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n266), .A2(KEYINPUT92), .A3(new_n267), .A4(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G131), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(G143), .B1(new_n254), .B2(G214), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT89), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(G143), .A2(G214), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n275), .A2(G237), .A3(G953), .ZN(new_n276));
  OAI21_X1  g090(.A(G131), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n274), .A2(new_n269), .A3(new_n267), .A4(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT92), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n265), .A2(KEYINPUT17), .A3(G131), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n253), .A2(new_n270), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(KEYINPUT18), .A2(G131), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n265), .B(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n217), .A2(KEYINPUT88), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT88), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n203), .A2(new_n205), .A3(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n285), .A2(G146), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n288), .B2(new_n218), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(G113), .B(G122), .ZN(new_n291));
  INV_X1    g105(.A(G104), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT93), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n282), .A2(new_n293), .A3(new_n289), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n293), .B1(new_n282), .B2(new_n289), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n299), .B2(KEYINPUT93), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n252), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(G475), .A2(G902), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n285), .A2(KEYINPUT19), .A3(new_n287), .ZN(new_n303));
  INV_X1    g117(.A(G146), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n217), .A2(KEYINPUT19), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT90), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n266), .A2(new_n269), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT90), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n303), .A2(new_n309), .A3(new_n304), .A4(new_n305), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n307), .A2(new_n222), .A3(new_n308), .A4(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n293), .B1(new_n311), .B2(new_n289), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n297), .B1(new_n312), .B2(KEYINPUT91), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT91), .ZN(new_n314));
  AOI211_X1 g128(.A(new_n314), .B(new_n293), .C1(new_n311), .C2(new_n289), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n302), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT20), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT20), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n318), .B(new_n302), .C1(new_n313), .C2(new_n315), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n301), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT9), .B(G234), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n321), .A2(new_n235), .A3(G953), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT94), .B1(new_n187), .B2(G143), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT94), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n256), .A3(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G134), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n187), .A2(G143), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT95), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT95), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n327), .A2(new_n332), .A3(new_n328), .A4(new_n329), .ZN(new_n333));
  INV_X1    g147(.A(G116), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G122), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G107), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(G122), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G122), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(G116), .ZN(new_n341));
  OAI21_X1  g155(.A(G107), .B1(new_n341), .B2(new_n335), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n331), .A2(new_n333), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT13), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n329), .B1(new_n327), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT13), .B1(new_n324), .B2(new_n326), .ZN(new_n347));
  OAI21_X1  g161(.A(G134), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT96), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(new_n338), .C1(new_n335), .C2(KEYINPUT14), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT14), .B1(new_n340), .B2(G116), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(new_n341), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT96), .B1(new_n338), .B2(KEYINPUT14), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n350), .B(G107), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n330), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n328), .B1(new_n327), .B2(new_n329), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n354), .B(new_n339), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT97), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n339), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n337), .B1(new_n352), .B2(new_n349), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n338), .A2(KEYINPUT14), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n338), .B1(new_n335), .B2(KEYINPUT14), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT96), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n360), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n327), .A2(new_n329), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G134), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n330), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n365), .A2(KEYINPUT97), .A3(new_n368), .ZN(new_n369));
  AOI221_X4 g183(.A(new_n323), .B1(new_n344), .B2(new_n348), .C1(new_n359), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n359), .A2(new_n369), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n344), .A2(new_n348), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n322), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n236), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G478), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT15), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(KEYINPUT98), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n357), .A2(new_n358), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT97), .B1(new_n365), .B2(new_n368), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n372), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n323), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n371), .A2(new_n322), .A3(new_n372), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT98), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(new_n236), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n377), .B1(new_n387), .B2(new_n376), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n228), .A2(G952), .ZN(new_n389));
  INV_X1    g203(.A(G234), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n389), .B1(new_n390), .B2(new_n261), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AOI211_X1 g206(.A(new_n236), .B(new_n228), .C1(G234), .C2(G237), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT21), .B(G898), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n320), .A2(new_n388), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G214), .B1(G237), .B2(G902), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G210), .B1(G237), .B2(G902), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT85), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n304), .A2(G143), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n256), .A2(G146), .ZN(new_n404));
  AND4_X1   g218(.A1(KEYINPUT0), .A2(new_n403), .A3(new_n404), .A4(G128), .ZN(new_n405));
  XNOR2_X1  g219(.A(G143), .B(G146), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT0), .B(G128), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT64), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n404), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n187), .A2(KEYINPUT0), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT0), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G128), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT64), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n409), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n405), .B1(new_n408), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n402), .B1(new_n416), .B2(new_n204), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT1), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(G143), .B2(new_n304), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n409), .B1(new_n419), .B2(new_n187), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n406), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n204), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n408), .A2(new_n415), .ZN(new_n425));
  INV_X1    g239(.A(new_n405), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n427), .B2(G125), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n417), .B1(new_n428), .B2(new_n402), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n430));
  INV_X1    g244(.A(G224), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n430), .B1(new_n431), .B2(G953), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n228), .A2(KEYINPUT87), .A3(G224), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT86), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n429), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT3), .B1(new_n292), .B2(G107), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT3), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n337), .A3(G104), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n292), .A2(G107), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G101), .ZN(new_n443));
  INV_X1    g257(.A(G101), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n438), .A2(new_n440), .A3(new_n444), .A4(new_n441), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(KEYINPUT4), .A3(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(G116), .A2(G119), .ZN(new_n447));
  NOR2_X1   g261(.A1(G116), .A2(G119), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT2), .B(G113), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT4), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n442), .A2(new_n452), .A3(G101), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n446), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n292), .A2(G107), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n337), .A2(G104), .ZN(new_n456));
  OAI21_X1  g270(.A(G101), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n445), .A2(new_n457), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n449), .A2(new_n450), .ZN(new_n459));
  INV_X1    g273(.A(G113), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n334), .A2(KEYINPUT5), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n460), .B1(new_n461), .B2(new_n189), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT5), .B1(new_n447), .B2(new_n448), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n462), .A2(KEYINPUT84), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT84), .B1(new_n462), .B2(new_n463), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n458), .B(new_n459), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n454), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G110), .B(G122), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n454), .A2(new_n466), .A3(new_n468), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(KEYINPUT6), .A3(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n417), .B(new_n435), .C1(new_n428), .C2(new_n402), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n467), .A2(new_n474), .A3(new_n469), .ZN(new_n475));
  AND4_X1   g289(.A1(new_n437), .A2(new_n472), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n445), .A2(new_n457), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n459), .B(new_n477), .C1(new_n464), .C2(new_n465), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n468), .B(KEYINPUT8), .Z(new_n479));
  NAND2_X1  g293(.A1(new_n462), .A2(new_n463), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n459), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n481), .B2(new_n458), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n423), .B1(new_n416), .B2(new_n204), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n432), .A2(KEYINPUT7), .A3(new_n433), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n478), .A2(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n471), .B(new_n485), .C1(new_n429), .C2(new_n484), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n236), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n401), .B1(new_n476), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n437), .A2(new_n472), .A3(new_n473), .A4(new_n475), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n489), .A2(new_n236), .A3(new_n400), .A4(new_n486), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n399), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT83), .B(G469), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n420), .A2(new_n422), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT82), .B1(new_n458), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT1), .B1(new_n256), .B2(G146), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n187), .B1(new_n495), .B2(KEYINPUT80), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT80), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n419), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n406), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n421), .A2(new_n403), .A3(new_n404), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n458), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n495), .A2(G128), .B1(new_n403), .B2(new_n404), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(new_n500), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT82), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(new_n477), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n494), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT11), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n328), .B2(G137), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n231), .A2(KEYINPUT11), .A3(G134), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n328), .A2(G137), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n271), .A2(KEYINPUT65), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n512), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n514), .A2(new_n508), .A3(new_n509), .A4(new_n510), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n506), .A2(KEYINPUT12), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT12), .B1(new_n506), .B2(new_n516), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT10), .B1(new_n502), .B2(new_n500), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT81), .B1(new_n520), .B2(new_n477), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT81), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n458), .A2(new_n493), .A3(new_n522), .A4(KEYINPUT10), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT10), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n501), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n516), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n416), .A2(new_n446), .A3(new_n453), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n524), .A2(new_n526), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G110), .B(G140), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT79), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n228), .A2(G227), .ZN(new_n532));
  XOR2_X1   g346(.A(new_n531), .B(new_n532), .Z(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n519), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n516), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n533), .B1(new_n537), .B2(new_n529), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n236), .B(new_n492), .C1(new_n535), .C2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n529), .B1(new_n517), .B2(new_n518), .ZN(new_n540));
  INV_X1    g354(.A(new_n533), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n529), .A2(new_n533), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n537), .ZN(new_n544));
  AOI21_X1  g358(.A(G902), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G469), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n539), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(G221), .B1(new_n321), .B2(G902), .ZN(new_n548));
  XOR2_X1   g362(.A(new_n548), .B(KEYINPUT78), .Z(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n491), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n397), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT71), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n425), .A2(new_n516), .A3(new_n426), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT66), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n508), .A2(new_n509), .A3(new_n271), .A4(new_n510), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n328), .A2(G137), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n231), .A2(G134), .ZN(new_n558));
  OAI21_X1  g372(.A(G131), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n555), .B1(new_n503), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n493), .A2(KEYINPUT66), .A3(new_n556), .A4(new_n559), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n554), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT30), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT30), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n493), .A2(new_n556), .A3(new_n559), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n554), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n451), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT29), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n503), .A2(new_n560), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n571), .A2(KEYINPUT66), .B1(new_n416), .B2(new_n516), .ZN(new_n572));
  INV_X1    g386(.A(new_n451), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n572), .A2(KEYINPUT67), .A3(new_n573), .A4(new_n561), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n554), .A2(new_n561), .A3(new_n562), .A4(new_n573), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT67), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT26), .B(G101), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n254), .A2(G210), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n569), .A2(new_n570), .A3(new_n578), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n236), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT28), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n563), .A2(new_n451), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT69), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT69), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n563), .A2(new_n589), .A3(new_n451), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n586), .B1(new_n591), .B2(new_n578), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n554), .A2(new_n566), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n586), .B1(new_n593), .B2(new_n451), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT70), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT29), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n451), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n574), .A2(new_n577), .A3(KEYINPUT28), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n570), .ZN(new_n601));
  INV_X1    g415(.A(new_n583), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n585), .B1(new_n597), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(G472), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n553), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n563), .A2(new_n589), .A3(new_n451), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n589), .B1(new_n563), .B2(new_n451), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n574), .A2(new_n577), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT28), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n596), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n603), .B1(new_n614), .B2(KEYINPUT29), .ZN(new_n615));
  OAI211_X1 g429(.A(KEYINPUT71), .B(G472), .C1(new_n615), .C2(new_n585), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n607), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n602), .B1(new_n599), .B2(new_n600), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n554), .A2(new_n565), .A3(new_n566), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(KEYINPUT30), .B2(new_n563), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n578), .B(new_n602), .C1(new_n621), .C2(new_n573), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT31), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n568), .A2(new_n451), .B1(new_n577), .B2(new_n574), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT31), .B1(new_n625), .B2(new_n602), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n619), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(G472), .A2(G902), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(KEYINPUT32), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT72), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT32), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n622), .A2(new_n623), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n625), .A2(KEYINPUT31), .A3(new_n602), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n618), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n628), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n627), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n628), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n631), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n251), .B(new_n552), .C1(new_n617), .C2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G101), .ZN(G3));
  OAI21_X1  g455(.A(G472), .B1(new_n635), .B2(G902), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n540), .A2(new_n541), .B1(new_n543), .B2(new_n537), .ZN(new_n643));
  OAI21_X1  g457(.A(G469), .B1(new_n643), .B2(G902), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n549), .B1(new_n644), .B2(new_n539), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n627), .A2(new_n628), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n642), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n249), .A2(new_n244), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n247), .A3(new_n237), .ZN(new_n649));
  INV_X1    g463(.A(new_n243), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n491), .A2(new_n649), .A3(new_n650), .A4(new_n396), .ZN(new_n651));
  INV_X1    g465(.A(new_n301), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n311), .A2(new_n289), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n294), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n314), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n312), .A2(KEYINPUT91), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n297), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n318), .B1(new_n657), .B2(new_n302), .ZN(new_n658));
  INV_X1    g472(.A(new_n319), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n652), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n385), .B1(new_n384), .B2(new_n236), .ZN(new_n661));
  AOI211_X1 g475(.A(KEYINPUT98), .B(G902), .C1(new_n382), .C2(new_n383), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n375), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT33), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n384), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n375), .A2(G902), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n383), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n373), .A2(KEYINPUT99), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT99), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n359), .A2(new_n369), .B1(new_n348), .B2(new_n344), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(new_n322), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n669), .A2(KEYINPUT33), .A3(new_n672), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n665), .B(new_n666), .C1(new_n668), .C2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n663), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n660), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n647), .A2(new_n651), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT34), .B(G104), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT101), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n677), .B(new_n679), .ZN(G6));
  OAI21_X1  g494(.A(new_n376), .B1(new_n661), .B2(new_n662), .ZN(new_n681));
  INV_X1    g495(.A(new_n377), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n301), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(new_n658), .B2(new_n659), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n317), .A2(KEYINPUT102), .A3(new_n319), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n687), .A2(new_n647), .A3(new_n651), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT35), .B(G107), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G9));
  AND2_X1   g504(.A1(new_n225), .A2(new_n227), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n232), .A2(KEYINPUT36), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n238), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n649), .A2(new_n695), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n642), .A2(new_n646), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n552), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT37), .B(G110), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G12));
  INV_X1    g514(.A(G900), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n392), .B1(new_n393), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n683), .A2(new_n685), .A3(new_n686), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n645), .A2(new_n491), .A3(new_n696), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n706), .B1(new_n617), .B2(new_n639), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  NAND2_X1  g522(.A1(new_n488), .A2(new_n490), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(KEYINPUT103), .Z(new_n710));
  XOR2_X1   g524(.A(new_n710), .B(KEYINPUT38), .Z(new_n711));
  XOR2_X1   g525(.A(new_n702), .B(KEYINPUT39), .Z(new_n712));
  NAND2_X1  g526(.A1(new_n645), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n713), .B(KEYINPUT40), .Z(new_n714));
  INV_X1    g528(.A(new_n625), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n602), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n591), .A2(new_n578), .A3(new_n583), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n236), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G472), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n631), .A2(new_n637), .A3(new_n638), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n681), .A2(new_n682), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n660), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n722), .A2(new_n399), .A3(new_n696), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n711), .A2(new_n714), .A3(new_n720), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G143), .ZN(G45));
  NAND3_X1  g539(.A1(new_n660), .A2(new_n675), .A3(new_n703), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n705), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(new_n617), .B2(new_n639), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G146), .ZN(G48));
  AOI211_X1 g543(.A(new_n395), .B(new_n399), .C1(new_n488), .C2(new_n490), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n446), .A2(new_n453), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n731), .A2(new_n416), .B1(new_n525), .B2(new_n501), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n527), .B1(new_n732), .B2(new_n524), .ZN(new_n733));
  INV_X1    g547(.A(new_n529), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n541), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n529), .B(new_n533), .C1(new_n517), .C2(new_n518), .ZN(new_n736));
  AOI21_X1  g550(.A(G902), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n546), .ZN(new_n738));
  INV_X1    g552(.A(new_n492), .ZN(new_n739));
  AOI211_X1 g553(.A(G902), .B(new_n739), .C1(new_n735), .C2(new_n736), .ZN(new_n740));
  INV_X1    g554(.A(new_n548), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AND4_X1   g556(.A1(new_n660), .A2(new_n730), .A3(new_n742), .A4(new_n675), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n251), .B(new_n743), .C1(new_n617), .C2(new_n639), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT41), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G113), .ZN(G15));
  NAND2_X1  g560(.A1(new_n638), .A2(new_n637), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n633), .A2(new_n634), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n636), .B1(new_n748), .B2(new_n619), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT72), .B1(new_n749), .B2(KEYINPUT32), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n607), .A2(new_n616), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n730), .A2(new_n742), .A3(new_n251), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n687), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G116), .ZN(G18));
  NAND4_X1  g571(.A1(new_n320), .A2(new_n696), .A3(new_n388), .A4(new_n396), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n742), .A2(new_n491), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n753), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G119), .ZN(G21));
  NOR2_X1   g576(.A1(new_n624), .A2(new_n626), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n602), .B1(new_n612), .B2(new_n613), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n628), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n251), .A2(new_n642), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n396), .A3(new_n742), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(new_n320), .B2(new_n388), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n660), .A2(KEYINPUT104), .A3(new_n721), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n771), .A3(new_n491), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT105), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n770), .A2(new_n771), .A3(KEYINPUT105), .A4(new_n491), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n768), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n340), .ZN(G24));
  NAND3_X1  g591(.A1(new_n642), .A2(new_n765), .A3(new_n696), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n778), .A2(new_n759), .A3(new_n726), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n204), .ZN(G27));
  NAND3_X1  g594(.A1(new_n488), .A2(new_n398), .A3(new_n490), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT106), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n488), .A2(KEYINPUT106), .A3(new_n398), .A4(new_n490), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n251), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n547), .A2(new_n548), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n726), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n788), .B(new_n789), .C1(new_n617), .C2(new_n639), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT42), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT32), .B1(new_n627), .B2(new_n628), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n607), .A2(new_n616), .B1(KEYINPUT107), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n629), .A2(KEYINPUT107), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n637), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n786), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n785), .A2(new_n726), .A3(new_n791), .A4(new_n787), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n790), .A2(new_n791), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n271), .ZN(G33));
  INV_X1    g613(.A(new_n704), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n753), .A2(new_n800), .A3(new_n788), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  NAND2_X1  g616(.A1(new_n675), .A2(new_n320), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT43), .Z(new_n804));
  OR2_X1    g618(.A1(new_n804), .A2(KEYINPUT108), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n642), .A2(new_n646), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(KEYINPUT108), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n805), .A2(new_n806), .A3(new_n696), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n643), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT45), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n546), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n812), .B2(new_n811), .ZN(new_n814));
  NAND2_X1  g628(.A1(G469), .A2(G902), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT46), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n740), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(new_n817), .B2(new_n816), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n548), .A3(new_n712), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n810), .A2(new_n785), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n808), .A2(new_n809), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n822), .A2(KEYINPUT109), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(KEYINPUT109), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT110), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G137), .ZN(G39));
  NAND2_X1  g641(.A1(new_n819), .A2(new_n548), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT47), .ZN(new_n829));
  OR4_X1    g643(.A1(new_n753), .A2(new_n251), .A3(new_n726), .A4(new_n785), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(new_n202), .ZN(G42));
  NAND2_X1  g646(.A1(new_n298), .A2(new_n300), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n702), .B1(new_n833), .B2(G475), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n685), .A2(new_n388), .A3(new_n686), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT111), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n834), .A2(new_n681), .A3(new_n682), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT111), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n839), .A3(new_n685), .A4(new_n686), .ZN(new_n840));
  INV_X1    g654(.A(new_n785), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n836), .A2(new_n837), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n753), .A3(new_n645), .A4(new_n696), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n785), .B1(new_n835), .B2(KEYINPUT111), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n837), .B1(new_n844), .B2(new_n840), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OR4_X1    g660(.A1(new_n726), .A2(new_n778), .A3(new_n785), .A4(new_n787), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n801), .A2(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n846), .A2(new_n798), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  INV_X1    g664(.A(new_n779), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n707), .A2(new_n851), .A3(new_n728), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n787), .A2(new_n696), .A3(new_n702), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n720), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n774), .B2(new_n775), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n850), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n720), .A2(new_n853), .ZN(new_n857));
  INV_X1    g671(.A(new_n491), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n722), .B2(new_n769), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT105), .B1(new_n859), .B2(new_n771), .ZN(new_n860));
  INV_X1    g674(.A(new_n775), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n857), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n779), .B1(new_n753), .B2(new_n706), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n862), .A2(KEYINPUT52), .A3(new_n728), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n856), .A2(new_n864), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n755), .A2(new_n760), .B1(new_n617), .B2(new_n639), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(new_n744), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n647), .A2(new_n651), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n676), .B1(new_n660), .B2(new_n388), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n868), .A2(new_n869), .B1(new_n552), .B2(new_n697), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n640), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n742), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n766), .A2(new_n395), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n873), .B1(new_n860), .B2(new_n861), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n867), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n849), .A2(new_n865), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT113), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n866), .A2(new_n744), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n881), .B1(new_n882), .B2(new_n776), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n874), .A2(KEYINPUT113), .A3(new_n744), .A4(new_n866), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n871), .A2(KEYINPUT53), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n849), .A2(new_n865), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n879), .A2(new_n880), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n877), .B(new_n878), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n889), .B1(KEYINPUT54), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n804), .A2(new_n392), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n767), .ZN(new_n893));
  NOR4_X1   g707(.A1(new_n893), .A2(new_n398), .A3(new_n711), .A4(new_n872), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT50), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(KEYINPUT114), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n785), .A2(new_n872), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n778), .ZN(new_n899));
  INV_X1    g713(.A(new_n720), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n251), .A3(new_n392), .A4(new_n897), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n901), .A2(new_n660), .A3(new_n675), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g717(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n904));
  OAI211_X1 g718(.A(new_n896), .B(new_n903), .C1(new_n894), .C2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n539), .B1(new_n546), .B2(new_n737), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n907), .A2(new_n550), .ZN(new_n908));
  AOI211_X1 g722(.A(new_n785), .B(new_n893), .C1(new_n829), .C2(new_n908), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n906), .B1(new_n905), .B2(new_n909), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n892), .A2(new_n796), .A3(new_n897), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT48), .Z(new_n913));
  OAI221_X1 g727(.A(new_n389), .B1(new_n676), .B2(new_n901), .C1(new_n893), .C2(new_n759), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n891), .A2(new_n910), .A3(new_n911), .A4(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(G952), .B2(G953), .ZN(new_n917));
  INV_X1    g731(.A(new_n711), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n907), .B(KEYINPUT49), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n251), .A2(new_n398), .A3(new_n550), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n803), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n900), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n917), .A2(new_n922), .ZN(G75));
  NAND2_X1  g737(.A1(new_n437), .A2(new_n473), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n472), .A2(new_n475), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n489), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT115), .Z(new_n928));
  INV_X1    g742(.A(KEYINPUT55), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n879), .A2(new_n887), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n236), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(G210), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI211_X1 g749(.A(KEYINPUT55), .B(KEYINPUT56), .C1(new_n932), .C2(G210), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n928), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n228), .A2(G952), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT116), .Z(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n935), .A2(new_n936), .A3(new_n928), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(G51));
  NOR3_X1   g756(.A1(new_n931), .A2(new_n236), .A3(new_n814), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n875), .B1(new_n856), .B2(new_n864), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT53), .B1(new_n944), .B2(new_n849), .ZN(new_n945));
  AND4_X1   g759(.A1(new_n849), .A2(new_n865), .A3(new_n885), .A4(new_n886), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT54), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n947), .A2(KEYINPUT118), .A3(new_n888), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT118), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n930), .A2(new_n949), .A3(KEYINPUT54), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n815), .B(KEYINPUT117), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT57), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n948), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT119), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n948), .A2(KEYINPUT119), .A3(new_n950), .A4(new_n952), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n735), .A2(new_n736), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT120), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n943), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n957), .A2(KEYINPUT120), .A3(new_n958), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n938), .B1(new_n961), .B2(new_n962), .ZN(G54));
  NAND3_X1  g777(.A1(new_n932), .A2(KEYINPUT58), .A3(G475), .ZN(new_n964));
  INV_X1    g778(.A(new_n657), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n966), .A2(new_n967), .A3(new_n938), .ZN(G60));
  OAI21_X1  g782(.A(new_n665), .B1(new_n668), .B2(new_n673), .ZN(new_n969));
  NAND2_X1  g783(.A1(G478), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT59), .Z(new_n971));
  OAI21_X1  g785(.A(new_n969), .B1(new_n891), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT121), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n948), .A2(new_n950), .ZN(new_n974));
  OR3_X1    g788(.A1(new_n974), .A2(new_n969), .A3(new_n971), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n973), .A2(new_n939), .A3(new_n975), .ZN(G63));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT60), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n931), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n233), .A2(new_n234), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n939), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n693), .A2(new_n694), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT122), .Z(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT61), .ZN(G66));
  NOR3_X1   g799(.A1(new_n394), .A2(new_n431), .A3(new_n228), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n876), .B2(new_n228), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n925), .B1(G898), .B2(new_n228), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  INV_X1    g803(.A(new_n852), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n724), .A2(new_n990), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT62), .Z(new_n992));
  INV_X1    g806(.A(new_n831), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n785), .A2(new_n713), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n753), .A2(new_n251), .A3(new_n869), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n825), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(KEYINPUT124), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT124), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n825), .A2(new_n999), .A3(new_n996), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n994), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n621), .B(KEYINPUT123), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n303), .A2(new_n305), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n820), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1007), .B(new_n796), .C1(new_n860), .C2(new_n861), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n825), .A2(new_n993), .A3(new_n990), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n801), .ZN(new_n1010));
  NOR4_X1   g824(.A1(new_n1009), .A2(new_n798), .A3(new_n1010), .A4(new_n1004), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n228), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n701), .B1(new_n1005), .B2(G227), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1013), .B1(G227), .B2(new_n1005), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(G953), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1012), .A2(new_n1015), .ZN(G72));
  XNOR2_X1  g830(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n606), .A2(new_n236), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  OR3_X1    g833(.A1(new_n875), .A2(new_n798), .A3(new_n1010), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1019), .B1(new_n1009), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n715), .A2(new_n602), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n938), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1022), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1024), .A2(new_n716), .A3(new_n1019), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(KEYINPUT127), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n890), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1019), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1029), .B1(new_n1001), .B2(new_n876), .ZN(new_n1030));
  OR3_X1    g844(.A1(new_n1030), .A2(KEYINPUT126), .A3(new_n716), .ZN(new_n1031));
  OAI21_X1  g845(.A(KEYINPUT126), .B1(new_n1030), .B2(new_n716), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1028), .B1(new_n1031), .B2(new_n1032), .ZN(G57));
endmodule


