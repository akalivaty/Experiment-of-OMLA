//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(G29gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT86), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT86), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G29gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT14), .B1(new_n204), .B2(new_n203), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  NOR3_X1   g009(.A1(new_n210), .A2(G29gat), .A3(G36gat), .ZN(new_n211));
  NOR3_X1   g010(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(G43gat), .A2(G50gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT84), .ZN(new_n214));
  NAND2_X1  g013(.A1(G43gat), .A2(G50gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(G43gat), .A2(G50gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G43gat), .A2(G50gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT84), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n219), .A3(KEYINPUT15), .ZN(new_n220));
  OR3_X1    g019(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT15), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n212), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n203), .A3(KEYINPUT14), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n210), .B1(G29gat), .B2(G36gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT85), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT85), .B1(new_n223), .B2(new_n224), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n225), .A2(new_n226), .A3(new_n208), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT87), .B1(new_n227), .B2(new_n220), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT85), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(new_n211), .B2(new_n209), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT85), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n205), .A2(new_n207), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G36gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT87), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n216), .A2(new_n219), .A3(KEYINPUT15), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n222), .B1(new_n228), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G15gat), .B(G22gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT16), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(G1gat), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n241), .B(KEYINPUT88), .C1(G1gat), .C2(new_n239), .ZN(new_n242));
  INV_X1    g041(.A(G8gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n202), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n212), .A2(new_n220), .A3(new_n221), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n235), .B1(new_n234), .B2(new_n236), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n242), .B(G8gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(KEYINPUT89), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G229gat), .A2(G233gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT17), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(KEYINPUT17), .B(new_n246), .C1(new_n247), .C2(new_n248), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n244), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n252), .A2(new_n253), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT91), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n253), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(new_n260), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n252), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G113gat), .B(G141gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G169gat), .B(G197gat), .Z(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT12), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n245), .A2(new_n251), .B1(new_n244), .B2(new_n238), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n253), .B(KEYINPUT13), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n264), .B(new_n270), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n259), .B1(new_n258), .B2(new_n260), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n261), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n270), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n264), .B1(new_n271), .B2(new_n273), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n250), .B1(new_n249), .B2(new_n254), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n245), .A2(new_n251), .B1(new_n279), .B2(new_n256), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT18), .B1(new_n280), .B2(new_n253), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n277), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT90), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n258), .A2(new_n260), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n238), .A2(new_n244), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n252), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n272), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n288), .A3(new_n264), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(KEYINPUT90), .A3(new_n277), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n276), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT27), .B(G183gat), .ZN(new_n292));
  INV_X1    g091(.A(G190gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n294), .B(KEYINPUT28), .Z(new_n295));
  OAI21_X1  g094(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT67), .ZN(new_n297));
  NOR3_X1   g096(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n297), .A2(new_n299), .B1(G183gat), .B2(G190gat), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT24), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(G183gat), .A3(G190gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G183gat), .B(G190gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(new_n303), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n306), .A2(KEYINPUT64), .ZN(new_n307));
  INV_X1    g106(.A(G169gat), .ZN(new_n308));
  INV_X1    g107(.A(G176gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT23), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT23), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(G169gat), .B2(G176gat), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n310), .B(new_n312), .C1(new_n308), .C2(new_n309), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT65), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n313), .A2(KEYINPUT65), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n306), .A2(KEYINPUT64), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n307), .A2(new_n314), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT25), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n302), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n306), .A2(new_n313), .A3(new_n318), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n317), .A2(new_n302), .A3(new_n318), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n301), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n324));
  INV_X1    g123(.A(G120gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G113gat), .ZN(new_n326));
  INV_X1    g125(.A(G113gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G120gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n324), .B1(new_n331), .B2(KEYINPUT68), .ZN(new_n332));
  XOR2_X1   g131(.A(G127gat), .B(G134gat), .Z(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT69), .B1(new_n329), .B2(new_n330), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n335), .A2(new_n333), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n336), .B2(new_n332), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n323), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n337), .ZN(new_n339));
  AOI211_X1 g138(.A(new_n339), .B(new_n301), .C1(new_n321), .C2(new_n322), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT34), .ZN(new_n342));
  INV_X1    g141(.A(G227gat), .ZN(new_n343));
  INV_X1    g142(.A(G233gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n341), .A2(KEYINPUT72), .A3(new_n342), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n323), .A2(new_n337), .ZN(new_n348));
  INV_X1    g147(.A(new_n322), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n349), .A2(new_n319), .A3(new_n320), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n339), .B1(new_n350), .B2(new_n301), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT34), .B1(new_n352), .B2(new_n345), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n348), .A2(new_n351), .A3(new_n342), .A4(new_n346), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n347), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n352), .A2(new_n345), .ZN(new_n359));
  XOR2_X1   g158(.A(G71gat), .B(G99gat), .Z(new_n360));
  XNOR2_X1  g159(.A(G15gat), .B(G43gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n362), .A2(KEYINPUT70), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(KEYINPUT70), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(KEYINPUT33), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n359), .A2(KEYINPUT32), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n359), .A2(KEYINPUT32), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT33), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n359), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n369), .A3(new_n362), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n358), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n346), .B1(new_n348), .B2(new_n351), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT32), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n362), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n372), .A2(KEYINPUT33), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n366), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n357), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT36), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n371), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT71), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n357), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n376), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n370), .A2(new_n357), .A3(new_n380), .A4(new_n366), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT36), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G197gat), .B(G204gat), .ZN(new_n386));
  XOR2_X1   g185(.A(KEYINPUT73), .B(G218gat), .Z(new_n387));
  INV_X1    g186(.A(G211gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n386), .B1(new_n389), .B2(KEYINPUT22), .ZN(new_n390));
  XNOR2_X1  g189(.A(G211gat), .B(G218gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(KEYINPUT29), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n323), .A2(new_n395), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n350), .A2(new_n301), .A3(new_n394), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI22_X1  g197(.A1(new_n350), .A2(new_n301), .B1(KEYINPUT29), .B2(new_n394), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n323), .A2(new_n393), .ZN(new_n400));
  INV_X1    g199(.A(new_n392), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n398), .A2(new_n402), .A3(new_n406), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT30), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n398), .A2(new_n411), .A3(new_n402), .A4(new_n406), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G155gat), .A2(G162gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT74), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G155gat), .ZN(new_n417));
  INV_X1    g216(.A(G162gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(KEYINPUT74), .A2(G155gat), .A3(G162gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(G141gat), .B(G148gat), .Z(new_n422));
  INV_X1    g221(.A(KEYINPUT75), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n422), .A2(new_n423), .B1(KEYINPUT2), .B2(new_n414), .ZN(new_n424));
  XNOR2_X1  g223(.A(G141gat), .B(G148gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT75), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n421), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n419), .A2(KEYINPUT2), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n425), .B1(new_n428), .B2(new_n414), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT3), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n432), .B(new_n339), .C1(new_n433), .C2(new_n430), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n435));
  INV_X1    g234(.A(new_n430), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n435), .B1(new_n339), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n337), .A2(new_n430), .A3(KEYINPUT4), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n434), .A2(new_n437), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT77), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT5), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n337), .B(new_n430), .ZN(new_n443));
  INV_X1    g242(.A(new_n438), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n443), .A2(new_n444), .ZN(new_n447));
  OAI211_X1 g246(.A(KEYINPUT77), .B(new_n440), .C1(new_n447), .C2(new_n442), .ZN(new_n448));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT0), .ZN(new_n450));
  XOR2_X1   g249(.A(G57gat), .B(G85gat), .Z(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n446), .A2(new_n448), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n446), .B2(new_n448), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT78), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n455), .B(new_n454), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n457), .A2(new_n458), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n413), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n432), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n392), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n430), .A2(KEYINPUT29), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n401), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G228gat), .A2(G233gat), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n468), .B1(new_n436), .B2(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n430), .A2(new_n431), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n401), .B2(new_n466), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n473), .A2(new_n465), .B1(G228gat), .B2(G233gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G78gat), .B(G106gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT31), .B(G50gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n476), .B(new_n477), .Z(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n478), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n480), .B1(new_n471), .B2(new_n474), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT79), .ZN(new_n482));
  INV_X1    g281(.A(G22gat), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n481), .B2(new_n482), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n479), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n482), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(G22gat), .ZN(new_n488));
  INV_X1    g287(.A(new_n479), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n462), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n456), .B(new_n409), .C1(new_n459), .C2(new_n460), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT82), .B(KEYINPUT38), .Z(new_n495));
  INV_X1    g294(.A(KEYINPUT37), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n401), .B1(new_n399), .B2(new_n400), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT81), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(new_n402), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n402), .A2(new_n498), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n407), .B1(new_n403), .B2(KEYINPUT37), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n495), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n495), .B1(new_n403), .B2(KEYINPUT37), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n504), .B(new_n407), .C1(KEYINPUT37), .C2(new_n403), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n494), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n434), .A2(new_n437), .A3(new_n439), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n444), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n508), .A2(KEYINPUT39), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(new_n453), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT39), .B1(new_n443), .B2(new_n444), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT80), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(KEYINPUT80), .B(KEYINPUT39), .C1(new_n443), .C2(new_n444), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n508), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(KEYINPUT40), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n516), .A2(new_n454), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n510), .A2(new_n515), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT40), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n410), .A2(new_n517), .A3(new_n412), .A4(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n486), .A2(new_n491), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n385), .B(new_n493), .C1(new_n506), .C2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n492), .B1(new_n382), .B2(new_n383), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n457), .A2(new_n458), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n457), .A2(new_n458), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n526), .A2(new_n455), .A3(new_n527), .A4(new_n454), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n528), .A2(new_n456), .B1(new_n412), .B2(new_n410), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT35), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n522), .A2(new_n371), .A3(new_n377), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT35), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n413), .A2(new_n461), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n291), .B1(new_n524), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(KEYINPUT41), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(KEYINPUT93), .Z(new_n541));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  NAND2_X1  g345(.A1(G99gat), .A2(G106gat), .ZN(new_n547));
  INV_X1    g346(.A(G85gat), .ZN(new_n548));
  INV_X1    g347(.A(G92gat), .ZN(new_n549));
  AOI22_X1  g348(.A1(KEYINPUT8), .A2(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G99gat), .B(G106gat), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n546), .A3(new_n550), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n255), .A2(new_n256), .A3(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G190gat), .B(G218gat), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n556), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n249), .A2(new_n560), .B1(KEYINPUT41), .B2(new_n539), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n559), .B1(new_n557), .B2(new_n561), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n544), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n564), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(new_n543), .A3(new_n562), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G71gat), .A2(G78gat), .ZN(new_n569));
  OR2_X1    g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT9), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G64gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(G57gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(G57gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(KEYINPUT92), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT92), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n577), .A2(new_n573), .A3(G57gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n572), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(G57gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(G64gat), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT9), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n569), .A3(new_n570), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G127gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n244), .B1(new_n585), .B2(new_n584), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(new_n417), .ZN(new_n595));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n591), .A2(new_n592), .A3(new_n597), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n568), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n553), .A2(new_n555), .A3(new_n579), .A4(new_n583), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT94), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n604), .A3(KEYINPUT10), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n556), .A2(new_n584), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT10), .B1(new_n603), .B2(new_n604), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n602), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n603), .A2(new_n604), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n613), .A2(KEYINPUT95), .A3(new_n606), .A4(new_n605), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n609), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n606), .A2(new_n603), .ZN(new_n616));
  INV_X1    g415(.A(new_n610), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  NAND3_X1  g420(.A1(new_n615), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n613), .A2(new_n606), .A3(new_n605), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n618), .B1(new_n624), .B2(new_n617), .ZN(new_n625));
  INV_X1    g424(.A(new_n621), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n622), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n623), .B1(new_n622), .B2(new_n627), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n601), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n538), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n461), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G1gat), .ZN(G1324gat));
  INV_X1    g436(.A(new_n413), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n538), .A2(new_n638), .A3(new_n632), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n639), .A2(G8gat), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n640), .A2(KEYINPUT97), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT16), .B(G8gat), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OR3_X1    g442(.A1(new_n639), .A2(KEYINPUT42), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT42), .B1(new_n639), .B2(new_n643), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n640), .A2(KEYINPUT97), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n641), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT98), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT98), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n641), .A2(new_n646), .A3(new_n650), .A4(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(G1325gat));
  NAND2_X1  g451(.A1(new_n371), .A2(new_n377), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(G15gat), .B1(new_n634), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT99), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n379), .A2(new_n384), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n657), .A2(G15gat), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n656), .B1(new_n634), .B2(new_n658), .ZN(G1326gat));
  NOR2_X1   g458(.A1(new_n633), .A2(new_n522), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT43), .B(G22gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  NAND2_X1  g461(.A1(new_n599), .A2(new_n600), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT100), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n664), .A2(new_n291), .A3(new_n630), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n493), .B1(new_n506), .B2(new_n523), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n533), .B1(new_n525), .B2(new_n529), .ZN(new_n668));
  OAI22_X1  g467(.A1(new_n667), .A2(new_n657), .B1(new_n668), .B2(new_n535), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n669), .B2(new_n568), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n568), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n565), .A2(new_n567), .A3(KEYINPUT101), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(KEYINPUT44), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n524), .B2(new_n537), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n665), .B1(new_n670), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI211_X1 g479(.A(KEYINPUT102), .B(new_n665), .C1(new_n670), .C2(new_n677), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n635), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n232), .ZN(new_n683));
  INV_X1    g482(.A(new_n232), .ZN(new_n684));
  INV_X1    g483(.A(new_n568), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n663), .A2(new_n630), .A3(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n538), .A2(new_n635), .A3(new_n684), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT45), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT103), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n683), .A2(new_n691), .A3(new_n688), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(G1328gat));
  AND2_X1   g492(.A1(new_n538), .A2(new_n686), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n203), .A3(new_n638), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT46), .Z(new_n696));
  AND3_X1   g495(.A1(new_n680), .A2(new_n638), .A3(new_n681), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n203), .B2(new_n697), .ZN(G1329gat));
  OAI21_X1  g497(.A(G43gat), .B1(new_n678), .B2(new_n385), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n653), .A2(G43gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(KEYINPUT47), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n680), .A2(new_n657), .A3(new_n681), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n703), .A2(G43gat), .B1(new_n694), .B2(new_n700), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n704), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g504(.A(G50gat), .B1(new_n678), .B2(new_n522), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n522), .A2(G50gat), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n694), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(KEYINPUT48), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n680), .A2(new_n492), .A3(new_n681), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n710), .A2(G50gat), .B1(new_n694), .B2(new_n707), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT104), .B(KEYINPUT48), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n709), .B1(new_n711), .B2(new_n712), .ZN(G1331gat));
  NAND2_X1  g512(.A1(new_n291), .A2(new_n601), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n669), .A2(new_n630), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n635), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT105), .B(G57gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1332gat));
  AND2_X1   g518(.A1(new_n638), .A2(KEYINPUT106), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n638), .A2(KEYINPUT106), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT49), .B(G64gat), .Z(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n723), .B2(new_n725), .ZN(G1333gat));
  NAND2_X1  g525(.A1(new_n716), .A2(new_n657), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n653), .A2(G71gat), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n727), .A2(G71gat), .B1(new_n716), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g529(.A1(new_n716), .A2(new_n492), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g531(.A1(new_n670), .A2(new_n677), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n261), .A2(new_n274), .ZN(new_n734));
  INV_X1    g533(.A(new_n275), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n290), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT90), .B1(new_n289), .B2(new_n277), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n739), .A2(new_n663), .A3(new_n631), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n733), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n635), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G85gat), .ZN(new_n744));
  INV_X1    g543(.A(new_n663), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n669), .A2(new_n291), .A3(new_n745), .A4(new_n568), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n631), .B1(new_n748), .B2(KEYINPUT107), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(KEYINPUT107), .B2(new_n748), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n635), .A2(new_n548), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n744), .B1(new_n750), .B2(new_n751), .ZN(G1336gat));
  AOI21_X1  g551(.A(new_n549), .B1(new_n742), .B2(new_n638), .ZN(new_n753));
  INV_X1    g552(.A(new_n722), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n754), .A2(G92gat), .A3(new_n631), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n753), .B1(new_n748), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n549), .B1(new_n742), .B2(new_n722), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n748), .A2(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n757), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n756), .A2(new_n757), .B1(new_n758), .B2(new_n760), .ZN(G1337gat));
  NAND2_X1  g560(.A1(new_n742), .A2(new_n657), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G99gat), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n653), .A2(G99gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n750), .B2(new_n764), .ZN(G1338gat));
  NAND2_X1  g564(.A1(new_n742), .A2(new_n492), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G106gat), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n522), .A2(G106gat), .A3(new_n631), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT108), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n748), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT53), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT53), .B1(new_n748), .B2(new_n768), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n767), .A2(new_n773), .A3(KEYINPUT109), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT109), .B1(new_n767), .B2(new_n773), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n772), .B1(new_n774), .B2(new_n775), .ZN(G1339gat));
  NAND2_X1  g575(.A1(new_n715), .A2(new_n631), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n624), .B2(new_n617), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n615), .A2(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n607), .A2(new_n617), .A3(new_n608), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n621), .B1(new_n781), .B2(new_n778), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(KEYINPUT55), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n622), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT55), .B1(new_n780), .B2(new_n782), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT111), .B1(new_n287), .B2(new_n272), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n280), .B2(new_n253), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n252), .A2(new_n257), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(KEYINPUT110), .A3(new_n262), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n271), .A2(new_n792), .A3(new_n273), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n787), .A2(new_n789), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n269), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n786), .A2(new_n736), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n674), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n736), .A2(new_n630), .A3(new_n795), .ZN(new_n798));
  INV_X1    g597(.A(new_n786), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n291), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n797), .B1(new_n800), .B2(new_n674), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n777), .B1(new_n801), .B2(new_n664), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n802), .A2(new_n522), .A3(new_n654), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n635), .B1(new_n720), .B2(new_n721), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n327), .B1(new_n806), .B2(new_n739), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n807), .B(KEYINPUT112), .Z(new_n808));
  AND2_X1   g607(.A1(new_n802), .A2(new_n635), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n809), .A2(new_n525), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n754), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n327), .A3(new_n739), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n808), .A2(new_n813), .ZN(G1340gat));
  INV_X1    g613(.A(new_n806), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n815), .A2(new_n325), .A3(new_n631), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n630), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n325), .B2(new_n817), .ZN(G1341gat));
  NOR3_X1   g617(.A1(new_n811), .A2(G127gat), .A3(new_n745), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n806), .A2(new_n664), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(G127gat), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT113), .ZN(G1342gat));
  INV_X1    g621(.A(G134gat), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n638), .A2(new_n685), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n810), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n826));
  OAI21_X1  g625(.A(G134gat), .B1(new_n815), .B2(new_n685), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(G1343gat));
  INV_X1    g628(.A(G141gat), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n809), .B(KEYINPUT115), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n657), .A2(new_n522), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT116), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n754), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n830), .B1(new_n834), .B2(new_n291), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n804), .A2(new_n657), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT57), .B1(new_n802), .B2(new_n492), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n492), .A2(KEYINPUT57), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n780), .A2(new_n782), .ZN(new_n839));
  XOR2_X1   g638(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n840));
  OAI211_X1 g639(.A(new_n622), .B(new_n783), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n739), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n568), .B1(new_n843), .B2(new_n798), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n745), .B1(new_n844), .B2(new_n797), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n838), .B1(new_n845), .B2(new_n777), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n836), .B1(new_n837), .B2(new_n846), .ZN(new_n847));
  OR3_X1    g646(.A1(new_n847), .A2(new_n830), .A3(new_n291), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n835), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n849), .B(new_n850), .ZN(G1344gat));
  OAI211_X1 g650(.A(new_n630), .B(new_n836), .C1(new_n837), .C2(new_n846), .ZN(new_n852));
  INV_X1    g651(.A(G148gat), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(KEYINPUT59), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n852), .A2(KEYINPUT117), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT117), .B1(new_n852), .B2(new_n854), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n802), .A2(KEYINPUT57), .A3(new_n492), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n714), .B2(new_n630), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n291), .A2(KEYINPUT119), .A3(new_n631), .A4(new_n601), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND4_X1   g661(.A1(new_n736), .A2(new_n786), .A3(new_n568), .A4(new_n795), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n798), .B1(new_n291), .B2(new_n841), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(new_n685), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n745), .B1(new_n865), .B2(KEYINPUT120), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867));
  AOI211_X1 g666(.A(new_n867), .B(new_n863), .C1(new_n864), .C2(new_n685), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n862), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n871), .B(new_n862), .C1(new_n866), .C2(new_n868), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n492), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n858), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n836), .A2(new_n630), .ZN(new_n876));
  OAI21_X1  g675(.A(G148gat), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n857), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n834), .A2(G148gat), .A3(new_n631), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT122), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n881), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n522), .B1(new_n869), .B2(KEYINPUT121), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n885), .B2(new_n872), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n630), .B(new_n836), .C1(new_n886), .C2(new_n858), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n878), .B1(new_n887), .B2(G148gat), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n883), .B(new_n884), .C1(new_n888), .C2(new_n857), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n882), .A2(new_n889), .ZN(G1345gat));
  OR3_X1    g689(.A1(new_n834), .A2(G155gat), .A3(new_n745), .ZN(new_n891));
  INV_X1    g690(.A(new_n664), .ZN(new_n892));
  OAI21_X1  g691(.A(G155gat), .B1(new_n847), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n891), .A2(KEYINPUT123), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n847), .B2(new_n674), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n831), .A2(new_n833), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n824), .A2(new_n418), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(G1347gat));
  NOR2_X1   g701(.A1(new_n635), .A2(new_n413), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n803), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(new_n308), .A3(new_n291), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n802), .A2(new_n722), .A3(new_n461), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n525), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT124), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n739), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n905), .B1(new_n909), .B2(new_n308), .ZN(G1348gat));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n309), .A3(new_n630), .ZN(new_n911));
  OAI21_X1  g710(.A(G176gat), .B1(new_n904), .B2(new_n631), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1349gat));
  OAI21_X1  g712(.A(G183gat), .B1(new_n904), .B2(new_n892), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n663), .A2(new_n292), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n914), .B(KEYINPUT125), .C1(new_n907), .C2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g716(.A(G190gat), .B1(new_n904), .B2(new_n685), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT61), .ZN(new_n919));
  INV_X1    g718(.A(new_n674), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n908), .A2(new_n293), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1351gat));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n832), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(G197gat), .B1(new_n924), .B2(new_n739), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n385), .A2(new_n903), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n875), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n739), .A2(G197gat), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(G1352gat));
  INV_X1    g728(.A(new_n927), .ZN(new_n930));
  OAI21_X1  g729(.A(G204gat), .B1(new_n930), .B2(new_n631), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932));
  AOI21_X1  g731(.A(G204gat), .B1(new_n932), .B2(KEYINPUT62), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n924), .A2(new_n630), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n934), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n931), .A2(new_n936), .ZN(G1353gat));
  NAND2_X1  g736(.A1(new_n927), .A2(new_n663), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G211gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT63), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n941), .A3(G211gat), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n923), .A2(G211gat), .A3(new_n745), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT127), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n940), .A2(new_n942), .A3(new_n944), .ZN(G1354gat));
  AOI21_X1  g744(.A(G218gat), .B1(new_n924), .B2(new_n920), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n685), .A2(new_n387), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n927), .B2(new_n947), .ZN(G1355gat));
endmodule


