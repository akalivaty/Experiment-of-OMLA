//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT12), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT79), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(KEYINPUT79), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G104), .B(G107), .ZN(new_n193));
  INV_X1    g007(.A(G101), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT77), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n196), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(G107), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n197), .A2(new_n200), .A3(new_n194), .A4(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n199), .A2(G104), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n196), .A2(G107), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n203), .B(G101), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n195), .A2(new_n202), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n210), .A2(G143), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G128), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n212), .A2(G128), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n214), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n207), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n214), .A2(KEYINPUT78), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n210), .A2(new_n219), .B1(new_n215), .B2(new_n217), .ZN(new_n225));
  XNOR2_X1  g039(.A(G143), .B(G146), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT78), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n209), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n224), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n223), .B1(new_n207), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n231));
  INV_X1    g045(.A(G134), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G137), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G137), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT11), .A3(G134), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(G137), .ZN(new_n238));
  OAI211_X1 g052(.A(KEYINPUT64), .B(new_n231), .C1(new_n232), .C2(G137), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n235), .A2(new_n237), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G131), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n237), .A2(new_n238), .ZN(new_n242));
  INV_X1    g056(.A(G131), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n242), .A2(new_n243), .A3(new_n235), .A4(new_n239), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  AOI211_X1 g059(.A(new_n190), .B(new_n192), .C1(new_n230), .C2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n230), .A2(KEYINPUT79), .A3(new_n189), .A4(new_n245), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT10), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n249), .B1(new_n229), .B2(new_n207), .ZN(new_n250));
  INV_X1    g064(.A(new_n239), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n236), .A2(G134), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT64), .B1(new_n252), .B2(new_n231), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n243), .B1(new_n254), .B2(new_n242), .ZN(new_n255));
  INV_X1    g069(.A(new_n244), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n197), .A2(new_n200), .A3(new_n201), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G101), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n226), .A2(new_n261), .ZN(new_n262));
  OR2_X1    g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n263), .A2(new_n261), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n262), .B1(new_n264), .B2(new_n226), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n258), .A2(new_n266), .A3(G101), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n260), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n195), .A2(new_n202), .A3(new_n206), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n249), .B1(new_n225), .B2(new_n214), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n250), .A2(new_n257), .A3(new_n268), .A4(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G110), .B(G140), .ZN(new_n273));
  INV_X1    g087(.A(G227), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G953), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n273), .B(new_n275), .Z(new_n276));
  NAND2_X1  g090(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n246), .A2(new_n248), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n250), .A2(new_n268), .A3(new_n271), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n245), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n276), .B1(new_n280), .B2(new_n272), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n187), .B(new_n188), .C1(new_n278), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n230), .A2(new_n245), .ZN(new_n283));
  INV_X1    g097(.A(new_n190), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n191), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(new_n272), .A3(new_n247), .ZN(new_n286));
  INV_X1    g100(.A(new_n276), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n277), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n280), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(G469), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(G469), .A2(G902), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n282), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT9), .B(G234), .Z(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G221), .B1(new_n295), .B2(G902), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G210), .B1(G237), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n265), .A2(G125), .ZN(new_n300));
  INV_X1    g114(.A(G125), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n221), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G224), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(G953), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n305), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n300), .A2(new_n307), .A3(new_n302), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n306), .B(new_n308), .C1(KEYINPUT7), .C2(new_n305), .ZN(new_n309));
  INV_X1    g123(.A(G119), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G116), .ZN(new_n311));
  INV_X1    g125(.A(G116), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G119), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT2), .B(G113), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT5), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n310), .A3(G116), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n318), .B(G113), .C1(new_n314), .C2(new_n317), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n269), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT81), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n316), .A2(new_n319), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(new_n207), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(G110), .B(G122), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT8), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n320), .A2(new_n269), .A3(new_n322), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n314), .A2(new_n315), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n316), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n260), .A2(new_n331), .A3(new_n267), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n321), .A2(new_n332), .A3(new_n326), .ZN(new_n333));
  OR3_X1    g147(.A1(new_n303), .A2(KEYINPUT7), .A3(new_n305), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n309), .A2(new_n329), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n188), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n306), .A2(new_n308), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n321), .A2(new_n332), .A3(new_n326), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n326), .B(KEYINPUT80), .Z(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n340), .B1(new_n321), .B2(new_n332), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT6), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n321), .A2(new_n332), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n339), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n337), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n299), .B1(new_n336), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n337), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n345), .B1(new_n344), .B2(new_n333), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n341), .A2(KEYINPUT6), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n352), .A2(new_n188), .A3(new_n298), .A4(new_n335), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n353), .A3(KEYINPUT82), .ZN(new_n354));
  OAI21_X1  g168(.A(G214), .B1(G237), .B2(G902), .ZN(new_n355));
  INV_X1    g169(.A(new_n336), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n356), .A2(new_n352), .A3(new_n357), .A4(new_n298), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n354), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n312), .A2(G122), .ZN(new_n360));
  INV_X1    g174(.A(G122), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G116), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n362), .A3(new_n199), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G128), .B(G143), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(G134), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT14), .B1(new_n361), .B2(G116), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT85), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT85), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n360), .A2(new_n369), .A3(KEYINPUT14), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n362), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n360), .A2(KEYINPUT14), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT86), .A4(new_n362), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n364), .B(new_n366), .C1(new_n376), .C2(G107), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n360), .A2(new_n362), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G107), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n379), .A2(new_n363), .B1(new_n232), .B2(new_n365), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n365), .A2(KEYINPUT13), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n212), .A2(G128), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n381), .B(G134), .C1(KEYINPUT13), .C2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n380), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n380), .B2(new_n383), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G217), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n295), .A2(new_n389), .A3(G953), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n377), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n376), .A2(G107), .ZN(new_n393));
  INV_X1    g207(.A(new_n366), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n363), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n387), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n385), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n390), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n188), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G478), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT15), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n391), .B1(new_n377), .B2(new_n388), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n395), .A2(new_n397), .A3(new_n390), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT87), .A3(new_n188), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n401), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n399), .A2(new_n403), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n411));
  INV_X1    g225(.A(G953), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G952), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(G234), .B2(G237), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  XOR2_X1   g229(.A(KEYINPUT21), .B(G898), .Z(new_n416));
  NAND2_X1  g230(.A1(G234), .A2(G237), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(G902), .A3(G953), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n415), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G475), .ZN(new_n420));
  XNOR2_X1  g234(.A(G113), .B(G122), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(G104), .ZN(new_n424));
  NOR2_X1   g238(.A1(G237), .A2(G953), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(G143), .A3(G214), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(G143), .B1(new_n425), .B2(G214), .ZN(new_n428));
  OAI21_X1  g242(.A(G131), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n428), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n243), .A3(new_n426), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT17), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n301), .A2(KEYINPUT16), .A3(G140), .ZN(new_n434));
  XNOR2_X1  g248(.A(G125), .B(G140), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(KEYINPUT16), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n436), .A2(G146), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(G146), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n430), .A2(new_n426), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(KEYINPUT17), .A3(G131), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n433), .A2(new_n437), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n435), .B(new_n210), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT18), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(new_n243), .ZN(new_n444));
  OAI221_X1 g258(.A(new_n442), .B1(new_n439), .B2(new_n444), .C1(new_n429), .C2(new_n443), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n424), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n435), .B(KEYINPUT19), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n210), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT75), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n438), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n429), .A2(new_n431), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n436), .A2(KEYINPUT75), .A3(G146), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n449), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n424), .B1(new_n445), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n420), .B(new_n188), .C1(new_n447), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT20), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n454), .A2(new_n445), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n446), .B1(new_n458), .B2(new_n424), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n420), .A4(new_n188), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n424), .B1(new_n445), .B2(new_n441), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n188), .B1(new_n447), .B2(new_n462), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n457), .A2(new_n461), .B1(G475), .B2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n410), .A2(new_n411), .A3(new_n419), .A4(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n408), .A2(new_n464), .A3(new_n419), .A4(new_n409), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT88), .ZN(new_n467));
  AOI211_X1 g281(.A(new_n297), .B(new_n359), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n211), .A2(new_n213), .B1(new_n263), .B2(new_n261), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n211), .A2(new_n213), .A3(new_n261), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n241), .B2(new_n244), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT65), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n252), .A2(new_n238), .A3(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(G131), .C1(new_n473), .C2(new_n252), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n244), .A2(new_n221), .A3(new_n475), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n472), .A2(new_n476), .A3(new_n331), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n265), .B1(new_n255), .B2(new_n256), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT30), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n244), .A2(new_n221), .A3(new_n475), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT30), .B1(new_n472), .B2(new_n476), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n477), .B1(new_n483), .B2(new_n331), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT26), .B(G101), .Z(new_n486));
  NAND2_X1  g300(.A1(new_n425), .A2(G210), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT29), .ZN(new_n492));
  INV_X1    g306(.A(new_n331), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n478), .B2(new_n480), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT28), .B1(new_n494), .B2(new_n477), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT68), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n477), .B2(KEYINPUT28), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n478), .A2(new_n493), .A3(new_n480), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT28), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(KEYINPUT68), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n491), .B(new_n492), .C1(new_n490), .C2(new_n501), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n503), .A2(new_n497), .A3(new_n500), .A4(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n490), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT29), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n502), .B(new_n188), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G472), .ZN(new_n509));
  NOR2_X1   g323(.A1(G472), .A2(G902), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT70), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n479), .B1(new_n478), .B2(new_n480), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n472), .A2(new_n476), .A3(KEYINPUT30), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n331), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n498), .A3(new_n506), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(KEYINPUT31), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT67), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n484), .A2(KEYINPUT67), .A3(new_n506), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n516), .B1(new_n520), .B2(KEYINPUT31), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT69), .B1(new_n501), .B2(new_n490), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n501), .A2(KEYINPUT69), .A3(new_n490), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI211_X1 g339(.A(KEYINPUT32), .B(new_n511), .C1(new_n521), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT32), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT67), .B1(new_n484), .B2(new_n506), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n493), .B1(new_n481), .B2(new_n482), .ZN(new_n529));
  NOR4_X1   g343(.A1(new_n529), .A2(new_n517), .A3(new_n477), .A4(new_n490), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT31), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n516), .ZN(new_n532));
  INV_X1    g346(.A(new_n524), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n531), .B(new_n532), .C1(new_n522), .C2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n511), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n527), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n509), .B1(new_n526), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT76), .ZN(new_n538));
  XOR2_X1   g352(.A(G119), .B(G128), .Z(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT24), .B(G110), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT23), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(new_n310), .B2(G128), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT73), .B1(new_n310), .B2(G128), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n541), .B1(new_n545), .B2(G110), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n546), .A2(KEYINPUT74), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n451), .A2(new_n453), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n435), .A2(new_n210), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(KEYINPUT74), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n437), .A2(new_n438), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n545), .A2(G110), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n552), .B(new_n553), .C1(new_n539), .C2(new_n540), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n412), .A2(G221), .A3(G234), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT22), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(G137), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n551), .A2(new_n554), .A3(new_n558), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n538), .B(KEYINPUT25), .C1(new_n562), .C2(G902), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n389), .B1(G234), .B2(new_n188), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n565), .A2(KEYINPUT72), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(KEYINPUT72), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT76), .B(KEYINPUT25), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n560), .A2(new_n188), .A3(new_n561), .A4(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n563), .A2(new_n566), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n564), .A2(G902), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n560), .A2(new_n561), .A3(new_n571), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n468), .A2(new_n537), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G101), .ZN(G3));
  AOI21_X1  g389(.A(new_n511), .B1(new_n521), .B2(new_n525), .ZN(new_n576));
  INV_X1    g390(.A(G472), .ZN(new_n577));
  AOI21_X1  g391(.A(G902), .B1(new_n521), .B2(new_n525), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n577), .B1(new_n578), .B2(KEYINPUT89), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n534), .A2(new_n188), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT89), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n576), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n464), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n406), .A2(KEYINPUT33), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n406), .A2(KEYINPUT33), .ZN(new_n586));
  AOI211_X1 g400(.A(new_n402), .B(G902), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n401), .A2(new_n402), .A3(new_n407), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n355), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n348), .B2(new_n353), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n419), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n297), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n573), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n583), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G104), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n596), .B(new_n598), .ZN(G6));
  INV_X1    g413(.A(new_n457), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n461), .B1(new_n600), .B2(KEYINPUT91), .ZN(new_n601));
  OR3_X1    g415(.A1(new_n456), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n601), .A2(new_n602), .B1(G475), .B2(new_n463), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n408), .A2(new_n409), .ZN(new_n604));
  AND4_X1   g418(.A1(new_n419), .A2(new_n603), .A3(new_n604), .A4(new_n591), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n583), .A2(new_n595), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT35), .B(G107), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  NOR2_X1   g422(.A1(new_n559), .A2(KEYINPUT36), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT92), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(new_n555), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n571), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n570), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT93), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT93), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n570), .A2(new_n615), .A3(new_n612), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n468), .A2(new_n583), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT37), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G110), .ZN(G12));
  OR3_X1    g434(.A1(new_n418), .A2(KEYINPUT94), .A3(G900), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT94), .B1(new_n418), .B2(G900), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n415), .A3(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n603), .A2(new_n604), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n591), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n297), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n537), .A2(new_n617), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G128), .ZN(G30));
  NAND2_X1  g442(.A1(new_n354), .A2(new_n358), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT95), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT38), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n355), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n623), .B(KEYINPUT39), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n594), .A2(new_n633), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n464), .B(new_n410), .C1(new_n634), .C2(KEYINPUT40), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(KEYINPUT40), .B2(new_n634), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n490), .B1(new_n494), .B2(new_n477), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n637), .A2(KEYINPUT96), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n577), .B1(new_n637), .B2(KEYINPUT96), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n638), .B(new_n639), .C1(new_n528), .C2(new_n530), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n641));
  NAND2_X1  g455(.A1(G472), .A2(G902), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n641), .B1(new_n640), .B2(new_n642), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n526), .B2(new_n536), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NOR4_X1   g461(.A1(new_n632), .A2(new_n636), .A3(new_n613), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n212), .ZN(G45));
  INV_X1    g463(.A(new_n623), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n589), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n537), .A2(new_n617), .A3(new_n626), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT98), .B(G146), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G48));
  AND2_X1   g468(.A1(new_n537), .A2(new_n573), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n278), .A2(new_n281), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n188), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G469), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n296), .A3(new_n282), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n655), .A2(new_n593), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT41), .B(G113), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT99), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(G15));
  NAND4_X1  g478(.A1(new_n537), .A2(new_n573), .A3(new_n605), .A4(new_n660), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G116), .ZN(G18));
  NAND2_X1  g480(.A1(new_n465), .A2(new_n467), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n659), .A2(new_n625), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n537), .A2(new_n617), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT100), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G119), .ZN(G21));
  NAND2_X1  g485(.A1(new_n505), .A2(new_n490), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n511), .B1(new_n521), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n580), .B2(G472), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n674), .A2(new_n573), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n604), .A2(new_n584), .A3(new_n591), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n604), .A2(new_n591), .A3(KEYINPUT101), .A4(new_n584), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n675), .A2(new_n419), .A3(new_n660), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G122), .ZN(G24));
  NAND4_X1  g496(.A1(new_n674), .A2(new_n668), .A3(new_n651), .A4(new_n613), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G125), .ZN(G27));
  NAND2_X1  g498(.A1(new_n629), .A2(new_n355), .ZN(new_n685));
  INV_X1    g499(.A(new_n296), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n292), .B(KEYINPUT102), .Z(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n286), .A2(new_n287), .B1(new_n280), .B2(new_n289), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n688), .B1(new_n689), .B2(G469), .ZN(new_n690));
  AOI211_X1 g504(.A(KEYINPUT103), .B(new_n686), .C1(new_n690), .C2(new_n282), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n282), .A2(new_n291), .A3(new_n687), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n692), .B1(new_n693), .B2(new_n296), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n685), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  AND4_X1   g509(.A1(new_n537), .A2(new_n573), .A3(new_n651), .A4(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT105), .B1(new_n696), .B2(KEYINPUT42), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n537), .A2(new_n573), .A3(new_n651), .A4(new_n695), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n698), .A2(new_n702), .A3(new_n700), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n702), .B1(new_n698), .B2(new_n700), .ZN(new_n704));
  OAI22_X1  g518(.A1(new_n697), .A2(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G131), .ZN(G33));
  NAND4_X1  g520(.A1(new_n537), .A2(new_n573), .A3(new_n624), .A4(new_n695), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G134), .ZN(G36));
  NAND2_X1  g522(.A1(new_n689), .A2(KEYINPUT45), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(KEYINPUT106), .Z(new_n710));
  OAI211_X1 g524(.A(new_n710), .B(G469), .C1(KEYINPUT45), .C2(new_n689), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n687), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n711), .A2(KEYINPUT46), .A3(new_n687), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n282), .A3(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n716), .A2(new_n296), .ZN(new_n717));
  INV_X1    g531(.A(new_n613), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n583), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n719), .B(KEYINPUT108), .Z(new_n720));
  OR2_X1    g534(.A1(new_n587), .A2(new_n588), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n464), .B(KEYINPUT107), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n723), .A2(new_n464), .B1(new_n725), .B2(KEYINPUT43), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n633), .B(new_n717), .C1(new_n728), .C2(KEYINPUT44), .ZN(new_n729));
  INV_X1    g543(.A(new_n685), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n730), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT109), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G137), .ZN(G39));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n716), .A2(new_n296), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT110), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n737), .A2(KEYINPUT110), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n736), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n737), .A2(KEYINPUT110), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(KEYINPUT47), .A3(new_n738), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n537), .ZN(new_n745));
  NOR4_X1   g559(.A1(new_n573), .A2(new_n589), .A3(new_n685), .A4(new_n650), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT111), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G140), .ZN(G42));
  NOR4_X1   g563(.A1(new_n631), .A2(new_n686), .A3(new_n590), .A4(new_n725), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n658), .A2(new_n282), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n751), .B(KEYINPUT49), .Z(new_n752));
  NAND4_X1  g566(.A1(new_n750), .A2(new_n573), .A3(new_n647), .A4(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n726), .A2(new_n414), .A3(new_n675), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n751), .A2(new_n296), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n730), .B(new_n754), .C1(new_n744), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n659), .A2(new_n685), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n647), .A2(new_n573), .A3(new_n414), .A4(new_n757), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n758), .A2(new_n584), .A3(new_n721), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n660), .A2(new_n590), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n631), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n762), .B(new_n754), .C1(new_n760), .C2(new_n761), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT50), .Z(new_n764));
  NAND3_X1  g578(.A1(new_n726), .A2(new_n414), .A3(new_n757), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT116), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n674), .A2(new_n613), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n756), .A2(new_n759), .A3(new_n764), .A4(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n413), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n354), .A2(new_n419), .A3(new_n355), .A4(new_n358), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n604), .A2(new_n464), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OR3_X1    g590(.A1(new_n774), .A2(new_n775), .A3(new_n773), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n583), .A2(new_n595), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n589), .A2(new_n774), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n583), .A2(new_n595), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n778), .A2(new_n618), .A3(new_n574), .A4(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n767), .A2(new_n651), .A3(new_n695), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n707), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n730), .A2(new_n603), .A3(new_n410), .A4(new_n623), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n537), .A2(new_n617), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n786), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n787), .A2(new_n788), .A3(new_n594), .A4(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n627), .A2(new_n683), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n686), .B(new_n650), .C1(new_n690), .C2(new_n282), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n646), .A2(new_n680), .A3(new_n718), .A4(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n791), .A2(new_n792), .A3(new_n652), .A4(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n627), .A2(new_n652), .A3(new_n794), .A4(new_n683), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT52), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n784), .A2(new_n790), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n661), .A2(new_n665), .A3(new_n669), .A4(new_n681), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n705), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n772), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n790), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n802), .A2(new_n781), .A3(new_n783), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n796), .B(new_n792), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n661), .A2(new_n665), .A3(new_n669), .A4(new_n681), .ZN(new_n805));
  OAI21_X1  g619(.A(KEYINPUT104), .B1(new_n696), .B2(KEYINPUT42), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n698), .A2(new_n702), .A3(new_n700), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n696), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n805), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n803), .B(new_n804), .C1(new_n812), .C2(KEYINPUT114), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n705), .A2(KEYINPUT114), .A3(new_n799), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT53), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n801), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n812), .A2(new_n803), .A3(new_n804), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT53), .ZN(new_n818));
  MUX2_X1   g632(.A(new_n816), .B(new_n818), .S(KEYINPUT54), .Z(new_n819));
  OAI211_X1 g633(.A(new_n771), .B(new_n819), .C1(new_n770), .C2(new_n769), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n754), .A2(new_n668), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n758), .A2(new_n589), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n766), .A2(new_n655), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT48), .Z(new_n824));
  NOR4_X1   g638(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(G952), .A2(G953), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n753), .B1(new_n825), .B2(new_n826), .ZN(G75));
  AOI21_X1  g641(.A(KEYINPUT114), .B1(new_n705), .B2(new_n799), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n798), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n772), .B1(new_n812), .B2(KEYINPUT114), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n829), .A2(new_n830), .B1(new_n772), .B2(new_n817), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n188), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT56), .B1(new_n832), .B2(G210), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n350), .A2(new_n351), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(new_n349), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT55), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n833), .B(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n412), .A2(G952), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(G51));
  XNOR2_X1  g653(.A(new_n816), .B(KEYINPUT54), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n687), .B(KEYINPUT57), .Z(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n656), .ZN(new_n843));
  OR3_X1    g657(.A1(new_n831), .A2(new_n188), .A3(new_n711), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n838), .B1(new_n843), .B2(new_n844), .ZN(G54));
  NAND3_X1  g659(.A1(new_n832), .A2(KEYINPUT58), .A3(G475), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(new_n459), .Z(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n838), .ZN(G60));
  NAND2_X1  g662(.A1(new_n585), .A2(new_n586), .ZN(new_n849));
  NAND2_X1  g663(.A1(G478), .A2(G902), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT59), .Z(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n840), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n586), .B(new_n585), .C1(new_n819), .C2(new_n851), .ZN(new_n856));
  INV_X1    g670(.A(new_n838), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n840), .A2(KEYINPUT117), .A3(new_n849), .A4(new_n852), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n855), .A2(new_n856), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n859), .B(new_n860), .ZN(G63));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n862));
  XNOR2_X1  g676(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n864));
  NAND2_X1  g678(.A1(G217), .A2(G902), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT60), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n864), .B1(new_n831), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n866), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n816), .A2(KEYINPUT120), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n562), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n611), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n867), .B2(new_n869), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n800), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n778), .A2(new_n618), .A3(new_n574), .ZN(new_n877));
  INV_X1    g691(.A(new_n783), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n790), .A4(new_n780), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n795), .A2(new_n797), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n876), .A2(new_n881), .A3(KEYINPUT53), .A4(new_n814), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n864), .B(new_n866), .C1(new_n882), .C2(new_n801), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT120), .B1(new_n816), .B2(new_n868), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n873), .B(new_n611), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n857), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n862), .B(new_n863), .C1(new_n874), .C2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n611), .B1(new_n883), .B2(new_n884), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT121), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(new_n857), .A3(new_n885), .A4(new_n870), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n862), .B1(new_n891), .B2(new_n863), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n870), .A2(KEYINPUT123), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n867), .A2(new_n894), .A3(new_n562), .A4(new_n869), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n872), .A2(new_n838), .ZN(new_n897));
  AND4_X1   g711(.A1(KEYINPUT124), .A2(new_n896), .A3(KEYINPUT61), .A4(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n893), .B2(new_n895), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT124), .B1(new_n900), .B2(new_n897), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n888), .A2(new_n892), .B1(new_n898), .B2(new_n901), .ZN(G66));
  INV_X1    g716(.A(new_n416), .ZN(new_n903));
  OAI21_X1  g717(.A(G953), .B1(new_n903), .B2(new_n304), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n805), .A2(new_n781), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n904), .B1(new_n905), .B2(G953), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n834), .B1(G898), .B2(new_n412), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n906), .B(new_n907), .ZN(G69));
  INV_X1    g722(.A(G900), .ZN(new_n909));
  OAI21_X1  g723(.A(G953), .B1(new_n274), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT126), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n589), .A2(new_n775), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n655), .A2(new_n912), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n913), .A2(new_n634), .A3(new_n685), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n791), .A2(new_n652), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n648), .A2(new_n915), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT62), .Z(new_n917));
  NOR2_X1   g731(.A1(new_n733), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n748), .A2(new_n914), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n448), .B(KEYINPUT125), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n483), .B(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n919), .A2(new_n412), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n717), .A2(new_n655), .A3(new_n633), .A4(new_n680), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n707), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n733), .A2(new_n915), .A3(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n748), .A2(new_n705), .A3(new_n925), .A4(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n921), .B1(new_n928), .B2(new_n412), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n911), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n909), .B1(new_n921), .B2(new_n274), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n930), .B1(new_n412), .B2(new_n931), .ZN(G72));
  XOR2_X1   g746(.A(new_n642), .B(KEYINPUT63), .Z(new_n933));
  INV_X1    g747(.A(new_n905), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n928), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n484), .A3(new_n490), .ZN(new_n936));
  INV_X1    g750(.A(new_n818), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n520), .A2(new_n491), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n938), .A3(new_n933), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n933), .B1(new_n919), .B2(new_n934), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n485), .A3(new_n506), .ZN(new_n941));
  AND4_X1   g755(.A1(new_n857), .A2(new_n936), .A3(new_n939), .A4(new_n941), .ZN(G57));
endmodule


