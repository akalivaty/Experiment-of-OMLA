//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G20), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  NOR2_X1   g0013(.A1(G58), .A2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT65), .B(G244), .Z(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n209), .B1(new_n213), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G50), .B(G58), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(KEYINPUT13), .ZN(new_n245));
  OR2_X1    g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G232), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G1698), .ZN(new_n250));
  OAI211_X1 g0050(.A(new_n248), .B(new_n250), .C1(G226), .C2(G1698), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G97), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G45), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n203), .A2(G274), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G238), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n255), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n265), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n245), .B1(new_n257), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n255), .B1(new_n251), .B2(new_n252), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n272), .A2(new_n269), .A3(KEYINPUT13), .ZN(new_n273));
  OAI21_X1  g0073(.A(G169), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT14), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n257), .A2(new_n245), .A3(new_n270), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT13), .B1(new_n272), .B2(new_n269), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT14), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(new_n279), .A3(G169), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT74), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(KEYINPUT74), .B(KEYINPUT13), .C1(new_n272), .C2(new_n269), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n282), .A2(new_n276), .A3(G179), .A4(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n275), .A2(new_n280), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n210), .ZN(new_n287));
  INV_X1    g0087(.A(G50), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n288), .A2(G20), .A3(G33), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT75), .ZN(new_n290));
  INV_X1    g0090(.A(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n293), .A2(new_n218), .B1(new_n204), .B2(G68), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n287), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT11), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(KEYINPUT11), .B(new_n287), .C1(new_n290), .C2(new_n294), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT12), .B1(new_n299), .B2(G68), .ZN(new_n300));
  OR3_X1    g0100(.A1(new_n299), .A2(KEYINPUT12), .A3(G68), .ZN(new_n301));
  INV_X1    g0101(.A(new_n299), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(new_n287), .ZN(new_n303));
  INV_X1    g0103(.A(G68), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n203), .B2(G20), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n300), .A2(new_n301), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n297), .A2(new_n298), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n285), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n307), .B1(new_n278), .B2(G200), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n282), .A2(new_n276), .A3(G190), .A4(new_n283), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g0112(.A(new_n312), .B(KEYINPUT76), .Z(new_n313));
  NAND3_X1  g0113(.A1(new_n248), .A2(G223), .A3(G1698), .ZN(new_n314));
  INV_X1    g0114(.A(G1698), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n248), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G222), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n314), .B1(new_n218), .B2(new_n248), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n256), .ZN(new_n319));
  INV_X1    g0119(.A(new_n265), .ZN(new_n320));
  INV_X1    g0120(.A(G226), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n268), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT69), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OR3_X1    g0123(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT69), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(G179), .ZN(new_n326));
  NOR2_X1   g0126(.A1(G20), .A2(G33), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G150), .ZN(new_n328));
  NOR3_X1   g0128(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n329));
  NOR2_X1   g0129(.A1(KEYINPUT8), .A2(G58), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT70), .B(G58), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(KEYINPUT8), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n328), .B1(new_n204), .B2(new_n329), .C1(new_n333), .C2(new_n293), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(new_n287), .B1(new_n288), .B2(new_n302), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n303), .A2(KEYINPUT71), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n303), .A2(KEYINPUT71), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n203), .A2(G20), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n335), .B1(new_n288), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n325), .A2(new_n341), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n326), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n248), .A2(G238), .A3(G1698), .ZN(new_n344));
  INV_X1    g0144(.A(G107), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n344), .B1(new_n345), .B2(new_n248), .C1(new_n316), .C2(new_n249), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n256), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n268), .A2(new_n217), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n320), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n287), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(new_n292), .B1(G20), .B2(G77), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT8), .B(G58), .Z(new_n358));
  OR2_X1    g0158(.A1(new_n327), .A2(KEYINPUT72), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n327), .A2(KEYINPUT72), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n354), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n303), .A2(G77), .A3(new_n338), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT73), .B1(new_n302), .B2(new_n218), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n302), .A2(KEYINPUT73), .A3(new_n218), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n350), .B2(new_n341), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n353), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n350), .A2(G200), .ZN(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n370), .B(new_n367), .C1(new_n371), .C2(new_n350), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT9), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n340), .B(new_n374), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n325), .A2(new_n371), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n325), .A2(G200), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT10), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n340), .B(KEYINPUT9), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT10), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(new_n377), .A4(new_n376), .ZN(new_n382));
  AOI211_X1 g0182(.A(new_n343), .B(new_n373), .C1(new_n379), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n321), .A2(G1698), .ZN(new_n384));
  AND2_X1   g0184(.A1(KEYINPUT3), .A2(G33), .ZN(new_n385));
  NOR2_X1   g0185(.A1(KEYINPUT3), .A2(G33), .ZN(new_n386));
  OAI221_X1 g0186(.A(new_n384), .B1(G223), .B2(G1698), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G87), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n256), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n255), .A2(G232), .A3(new_n267), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n265), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n371), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G200), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n255), .B1(new_n387), .B2(new_n388), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n265), .A2(new_n391), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT79), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n393), .A2(new_n397), .A3(KEYINPUT79), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n248), .B2(G20), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n385), .A2(new_n386), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n304), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n327), .A2(G159), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT77), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT77), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n327), .A2(new_n409), .A3(G159), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n214), .B1(new_n331), .B2(G68), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n204), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT16), .B1(new_n406), .B2(new_n413), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n248), .A2(new_n402), .A3(G20), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT7), .B1(new_n404), .B2(new_n204), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(KEYINPUT70), .A2(G58), .ZN(new_n418));
  NOR2_X1   g0218(.A1(KEYINPUT70), .A2(G58), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n215), .B1(new_n420), .B2(new_n304), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(G20), .B1(new_n408), .B2(new_n410), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT16), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n417), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n354), .B1(new_n414), .B2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n336), .A2(new_n332), .A3(new_n337), .A4(new_n338), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n333), .A2(new_n302), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n401), .A2(KEYINPUT17), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT17), .B1(new_n401), .B2(new_n429), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n428), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n414), .A2(new_n424), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(new_n354), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n395), .A2(new_n396), .A3(G179), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n390), .A2(new_n392), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n436), .B1(new_n341), .B2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n435), .A2(KEYINPUT78), .A3(KEYINPUT18), .A4(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(KEYINPUT18), .B(new_n438), .C1(new_n425), .C2(new_n428), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT78), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n438), .B1(new_n425), .B2(new_n428), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n439), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n432), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n313), .A2(new_n383), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT21), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT5), .B(G41), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n258), .A2(G1), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(G274), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n451), .A2(new_n452), .B1(new_n211), .B2(new_n254), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(G270), .B2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(G264), .B(G1698), .C1(new_n385), .C2(new_n386), .ZN(new_n457));
  OAI211_X1 g0257(.A(G257), .B(new_n315), .C1(new_n385), .C2(new_n386), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n246), .A2(G303), .A3(new_n247), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n460), .A2(KEYINPUT84), .A3(new_n256), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT84), .B1(new_n460), .B2(new_n256), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G169), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n299), .A2(G116), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n203), .A2(G33), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n299), .A2(new_n466), .A3(new_n210), .A4(new_n286), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n468), .B2(G116), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  AND2_X1   g0271(.A1(KEYINPUT81), .A2(G97), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT81), .A2(G97), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n204), .B(new_n471), .C1(new_n474), .C2(G33), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G20), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n287), .A2(KEYINPUT85), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT85), .B1(new_n287), .B2(new_n477), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT20), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n475), .B(KEYINPUT20), .C1(new_n479), .C2(new_n480), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n470), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n450), .B1(new_n464), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n484), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n287), .A2(new_n477), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT85), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n478), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT20), .B1(new_n491), .B2(new_n475), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n469), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n455), .A2(G270), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n453), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n460), .A2(new_n256), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT84), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n460), .A2(KEYINPUT84), .A3(new_n256), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n493), .A2(G179), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n493), .A2(KEYINPUT21), .A3(G169), .A4(new_n463), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n456), .B(G190), .C1(new_n461), .C2(new_n462), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n485), .B(new_n503), .C1(new_n500), .C2(new_n394), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n486), .A2(new_n501), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(G257), .B(G1698), .C1(new_n385), .C2(new_n386), .ZN(new_n507));
  OAI211_X1 g0307(.A(G250), .B(new_n315), .C1(new_n385), .C2(new_n386), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G294), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(new_n256), .B1(new_n455), .B2(G264), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n453), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n341), .ZN(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n248), .A2(new_n514), .A3(new_n204), .A4(G87), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n204), .B(G87), .C1(new_n385), .C2(new_n386), .ZN(new_n516));
  XOR2_X1   g0316(.A(KEYINPUT86), .B(KEYINPUT22), .Z(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(G20), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT23), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n204), .B2(G107), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n345), .A2(KEYINPUT23), .A3(G20), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n515), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT24), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT24), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n515), .A2(new_n518), .A3(new_n527), .A4(new_n524), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n354), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n302), .A2(KEYINPUT25), .A3(new_n345), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT25), .B1(new_n302), .B2(new_n345), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n530), .A2(new_n531), .B1(new_n345), .B2(new_n467), .ZN(new_n532));
  OAI221_X1 g0332(.A(new_n513), .B1(G179), .B2(new_n512), .C1(new_n529), .C2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n529), .A2(new_n532), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n512), .A2(new_n394), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n511), .A2(new_n371), .A3(new_n453), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n345), .B1(new_n403), .B2(new_n405), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n327), .A2(G77), .ZN(new_n542));
  OR2_X1    g0342(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n543));
  NAND2_X1  g0343(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n544));
  AOI21_X1  g0344(.A(G107), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n473), .ZN(new_n546));
  NAND2_X1  g0346(.A1(KEYINPUT81), .A2(G97), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n544), .ZN(new_n549));
  NOR2_X1   g0349(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g0351(.A(G97), .B(G107), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n545), .A2(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n542), .B1(new_n553), .B2(new_n204), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n541), .B1(new_n554), .B2(KEYINPUT82), .ZN(new_n555));
  AND2_X1   g0355(.A1(G97), .A2(G107), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n543), .B(new_n544), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n345), .B1(new_n549), .B2(new_n550), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(new_n474), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(G20), .B1(G77), .B2(new_n327), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT82), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n354), .B1(new_n555), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(G97), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n302), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n467), .B2(new_n565), .ZN(new_n567));
  OAI211_X1 g0367(.A(G244), .B(new_n315), .C1(new_n385), .C2(new_n386), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT4), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT83), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT83), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(new_n572), .A3(new_n569), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n248), .A2(KEYINPUT4), .A3(G244), .A4(new_n315), .ZN(new_n574));
  OAI211_X1 g0374(.A(G250), .B(G1698), .C1(new_n385), .C2(new_n386), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n575), .A2(new_n471), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n571), .A2(new_n573), .A3(new_n574), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n256), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n451), .A2(new_n452), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(G257), .A3(new_n255), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n453), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n341), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  AOI211_X1 g0383(.A(new_n352), .B(new_n581), .C1(new_n577), .C2(new_n256), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n564), .A2(new_n567), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n541), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n561), .B2(new_n562), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n554), .A2(KEYINPUT82), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n287), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n567), .ZN(new_n590));
  AOI21_X1  g0390(.A(G200), .B1(new_n578), .B2(new_n582), .ZN(new_n591));
  AOI211_X1 g0391(.A(G190), .B(new_n581), .C1(new_n577), .C2(new_n256), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n589), .B(new_n590), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n356), .A2(new_n299), .ZN(new_n594));
  INV_X1    g0394(.A(G87), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n467), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n546), .A2(new_n595), .A3(new_n345), .A4(new_n547), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT19), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n204), .B1(new_n252), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n598), .B1(new_n474), .B2(new_n293), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n248), .A2(new_n204), .A3(G68), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI211_X1 g0403(.A(new_n594), .B(new_n596), .C1(new_n603), .C2(new_n287), .ZN(new_n604));
  OAI211_X1 g0404(.A(G244), .B(G1698), .C1(new_n385), .C2(new_n386), .ZN(new_n605));
  OAI211_X1 g0405(.A(G238), .B(new_n315), .C1(new_n385), .C2(new_n386), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(new_n519), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n256), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n264), .A2(G45), .ZN(new_n609));
  OAI21_X1  g0409(.A(G250), .B1(new_n258), .B2(G1), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n256), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G200), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n611), .B1(new_n607), .B2(new_n256), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G190), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n604), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n603), .A2(new_n287), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n468), .A2(new_n356), .ZN(new_n619));
  INV_X1    g0419(.A(new_n594), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n613), .A2(new_n341), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n615), .A2(new_n352), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n585), .A2(new_n593), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n449), .A2(new_n506), .A3(new_n540), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n628), .B(KEYINPUT87), .ZN(G372));
  INV_X1    g0429(.A(new_n624), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n617), .A2(new_n624), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n631), .B1(new_n585), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n471), .B(new_n575), .C1(new_n568), .C2(new_n569), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n572), .B1(new_n568), .B2(new_n569), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n255), .B1(new_n636), .B2(new_n573), .ZN(new_n637));
  OAI21_X1  g0437(.A(G169), .B1(new_n637), .B2(new_n581), .ZN(new_n638));
  INV_X1    g0438(.A(new_n573), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n639), .A2(new_n634), .A3(new_n635), .ZN(new_n640));
  OAI211_X1 g0440(.A(G179), .B(new_n582), .C1(new_n640), .C2(new_n255), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n589), .A2(new_n590), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(KEYINPUT26), .A3(new_n625), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n630), .B1(new_n633), .B2(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n486), .A2(new_n533), .A3(new_n501), .A4(new_n502), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n585), .A2(new_n593), .A3(new_n625), .A4(new_n538), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n449), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT88), .ZN(new_n649));
  INV_X1    g0449(.A(new_n343), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n445), .A2(new_n440), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT89), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT89), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n445), .A2(new_n653), .A3(new_n440), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n311), .A2(new_n353), .A3(new_n368), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT90), .B1(new_n308), .B2(new_n657), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n658), .A2(new_n431), .A3(new_n430), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n308), .A2(new_n657), .A3(KEYINPUT90), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n656), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n379), .A2(new_n382), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n650), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n649), .A2(new_n665), .ZN(G369));
  NAND3_X1  g0466(.A1(new_n486), .A2(new_n501), .A3(new_n502), .ZN(new_n667));
  INV_X1    g0467(.A(G13), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n668), .A2(G1), .A3(G20), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT91), .B1(new_n670), .B2(KEYINPUT27), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(KEYINPUT91), .A3(KEYINPUT27), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(G213), .B1(new_n670), .B2(KEYINPUT27), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n485), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n667), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n505), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n540), .B1(new_n534), .B2(new_n677), .ZN(new_n683));
  INV_X1    g0483(.A(new_n533), .ZN(new_n684));
  INV_X1    g0484(.A(new_n677), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n667), .A2(new_n677), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n539), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n684), .B2(new_n677), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n207), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n203), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n597), .A2(G116), .ZN(new_n696));
  INV_X1    g0496(.A(new_n216), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n695), .A2(new_n696), .B1(new_n697), .B2(new_n694), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT28), .Z(new_n699));
  NAND2_X1  g0499(.A1(new_n647), .A2(new_n677), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G330), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n511), .A2(new_n615), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n500), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n705), .B1(new_n707), .B2(new_n641), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n511), .A2(new_n615), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n463), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n584), .A3(KEYINPUT30), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n578), .A2(new_n582), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n615), .A2(G179), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n712), .A2(new_n463), .A3(new_n512), .A4(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n708), .A2(new_n711), .A3(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n715), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT31), .B1(new_n715), .B2(new_n685), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n627), .A2(new_n506), .A3(new_n540), .A4(new_n677), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n704), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n703), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n699), .B1(new_n721), .B2(G1), .ZN(G364));
  NOR2_X1   g0522(.A1(new_n668), .A2(G20), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G45), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT92), .Z(new_n725));
  NAND2_X1  g0525(.A1(new_n695), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n682), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(G330), .B2(new_n680), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n210), .B1(G20), .B2(new_n341), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n204), .A2(new_n352), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G200), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G190), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(KEYINPUT33), .B(G317), .Z(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n204), .A2(G190), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR4_X1   g0544(.A1(new_n204), .A2(new_n371), .A3(new_n394), .A4(G179), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G329), .A2(new_n744), .B1(new_n745), .B2(G303), .ZN(new_n746));
  INV_X1    g0546(.A(G322), .ZN(new_n747));
  INV_X1    g0547(.A(new_n735), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n748), .A2(new_n371), .A3(G200), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n746), .B(new_n404), .C1(new_n747), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n736), .A2(new_n371), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n740), .B(new_n751), .C1(G326), .C2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n748), .A2(G190), .A3(G200), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n754), .A2(KEYINPUT97), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(KEYINPUT97), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR4_X1   g0558(.A1(new_n204), .A2(new_n394), .A3(G179), .A4(G190), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n759), .A2(KEYINPUT98), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(KEYINPUT98), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n758), .A2(G311), .B1(new_n763), .B2(G283), .ZN(new_n764));
  INV_X1    g0564(.A(G294), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n204), .B1(new_n742), .B2(G190), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n766), .A2(KEYINPUT99), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(KEYINPUT99), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n753), .B(new_n764), .C1(new_n765), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n745), .A2(G87), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n248), .B(new_n771), .C1(new_n750), .C2(new_n420), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n758), .B2(G77), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n762), .A2(new_n345), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n769), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G97), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n744), .A2(G159), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  INV_X1    g0579(.A(new_n752), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n288), .A2(new_n780), .B1(new_n738), .B2(new_n304), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n773), .A2(new_n775), .A3(new_n777), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n734), .B1(new_n770), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n204), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT94), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n734), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT96), .Z(new_n789));
  NAND2_X1  g0589(.A1(new_n207), .A2(new_n404), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT93), .Z(new_n791));
  AND2_X1   g0591(.A1(new_n259), .A2(new_n261), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n791), .B1(new_n216), .B2(new_n793), .C1(new_n240), .C2(new_n258), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n693), .A2(new_n404), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n795), .A2(G355), .B1(new_n476), .B2(new_n693), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n789), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n784), .A2(new_n726), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n787), .B(KEYINPUT100), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n680), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n729), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  NOR2_X1   g0602(.A1(new_n373), .A2(new_n685), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n585), .A2(new_n631), .A3(new_n632), .ZN(new_n804));
  AOI21_X1  g0604(.A(KEYINPUT26), .B1(new_n642), .B2(new_n625), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n624), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n646), .A2(new_n645), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n700), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n677), .A2(new_n367), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n372), .A2(new_n810), .B1(new_n353), .B2(new_n368), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n369), .A2(new_n685), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n808), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n720), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n727), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n758), .A2(G116), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n763), .A2(G87), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G283), .A2(new_n737), .B1(new_n752), .B2(G303), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n248), .B1(new_n749), .B2(G294), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G311), .A2(new_n744), .B1(new_n745), .B2(G107), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n818), .A2(new_n819), .A3(new_n823), .A4(new_n777), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n749), .A2(G143), .B1(new_n752), .B2(G137), .ZN(new_n825));
  INV_X1    g0625(.A(G150), .ZN(new_n826));
  INV_X1    g0626(.A(G159), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n738), .C1(new_n757), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n776), .A2(new_n331), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  INV_X1    g0632(.A(new_n745), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n248), .B1(new_n743), .B2(new_n832), .C1(new_n833), .C2(new_n288), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n763), .B2(G68), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n830), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n824), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n734), .B1(new_n839), .B2(KEYINPUT101), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(KEYINPUT101), .B2(new_n839), .ZN(new_n841));
  INV_X1    g0641(.A(new_n813), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n785), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n733), .A2(new_n785), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n726), .B1(new_n844), .B2(new_n218), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n841), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n817), .A2(new_n846), .ZN(G384));
  NOR2_X1   g0647(.A1(new_n723), .A2(new_n203), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT38), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n676), .B1(new_n425), .B2(new_n428), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n655), .B2(new_n432), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT102), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n393), .A2(new_n397), .A3(KEYINPUT79), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(new_n398), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n443), .B(new_n850), .C1(new_n435), .C2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n852), .B1(new_n855), .B2(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n401), .A2(new_n429), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(new_n443), .A4(new_n850), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n856), .B1(new_n861), .B2(new_n852), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n849), .B1(new_n851), .B2(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(KEYINPUT38), .B(new_n861), .C1(new_n447), .C2(new_n850), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT39), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n861), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n850), .B1(new_n432), .B2(new_n446), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n849), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n864), .A2(new_n868), .A3(KEYINPUT39), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n308), .A2(new_n685), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  OR3_X1    g0671(.A1(new_n865), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n655), .A2(new_n676), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n864), .A2(new_n868), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n685), .A2(new_n307), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n308), .A2(new_n311), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n311), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n307), .B(new_n685), .C1(new_n877), .C2(new_n285), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n812), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n808), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n873), .B1(new_n874), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n872), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n448), .B1(new_n701), .B2(new_n702), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n884), .A2(new_n664), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n883), .B(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n879), .A2(new_n842), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n718), .A2(new_n719), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT40), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n889), .A2(new_n890), .A3(new_n874), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n863), .A2(new_n864), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n890), .B1(new_n892), .B2(new_n889), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n449), .A2(new_n888), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n889), .A2(new_n890), .A3(new_n874), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n887), .A2(new_n888), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n864), .B2(new_n863), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(new_n899), .B2(new_n890), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(new_n449), .A3(new_n888), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n896), .A2(new_n901), .A3(G330), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n848), .B1(new_n886), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n886), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n213), .A2(new_n476), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT36), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n697), .B(G77), .C1(new_n304), .C2(new_n420), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(G50), .B2(new_n304), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(G1), .A3(new_n668), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n904), .A2(new_n909), .A3(new_n912), .ZN(G367));
  NOR2_X1   g0713(.A1(new_n677), .A2(new_n604), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n624), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n625), .B2(new_n914), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT103), .ZN(new_n917));
  INV_X1    g0717(.A(new_n799), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n791), .A2(new_n235), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n788), .B1(new_n693), .B2(new_n356), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n726), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(G137), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n833), .A2(new_n420), .B1(new_n923), .B2(new_n743), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(G143), .B2(new_n752), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n925), .B1(new_n827), .B2(new_n738), .C1(new_n757), .C2(new_n288), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n763), .A2(G77), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n248), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n926), .B1(new_n928), .B2(KEYINPUT109), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(KEYINPUT109), .B2(new_n928), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n769), .A2(new_n304), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(G150), .B2(new_n749), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT108), .Z(new_n933));
  INV_X1    g0733(.A(G303), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n404), .B1(new_n750), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(G317), .B2(new_n744), .ZN(new_n936));
  INV_X1    g0736(.A(G283), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n936), .B1(new_n937), .B2(new_n757), .C1(new_n474), .C2(new_n762), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n833), .A2(new_n476), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(KEYINPUT46), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G311), .B2(new_n752), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n939), .A2(KEYINPUT46), .B1(new_n737), .B2(G294), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n941), .B(new_n942), .C1(new_n345), .C2(new_n769), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n930), .A2(new_n933), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT47), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n733), .B1(new_n944), .B2(new_n945), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n919), .B(new_n922), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n725), .A2(G1), .ZN(new_n949));
  INV_X1    g0749(.A(new_n690), .ZN(new_n950));
  INV_X1    g0750(.A(new_n689), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n950), .B1(new_n687), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT106), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(new_n681), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n681), .B(new_n953), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n954), .B1(new_n955), .B2(new_n952), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n721), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT107), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n642), .A2(new_n685), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT105), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n960), .B(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n685), .B1(new_n564), .B2(new_n567), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n585), .A2(new_n593), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n691), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT45), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT44), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n965), .A2(new_n691), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n965), .B2(new_n691), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n968), .A2(new_n688), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n688), .B1(new_n968), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n721), .A2(new_n956), .A3(KEYINPUT107), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n959), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n721), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n694), .B(KEYINPUT41), .Z(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n949), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n965), .A2(new_n690), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT42), .Z(new_n983));
  AOI21_X1  g0783(.A(new_n533), .B1(new_n962), .B2(new_n964), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n677), .B1(new_n984), .B2(new_n642), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT43), .B1(new_n917), .B2(KEYINPUT104), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(KEYINPUT104), .B2(new_n917), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT43), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n986), .B(new_n988), .C1(new_n990), .C2(new_n917), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n688), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n965), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n992), .B(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n948), .B1(new_n981), .B2(new_n995), .ZN(G387));
  NAND3_X1  g0796(.A1(new_n683), .A2(new_n686), .A3(new_n918), .ZN(new_n997));
  INV_X1    g0797(.A(new_n795), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n998), .A2(new_n696), .B1(G107), .B2(new_n207), .ZN(new_n999));
  INV_X1    g0799(.A(new_n791), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n232), .B2(new_n793), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n696), .B(new_n258), .C1(new_n304), .C2(new_n218), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT110), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(KEYINPUT110), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n358), .A2(new_n288), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT50), .Z(new_n1006));
  NAND3_X1  g0806(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n999), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n727), .B1(new_n1008), .B2(new_n789), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n769), .A2(new_n355), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n404), .B1(new_n745), .B2(G77), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n826), .B2(new_n743), .C1(new_n750), .C2(new_n288), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(G159), .C2(new_n752), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n758), .A2(G68), .B1(new_n763), .B2(G97), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n333), .C2(new_n738), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G317), .A2(new_n749), .B1(new_n737), .B2(G311), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n747), .B2(new_n780), .C1(new_n757), .C2(new_n934), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT48), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n769), .A2(new_n937), .B1(new_n765), .B2(new_n833), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT111), .Z(new_n1020));
  NAND3_X1  g0820(.A1(new_n1018), .A2(KEYINPUT49), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n248), .B1(new_n744), .B2(G326), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(new_n476), .C2(new_n762), .ZN(new_n1023));
  AOI21_X1  g0823(.A(KEYINPUT49), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1015), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1009), .B1(new_n1025), .B2(new_n733), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n956), .A2(new_n949), .B1(new_n997), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n957), .A2(new_n694), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n721), .A2(new_n956), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(G393));
  INV_X1    g0830(.A(new_n694), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n975), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(new_n957), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1033), .A2(new_n977), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1000), .A2(new_n243), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n734), .B(new_n787), .C1(new_n207), .C2(new_n474), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n727), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n749), .A2(G159), .B1(new_n752), .B2(G150), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT51), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n758), .A2(new_n358), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n819), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n769), .A2(new_n218), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n404), .B1(new_n744), .B2(G143), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n833), .B2(new_n304), .C1(new_n738), .C2(new_n288), .ZN(new_n1044));
  OR4_X1    g0844(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n758), .A2(G294), .B1(G303), .B2(new_n737), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n476), .B2(new_n769), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT112), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n749), .A2(G311), .B1(new_n752), .B2(G317), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT52), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n404), .B1(new_n743), .B2(new_n747), .C1(new_n833), .C2(new_n937), .ZN(new_n1051));
  OR3_X1    g0851(.A1(new_n1050), .A2(new_n774), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1045), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1037), .B1(new_n1053), .B2(new_n733), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n787), .B2(new_n965), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n949), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n1032), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1034), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(G390));
  INV_X1    g0859(.A(KEYINPUT113), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n881), .B2(new_n870), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n812), .B1(new_n647), .B2(new_n803), .ZN(new_n1062));
  OAI211_X1 g0862(.A(KEYINPUT113), .B(new_n871), .C1(new_n1062), .C2(new_n879), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(new_n865), .C2(new_n869), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n892), .B(new_n871), .C1(new_n879), .C2(new_n1062), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n715), .A2(new_n685), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT31), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n715), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n626), .A2(new_n505), .A3(new_n539), .A4(new_n685), .ZN(new_n1072));
  OAI211_X1 g0872(.A(G330), .B(new_n813), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1073), .A2(new_n879), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1066), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1074), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1064), .A2(new_n1065), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n1056), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n785), .B1(new_n865), .B2(new_n869), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n844), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n727), .B1(new_n1081), .B2(new_n332), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n750), .A2(new_n476), .B1(new_n780), .B2(new_n937), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1042), .B(new_n1083), .C1(G107), .C2(new_n737), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n771), .A2(new_n404), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT116), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(new_n474), .C2(new_n757), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n762), .A2(new_n304), .B1(new_n765), .B2(new_n743), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT117), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n745), .A2(G150), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT53), .Z(new_n1091));
  XNOR2_X1  g0891(.A(KEYINPUT54), .B(G143), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1091), .B1(new_n762), .B2(new_n288), .C1(new_n757), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(G128), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1094), .A2(new_n780), .B1(new_n738), .B2(new_n923), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n404), .B1(new_n744), .B2(G125), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n750), .B2(new_n832), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n827), .B2(new_n769), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1087), .A2(new_n1089), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1082), .B1(new_n1100), .B2(new_n733), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1079), .B1(new_n1080), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1062), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n879), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n720), .B2(new_n813), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1103), .B1(new_n1105), .B2(new_n1074), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT114), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT115), .B1(new_n1073), .B2(new_n879), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1073), .A2(new_n879), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1073), .A2(KEYINPUT115), .A3(new_n879), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n1062), .A3(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(KEYINPUT114), .B(new_n1103), .C1(new_n1105), .C2(new_n1074), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1108), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n448), .A2(new_n815), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n884), .A2(new_n664), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1078), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1075), .A2(new_n1077), .A3(new_n1117), .A4(new_n1115), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n694), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1102), .A2(new_n1121), .ZN(G378));
  NAND2_X1  g0922(.A1(new_n340), .A2(new_n676), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n663), .A2(new_n343), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n662), .B2(new_n650), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OR3_X1    g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n900), .A2(new_n1131), .A3(G330), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n900), .B2(G330), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n883), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n1132), .A2(new_n1133), .B1(new_n1134), .B2(KEYINPUT120), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1129), .B(new_n1130), .C1(new_n894), .C2(new_n704), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT120), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n900), .A2(new_n1131), .A3(G330), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n883), .A4(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n949), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n727), .B1(new_n1081), .B2(G50), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n931), .B1(G116), .B2(new_n752), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT118), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n404), .A2(new_n262), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n749), .B2(G107), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G283), .A2(new_n744), .B1(new_n745), .B2(G77), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n565), .C2(new_n738), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n763), .A2(new_n331), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n757), .B2(new_n355), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1144), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(G50), .B1(new_n291), .B2(new_n262), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1151), .A2(KEYINPUT58), .B1(new_n1145), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n752), .A2(G125), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n833), .B2(new_n1092), .C1(new_n750), .C2(new_n1094), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G132), .B2(new_n737), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n923), .B2(new_n757), .C1(new_n826), .C2(new_n769), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1158));
  AOI211_X1 g0958(.A(G33), .B(G41), .C1(new_n744), .C2(G124), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(new_n827), .C2(new_n762), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1153), .B1(KEYINPUT58), .B2(new_n1151), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1142), .B1(new_n1162), .B2(new_n733), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n785), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1131), .B2(new_n1164), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT119), .Z(new_n1166));
  NAND2_X1  g0966(.A1(new_n1141), .A2(new_n1166), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1120), .A2(KEYINPUT121), .A3(new_n1117), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT121), .B1(new_n1120), .B2(new_n1117), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1140), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT121), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1064), .A2(new_n1065), .A3(new_n1076), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1076), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1118), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1117), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1173), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1120), .A2(KEYINPUT121), .A3(new_n1117), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n883), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1136), .A2(new_n1134), .A3(new_n1138), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1171), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1031), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1167), .B1(new_n1172), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(G375));
  OR2_X1    g0986(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1187), .A2(new_n980), .A3(new_n1118), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n879), .A2(new_n785), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n727), .B1(new_n1081), .B2(G68), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n758), .A2(G150), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n832), .A2(new_n780), .B1(new_n738), .B2(new_n1092), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n750), .A2(new_n923), .B1(new_n827), .B2(new_n833), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n248), .B1(new_n743), .B2(new_n1094), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n776), .A2(G50), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1191), .A2(new_n1195), .A3(new_n1149), .A4(new_n1196), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n476), .A2(new_n738), .B1(new_n780), .B2(new_n765), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n750), .A2(new_n937), .B1(new_n565), .B2(new_n833), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n404), .B1(new_n743), .B2(new_n934), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1201), .B(new_n927), .C1(new_n345), .C2(new_n757), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1197), .B1(new_n1202), .B2(new_n1010), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1190), .B1(new_n1203), .B2(new_n733), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1115), .A2(new_n949), .B1(new_n1189), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1188), .A2(new_n1205), .ZN(G381));
  OR3_X1    g1006(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(G390), .A2(G387), .A3(G381), .A4(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT122), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(G375), .A2(G378), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(G407));
  INV_X1    g1011(.A(G343), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(G213), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT123), .Z(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(G407), .A2(G213), .A3(new_n1215), .ZN(G409));
  AND2_X1   g1016(.A1(G387), .A2(new_n1058), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(G387), .A2(new_n1058), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(G393), .B(G396), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(G387), .A2(new_n1058), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT127), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1220), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1219), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1219), .A2(new_n1223), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1165), .B1(new_n1056), .B2(new_n1227), .C1(new_n1170), .C2(new_n979), .ZN(new_n1228));
  INV_X1    g1028(.A(G378), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT124), .B1(new_n1185), .B2(G378), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1183), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n694), .B(new_n1232), .C1(new_n1234), .C2(KEYINPUT57), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1167), .ZN(new_n1236));
  AND4_X1   g1036(.A1(KEYINPUT124), .A2(new_n1235), .A3(G378), .A4(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1230), .B1(new_n1231), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G384), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(KEYINPUT126), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1187), .A2(KEYINPUT125), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1241), .B(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n694), .A3(new_n1118), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1240), .B1(new_n1244), .B2(new_n1205), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT126), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(G384), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1244), .A2(KEYINPUT126), .A3(new_n1239), .A4(new_n1205), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1238), .A2(new_n1213), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT62), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1235), .A2(G378), .A3(new_n1236), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1185), .A2(KEYINPUT124), .A3(G378), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1214), .B1(new_n1256), .B2(new_n1230), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1251), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1250), .A2(new_n1251), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1214), .A2(G2897), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1247), .A2(new_n1248), .A3(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1212), .A2(G213), .A3(G2897), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1260), .B1(new_n1265), .B2(new_n1257), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1226), .B1(new_n1259), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1238), .A2(new_n1213), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1250), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1257), .A2(KEYINPUT63), .A3(new_n1249), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1226), .A2(KEYINPUT61), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1269), .A2(new_n1271), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1267), .A2(new_n1274), .ZN(G405));
  NAND2_X1  g1075(.A1(G375), .A2(new_n1229), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1226), .A2(new_n1256), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1256), .A2(new_n1276), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(new_n1225), .A3(new_n1224), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1249), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1280), .B(new_n1281), .ZN(G402));
endmodule


