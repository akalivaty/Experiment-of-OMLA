//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n440, new_n441, new_n445, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n590, new_n591, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n640, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  AND2_X1   g014(.A1(KEYINPUT64), .A2(G57), .ZN(new_n440));
  NOR2_X1   g015(.A1(KEYINPUT64), .A2(G57), .ZN(new_n441));
  NOR2_X1   g016(.A1(new_n440), .A2(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR3_X1   g029(.A1(G235), .A2(G238), .A3(G236), .ZN(new_n455));
  OAI21_X1  g030(.A(new_n455), .B1(new_n441), .B2(new_n440), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n454), .A2(new_n460), .B1(new_n461), .B2(new_n457), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT67), .Z(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n467), .A2(KEYINPUT68), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT68), .B1(new_n467), .B2(new_n470), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n464), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR3_X1   g050(.A1(new_n471), .A2(new_n472), .A3(new_n475), .ZN(G160));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n468), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n464), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G138), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT3), .B(G2104), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n490), .A2(new_n491), .A3(G138), .A4(new_n464), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n464), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT69), .A4(G2104), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n497), .A2(new_n501), .B1(new_n482), .B2(G126), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT70), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(new_n506), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n512), .B1(new_n513), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n519), .A2(G50), .A3(G543), .A4(new_n520), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT71), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n525), .A2(KEYINPUT71), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(G166));
  INV_X1    g103(.A(new_n523), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n519), .A2(G543), .A3(new_n520), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n529), .A2(G89), .B1(new_n530), .B2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(KEYINPUT73), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(KEYINPUT73), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n533), .A2(new_n537), .A3(new_n534), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n539));
  NOR3_X1   g114(.A1(new_n507), .A2(new_n508), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT72), .B1(new_n521), .B2(new_n506), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(G63), .A2(G651), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n536), .A2(new_n538), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n531), .A2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(new_n522), .A2(new_n539), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n521), .A2(KEYINPUT72), .A3(new_n506), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n547), .A2(G64), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n514), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n519), .A2(G543), .A3(new_n520), .ZN(new_n553));
  XOR2_X1   g128(.A(KEYINPUT74), .B(G90), .Z(new_n554));
  OAI22_X1  g129(.A1(new_n552), .A2(new_n553), .B1(new_n523), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n551), .A2(new_n555), .ZN(G171));
  NAND2_X1  g131(.A1(new_n542), .A2(G56), .ZN(new_n557));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n514), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G43), .ZN(new_n560));
  INV_X1    g135(.A(G81), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n560), .A2(new_n553), .B1(new_n523), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n553), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n515), .A2(new_n518), .B1(KEYINPUT6), .B2(new_n514), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n571), .A2(new_n572), .A3(G53), .A4(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n571), .A2(G91), .A3(new_n522), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n521), .B2(new_n506), .ZN(new_n577));
  AND2_X1   g152(.A1(G78), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n574), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(new_n555), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n549), .A2(new_n550), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT75), .B1(new_n551), .B2(new_n555), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G301));
  XNOR2_X1  g164(.A(new_n525), .B(KEYINPUT71), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n529), .A2(G88), .B1(G651), .B2(new_n511), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G303));
  INV_X1    g167(.A(G74), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n540), .B2(new_n541), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n571), .A2(G87), .A3(new_n522), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n571), .A2(G49), .A3(G543), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(KEYINPUT76), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n595), .A2(new_n600), .A3(new_n596), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G288));
  NAND4_X1  g178(.A1(new_n519), .A2(G86), .A3(new_n520), .A4(new_n522), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n571), .A2(KEYINPUT77), .A3(G86), .A4(new_n522), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(G61), .B1(new_n507), .B2(new_n508), .ZN(new_n609));
  NAND2_X1  g184(.A1(G73), .A2(G543), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n514), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n530), .B2(G48), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n612), .ZN(G305));
  NAND3_X1  g188(.A1(new_n547), .A2(G60), .A3(new_n548), .ZN(new_n614));
  NAND2_X1  g189(.A1(G72), .A2(G543), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G651), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n529), .A2(G85), .B1(new_n530), .B2(G47), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(G290));
  NAND2_X1  g194(.A1(G301), .A2(G868), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(KEYINPUT78), .ZN(new_n621));
  AND2_X1   g196(.A1(new_n620), .A2(KEYINPUT78), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n529), .A2(KEYINPUT10), .A3(G92), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT10), .ZN(new_n624));
  INV_X1    g199(.A(G92), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n523), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(G79), .A2(G543), .ZN(new_n628));
  INV_X1    g203(.A(G66), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n509), .B2(new_n629), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n530), .A2(G54), .B1(new_n630), .B2(G651), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(KEYINPUT79), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(KEYINPUT79), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n621), .B1(new_n622), .B2(new_n637), .ZN(G284));
  AOI21_X1  g213(.A(new_n621), .B1(new_n622), .B2(new_n637), .ZN(G321));
  NAND2_X1  g214(.A1(G299), .A2(new_n636), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G168), .B2(new_n636), .ZN(G297));
  OAI21_X1  g216(.A(new_n640), .B1(G168), .B2(new_n636), .ZN(G280));
  INV_X1    g217(.A(new_n635), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT80), .B(G559), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n643), .B1(G860), .B2(new_n645), .ZN(G148));
  NAND3_X1  g221(.A1(new_n633), .A2(new_n634), .A3(new_n645), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(G868), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g224(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g225(.A1(new_n490), .A2(new_n469), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT12), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT13), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n482), .A2(G123), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT81), .ZN(new_n656));
  OAI21_X1  g231(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n657));
  INV_X1    g232(.A(G111), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n657), .B1(new_n658), .B2(G2105), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n480), .B2(G135), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT82), .B(G2096), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n654), .A2(new_n663), .ZN(G156));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2435), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT84), .B(G2438), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2427), .B(G2430), .Z(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(KEYINPUT14), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1341), .B(G1348), .Z(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2451), .B(G2454), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2443), .B(G2446), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  OR2_X1    g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(G14), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n675), .B2(new_n678), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n679), .A2(new_n681), .ZN(G401));
  INV_X1    g257(.A(KEYINPUT18), .ZN(new_n683));
  XOR2_X1   g258(.A(G2084), .B(G2090), .Z(new_n684));
  XNOR2_X1  g259(.A(G2067), .B(G2678), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(KEYINPUT17), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n684), .A2(new_n685), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G2100), .ZN(new_n690));
  XOR2_X1   g265(.A(G2072), .B(G2078), .Z(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n686), .B2(KEYINPUT18), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(G2096), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n690), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G227));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT86), .Z(new_n699));
  XOR2_X1   g274(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n700));
  XNOR2_X1  g275(.A(G1971), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1956), .B(G2474), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1961), .B(G1966), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT20), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n703), .A2(new_n704), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n702), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n702), .B2(new_n708), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n699), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(G1991), .B(G1996), .Z(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n707), .A2(new_n710), .A3(new_n699), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(new_n712), .B2(new_n715), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n697), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n718), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n720), .A2(new_n696), .A3(new_n716), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n721), .ZN(G229));
  XOR2_X1   g297(.A(KEYINPUT31), .B(G11), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT99), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n661), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G28), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n728));
  AOI21_X1  g303(.A(G29), .B1(new_n727), .B2(KEYINPUT30), .ZN(new_n729));
  AOI211_X1 g304(.A(new_n724), .B(new_n726), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n725), .A2(G32), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n480), .A2(G141), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT96), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n469), .A2(G105), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT97), .Z(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT26), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n482), .A2(G129), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n731), .B1(new_n740), .B2(new_n725), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT27), .B(G1996), .Z(new_n742));
  INV_X1    g317(.A(G2078), .ZN(new_n743));
  NAND2_X1  g318(.A1(G164), .A2(G29), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G27), .B2(G29), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n741), .A2(new_n742), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n730), .B(new_n746), .C1(new_n743), .C2(new_n745), .ZN(new_n747));
  INV_X1    g322(.A(G16), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G21), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G168), .B2(new_n748), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1966), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT24), .ZN(new_n753));
  INV_X1    g328(.A(G34), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n753), .B2(new_n754), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G160), .B2(new_n725), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT95), .B(G2084), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n725), .A2(G35), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G162), .B2(new_n725), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT29), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n752), .B(new_n759), .C1(G2090), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n748), .A2(G4), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n643), .B2(new_n748), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G1348), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n725), .A2(G26), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  INV_X1    g345(.A(G116), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G2105), .ZN(new_n772));
  OAI211_X1 g347(.A(G128), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n490), .A2(KEYINPUT90), .A3(G128), .A4(G2105), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n480), .A2(KEYINPUT89), .A3(G140), .ZN(new_n778));
  OAI211_X1 g353(.A(G140), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT89), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  AND3_X1   g357(.A1(new_n777), .A2(KEYINPUT91), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(KEYINPUT91), .B1(new_n777), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n769), .B1(new_n786), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2067), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n765), .A2(G1348), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n766), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n762), .A2(G2090), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT101), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n725), .A2(G33), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n490), .A2(G127), .ZN(new_n794));
  NAND2_X1  g369(.A1(G115), .A2(G2104), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n464), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(KEYINPUT93), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(KEYINPUT93), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT25), .ZN(new_n799));
  NAND2_X1  g374(.A1(G103), .A2(G2104), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G2105), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n480), .A2(G139), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n797), .A2(new_n798), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n793), .B1(new_n806), .B2(new_n725), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(G2072), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n748), .A2(G20), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT102), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT23), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G299), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1956), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n807), .A2(G2072), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n792), .A2(new_n808), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n741), .A2(new_n742), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT98), .Z(new_n817));
  NOR2_X1   g392(.A1(G5), .A2(G16), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT100), .Z(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G171), .B2(G16), .ZN(new_n820));
  INV_X1    g395(.A(G1961), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n748), .A2(G19), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n563), .B2(new_n748), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(G1341), .Z(new_n825));
  NAND3_X1  g400(.A1(new_n817), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  NOR4_X1   g401(.A1(new_n763), .A2(new_n790), .A3(new_n815), .A4(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n748), .A2(G23), .ZN(new_n829));
  INV_X1    g404(.A(new_n598), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n748), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT33), .B(G1976), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G1971), .ZN(new_n834));
  NAND2_X1  g409(.A1(G166), .A2(G16), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G16), .B2(G22), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n833), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n748), .A2(G6), .ZN(new_n838));
  INV_X1    g413(.A(G305), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(new_n748), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT32), .B(G1981), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT88), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n840), .B(new_n842), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n837), .B(new_n843), .C1(new_n834), .C2(new_n836), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(KEYINPUT34), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(KEYINPUT34), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n748), .A2(G24), .ZN(new_n847));
  INV_X1    g422(.A(G290), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(new_n748), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT87), .B(G1986), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n849), .A2(new_n851), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n480), .A2(G131), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n482), .A2(G119), .ZN(new_n855));
  OR2_X1    g430(.A1(G95), .A2(G2105), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  MUX2_X1   g433(.A(G25), .B(new_n858), .S(G29), .Z(new_n859));
  XOR2_X1   g434(.A(KEYINPUT35), .B(G1991), .Z(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n859), .B(new_n861), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n852), .A2(new_n853), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n845), .A2(new_n846), .A3(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(KEYINPUT36), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(KEYINPUT36), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n828), .B1(new_n865), .B2(new_n866), .ZN(G311));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n864), .A2(KEYINPUT36), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n827), .B1(new_n868), .B2(new_n869), .ZN(G150));
  XNOR2_X1  g445(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n871));
  INV_X1    g446(.A(G559), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n635), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n635), .A2(new_n872), .A3(new_n871), .ZN(new_n875));
  INV_X1    g450(.A(G55), .ZN(new_n876));
  INV_X1    g451(.A(G93), .ZN(new_n877));
  OAI22_X1  g452(.A1(new_n876), .A2(new_n553), .B1(new_n523), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n547), .A2(G67), .A3(new_n548), .ZN(new_n880));
  NAND2_X1  g455(.A1(G80), .A2(G543), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G651), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n879), .A2(new_n883), .A3(KEYINPUT104), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n514), .B1(new_n880), .B2(new_n881), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n885), .B1(new_n886), .B2(new_n878), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n563), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n879), .A2(new_n883), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n889), .B(new_n885), .C1(new_n559), .C2(new_n562), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n874), .A2(new_n875), .A3(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n888), .A2(new_n890), .ZN(new_n893));
  INV_X1    g468(.A(new_n871), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n643), .A2(G559), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n895), .B2(new_n873), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT39), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT105), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n899), .B(KEYINPUT39), .C1(new_n892), .C2(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n891), .B1(new_n874), .B2(new_n875), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT39), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n895), .A2(new_n893), .A3(new_n873), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G860), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n889), .A2(G860), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT37), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(KEYINPUT106), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n907), .B1(new_n898), .B2(new_n900), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n915), .B2(new_n911), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(G145));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n661), .B(KEYINPUT107), .ZN(new_n919));
  INV_X1    g494(.A(G160), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n919), .A2(new_n920), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n486), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n923), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(G162), .A3(new_n921), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n652), .B(new_n858), .Z(new_n929));
  NAND2_X1  g504(.A1(new_n482), .A2(G130), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n930), .B(KEYINPUT108), .Z(new_n931));
  NAND2_X1  g506(.A1(new_n480), .A2(G142), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n464), .A2(G118), .ZN(new_n933));
  OAI21_X1  g508(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n931), .B(new_n932), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n929), .B(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(G164), .B1(new_n783), .B2(new_n784), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n777), .A2(new_n782), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT91), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n777), .A2(KEYINPUT91), .A3(new_n782), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n503), .A3(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n937), .A2(new_n942), .A3(new_n740), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n740), .B1(new_n937), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n806), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n783), .A2(new_n784), .A3(G164), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n503), .B1(new_n940), .B2(new_n941), .ZN(new_n947));
  OAI22_X1  g522(.A1(new_n946), .A2(new_n947), .B1(new_n733), .B2(new_n739), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n937), .A2(new_n942), .A3(new_n740), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n804), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n936), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n950), .A3(new_n936), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT109), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n945), .A2(new_n950), .A3(new_n936), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n953), .A2(KEYINPUT110), .A3(new_n955), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n928), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n927), .A2(new_n951), .ZN(new_n961));
  AOI21_X1  g536(.A(G37), .B1(new_n961), .B2(new_n956), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n918), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n959), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT110), .B1(new_n953), .B2(new_n955), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n965), .A2(new_n966), .A3(new_n951), .ZN(new_n967));
  OAI211_X1 g542(.A(KEYINPUT40), .B(new_n962), .C1(new_n967), .C2(new_n928), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n964), .A2(new_n968), .ZN(G395));
  NAND2_X1  g544(.A1(new_n889), .A2(new_n636), .ZN(new_n970));
  NAND2_X1  g545(.A1(G166), .A2(G305), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n839), .A2(G303), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(G290), .A2(new_n830), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n598), .A2(new_n617), .A3(new_n618), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n971), .A2(new_n972), .A3(new_n974), .A4(new_n975), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n977), .A2(KEYINPUT112), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT112), .B1(new_n977), .B2(new_n978), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT42), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n977), .A2(new_n978), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n647), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n647), .A2(new_n985), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n891), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n988), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(new_n893), .A3(new_n986), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n632), .A2(G299), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n627), .A2(new_n631), .B1(new_n574), .B2(new_n580), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT41), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT41), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n992), .B2(new_n993), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n989), .A2(new_n991), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n994), .B1(new_n989), .B2(new_n991), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n981), .B(new_n984), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n981), .A2(new_n984), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n893), .B1(new_n990), .B2(new_n986), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n987), .A2(new_n891), .A3(new_n988), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n999), .B(new_n1003), .C1(new_n1006), .C2(new_n994), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n970), .B1(new_n1008), .B2(new_n636), .ZN(G295));
  OAI21_X1  g584(.A(new_n970), .B1(new_n1008), .B2(new_n636), .ZN(G331));
  NAND2_X1  g585(.A1(new_n588), .A2(G168), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n584), .A2(new_n582), .B1(new_n531), .B2(new_n544), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n891), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1011), .A2(new_n890), .A3(new_n888), .A4(new_n1013), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1015), .A2(new_n994), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1012), .B1(new_n588), .B2(G168), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n893), .A2(new_n1018), .A3(KEYINPUT113), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n1014), .B2(new_n891), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1016), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n998), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1017), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n979), .A2(new_n980), .ZN(new_n1025));
  AOI21_X1  g600(.A(G37), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1015), .A2(new_n994), .A3(new_n1016), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT113), .B1(new_n893), .B2(new_n1018), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1014), .A2(new_n1020), .A3(new_n891), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1028), .A2(new_n1029), .B1(new_n893), .B2(new_n1018), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1027), .B1(new_n1030), .B2(new_n998), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n982), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n977), .A2(KEYINPUT112), .A3(new_n978), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT114), .B1(new_n979), .B2(new_n980), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1031), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT43), .B1(new_n1026), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1016), .A2(new_n994), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n998), .B1(new_n1016), .B2(new_n1015), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1037), .B(new_n1036), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G37), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1025), .B(new_n1027), .C1(new_n1030), .C2(new_n998), .ZN(new_n1045));
  AND4_X1   g620(.A1(KEYINPUT43), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT44), .B1(new_n1039), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT43), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1026), .B2(new_n1038), .ZN(new_n1050));
  AND4_X1   g625(.A1(new_n1049), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1052), .ZN(G397));
  INV_X1    g628(.A(G1384), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n489), .A2(new_n492), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n497), .A2(new_n501), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n482), .A2(G126), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1054), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT45), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n467), .A2(new_n470), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT68), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n475), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n467), .A2(KEYINPUT68), .A3(new_n470), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1064), .A2(new_n1065), .A3(G40), .A4(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1061), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1986), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(new_n848), .ZN(new_n1070));
  XOR2_X1   g645(.A(new_n1070), .B(KEYINPUT125), .Z(new_n1071));
  OR2_X1    g646(.A1(new_n1071), .A2(KEYINPUT48), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n785), .B(G2067), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n740), .B(G1996), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n858), .B(new_n860), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1068), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1077), .A2(KEYINPUT124), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(KEYINPUT124), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1071), .A2(KEYINPUT48), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1072), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n858), .A2(new_n861), .ZN(new_n1083));
  OAI22_X1  g658(.A1(new_n1082), .A2(new_n1083), .B1(G2067), .B2(new_n786), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1068), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1073), .A2(new_n740), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1068), .ZN(new_n1087));
  INV_X1    g662(.A(G1996), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1068), .A2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(KEYINPUT46), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT123), .B(KEYINPUT47), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1087), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1081), .A2(new_n1085), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT126), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1081), .A2(new_n1094), .A3(KEYINPUT126), .A4(new_n1085), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(G286), .A2(G8), .ZN(new_n1100));
  AOI21_X1  g675(.A(G1384), .B1(new_n493), .B2(new_n502), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT50), .ZN(new_n1102));
  OAI211_X1 g677(.A(G40), .B(G160), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g678(.A(KEYINPUT50), .B(G1384), .C1(new_n493), .C2(new_n502), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G2084), .ZN(new_n1106));
  AND4_X1   g681(.A1(G40), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1101), .A2(KEYINPUT45), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1061), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1966), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1105), .A2(new_n1106), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G8), .ZN(new_n1112));
  OAI211_X1 g687(.A(KEYINPUT51), .B(new_n1100), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1067), .B1(new_n1059), .B2(KEYINPUT50), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1106), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1114), .B(G8), .C1(new_n1119), .C2(G286), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1100), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g698(.A(KEYINPUT120), .B(new_n1100), .C1(new_n1115), .C2(new_n1118), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1113), .B(new_n1120), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT62), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1059), .A2(KEYINPUT50), .ZN(new_n1127));
  INV_X1    g702(.A(G2090), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n1107), .A4(new_n1117), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT115), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1116), .A2(new_n1131), .A3(new_n1128), .A4(new_n1117), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1109), .A2(new_n834), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(G303), .A2(G8), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT55), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(G8), .A3(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n595), .A2(G1976), .A3(new_n596), .A4(new_n597), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1139), .B(G8), .C1(new_n1059), .C2(new_n1067), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT116), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1107), .A2(new_n1101), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT116), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(G8), .A4(new_n1139), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(new_n1144), .A3(KEYINPUT52), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n1112), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT52), .ZN(new_n1148));
  INV_X1    g723(.A(G1976), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n599), .A2(new_n1149), .A3(new_n601), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .A4(new_n1139), .ZN(new_n1151));
  INV_X1    g726(.A(G1981), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n608), .A2(new_n612), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(G48), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n522), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1155));
  OAI22_X1  g730(.A1(new_n1154), .A2(new_n553), .B1(new_n1155), .B2(new_n514), .ZN(new_n1156));
  INV_X1    g731(.A(new_n604), .ZN(new_n1157));
  OAI21_X1  g732(.A(G1981), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT49), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1153), .A2(new_n1158), .A3(KEYINPUT49), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1161), .A2(new_n1147), .A3(new_n1162), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1145), .A2(new_n1151), .A3(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1135), .B(KEYINPUT55), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1105), .A2(new_n1128), .B1(new_n1109), .B2(new_n834), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1165), .B1(new_n1166), .B2(new_n1112), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1138), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT53), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n1109), .B2(G2078), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n821), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1169), .A2(G2078), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1061), .A2(new_n1107), .A3(new_n1108), .A4(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1171), .A2(KEYINPUT121), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT121), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1170), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n588), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1168), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT120), .B1(new_n1111), .B2(new_n1100), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1119), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1181), .A2(new_n1182), .A3(new_n1113), .A4(new_n1120), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1126), .A2(new_n1178), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1164), .A2(G168), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1137), .B1(new_n1134), .B2(G8), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT63), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1185), .A2(G168), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT63), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1112), .B1(new_n1133), .B2(new_n1129), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1190), .B1(new_n1191), .B2(new_n1137), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1138), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1163), .A2(new_n1149), .A3(new_n602), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1153), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1193), .A2(new_n1164), .B1(new_n1147), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1184), .A2(new_n1188), .A3(new_n1196), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1101), .A2(KEYINPUT45), .ZN(new_n1198));
  AOI211_X1 g773(.A(new_n1060), .B(G1384), .C1(new_n493), .C2(new_n502), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1172), .A2(G40), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1202));
  AOI211_X1 g777(.A(new_n475), .B(new_n1201), .C1(new_n1202), .C2(KEYINPUT122), .ZN(new_n1203));
  OAI211_X1 g778(.A(new_n1200), .B(new_n1203), .C1(KEYINPUT122), .C2(new_n1202), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1170), .A2(new_n1204), .A3(G301), .A4(new_n1171), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1170), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT121), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1171), .A2(KEYINPUT121), .A3(new_n1173), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1206), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1205), .B1(new_n1211), .B2(G301), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT54), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1170), .A2(new_n1204), .A3(new_n1171), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1213), .B1(new_n1215), .B2(G171), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1216), .B1(new_n588), .B2(new_n1176), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1168), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1214), .A2(new_n1217), .A3(new_n1125), .A4(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(G1956), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1220), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT57), .ZN(new_n1222));
  AND3_X1   g797(.A1(new_n574), .A2(new_n1222), .A3(new_n580), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1222), .B1(new_n574), .B2(new_n580), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g800(.A(KEYINPUT56), .B(G2072), .ZN(new_n1226));
  NAND4_X1  g801(.A1(new_n1061), .A2(new_n1107), .A3(new_n1108), .A4(new_n1226), .ZN(new_n1227));
  AND3_X1   g802(.A1(new_n1221), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1225), .B1(new_n1221), .B2(new_n1227), .ZN(new_n1229));
  OAI21_X1  g804(.A(KEYINPUT61), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g805(.A(new_n1225), .ZN(new_n1231));
  AND4_X1   g806(.A1(new_n1107), .A2(new_n1061), .A3(new_n1108), .A4(new_n1226), .ZN(new_n1232));
  AOI21_X1  g807(.A(G1956), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1231), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g809(.A(KEYINPUT61), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1221), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1230), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g813(.A(KEYINPUT117), .ZN(new_n1239));
  NAND4_X1  g814(.A1(new_n1200), .A2(new_n1239), .A3(new_n1088), .A4(new_n1107), .ZN(new_n1240));
  NAND4_X1  g815(.A1(new_n1061), .A2(new_n1088), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1241), .A2(KEYINPUT117), .ZN(new_n1242));
  XOR2_X1   g817(.A(KEYINPUT58), .B(G1341), .Z(new_n1243));
  NAND2_X1  g818(.A1(new_n1142), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g819(.A1(new_n1240), .A2(new_n1242), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1245), .A2(new_n563), .ZN(new_n1246));
  INV_X1    g821(.A(KEYINPUT118), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g824(.A(G1348), .ZN(new_n1250));
  OAI21_X1  g825(.A(new_n1250), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1251));
  INV_X1    g826(.A(G2067), .ZN(new_n1252));
  NAND2_X1  g827(.A1(new_n1146), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g828(.A1(new_n1251), .A2(KEYINPUT60), .A3(new_n1253), .ZN(new_n1254));
  AOI21_X1  g829(.A(KEYINPUT60), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1255));
  OAI21_X1  g830(.A(new_n1254), .B1(new_n1255), .B2(new_n632), .ZN(new_n1256));
  AND2_X1   g831(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1257));
  INV_X1    g832(.A(new_n632), .ZN(new_n1258));
  NAND3_X1  g833(.A1(new_n1257), .A2(KEYINPUT60), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g834(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  NAND4_X1  g835(.A1(new_n1245), .A2(new_n1247), .A3(KEYINPUT59), .A4(new_n563), .ZN(new_n1261));
  NAND4_X1  g836(.A1(new_n1238), .A2(new_n1249), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  NOR2_X1   g837(.A1(new_n1257), .A2(new_n632), .ZN(new_n1263));
  AOI21_X1  g838(.A(new_n1229), .B1(new_n1263), .B2(new_n1236), .ZN(new_n1264));
  AOI21_X1  g839(.A(KEYINPUT119), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g840(.A1(new_n1219), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g841(.A1(new_n1262), .A2(KEYINPUT119), .A3(new_n1264), .ZN(new_n1267));
  AOI21_X1  g842(.A(new_n1197), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g843(.A(new_n1076), .ZN(new_n1269));
  XNOR2_X1  g844(.A(G290), .B(new_n1069), .ZN(new_n1270));
  AOI211_X1 g845(.A(new_n1067), .B(new_n1061), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g846(.A(new_n1099), .B1(new_n1268), .B2(new_n1271), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g847(.A1(G319), .A2(new_n694), .ZN(new_n1274));
  AOI21_X1  g848(.A(new_n1274), .B1(new_n679), .B2(new_n681), .ZN(new_n1275));
  NAND3_X1  g849(.A1(new_n719), .A2(new_n721), .A3(new_n1275), .ZN(new_n1276));
  XNOR2_X1  g850(.A(new_n1276), .B(KEYINPUT127), .ZN(new_n1277));
  OAI21_X1  g851(.A(new_n1277), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1278));
  NOR2_X1   g852(.A1(new_n960), .A2(new_n963), .ZN(new_n1279));
  NOR2_X1   g853(.A1(new_n1278), .A2(new_n1279), .ZN(G308));
  OAI221_X1 g854(.A(new_n1277), .B1(new_n960), .B2(new_n963), .C1(new_n1050), .C2(new_n1051), .ZN(G225));
endmodule


