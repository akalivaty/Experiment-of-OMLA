//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n211), .B1(new_n212), .B2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G13), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n214), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI22_X1  g0022(.A1(new_n219), .A2(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(G87), .B2(G250), .ZN(new_n224));
  INV_X1    g0024(.A(G116), .ZN(new_n225));
  INV_X1    g0025(.A(G270), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(G50), .B2(G226), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  INV_X1    g0030(.A(G264), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n228), .B1(new_n201), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G238), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n202), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n212), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT1), .ZN(new_n236));
  NAND2_X1  g0036(.A1(G1), .A2(G13), .ZN(new_n237));
  INV_X1    g0037(.A(G20), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n206), .A2(new_n207), .ZN(new_n240));
  AOI211_X1 g0040(.A(new_n218), .B(new_n236), .C1(new_n239), .C2(new_n240), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G226), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G250), .B(G257), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G264), .B(G270), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G358));
  XOR2_X1   g0051(.A(G68), .B(G77), .Z(new_n252));
  XOR2_X1   g0052(.A(G50), .B(G58), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G107), .B(G116), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n237), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(G33), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n230), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n238), .A2(KEYINPUT23), .A3(G107), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n269), .A2(new_n271), .A3(new_n238), .A4(G87), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT22), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n267), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT23), .B1(new_n238), .B2(G107), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT90), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(KEYINPUT90), .B(KEYINPUT23), .C1(new_n238), .C2(G107), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G116), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT89), .ZN(new_n282));
  AND3_X1   g0082(.A1(new_n274), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT24), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT77), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(new_n268), .A3(G33), .ZN(new_n286));
  AOI21_X1  g0086(.A(KEYINPUT77), .B1(new_n270), .B2(KEYINPUT3), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n238), .A2(G87), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n289), .A2(new_n273), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n281), .A2(KEYINPUT89), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n283), .A2(new_n284), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n274), .A2(new_n293), .A3(new_n279), .A4(new_n282), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT24), .B1(new_n295), .B2(new_n291), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n266), .B1(new_n297), .B2(new_n260), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  OAI211_X1 g0099(.A(G1), .B(G13), .C1(new_n270), .C2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n285), .B1(new_n268), .B2(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n269), .ZN(new_n302));
  OR2_X1    g0102(.A1(G250), .A2(G1698), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n222), .A2(G1698), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n302), .A2(new_n286), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G294), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n300), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n299), .A2(KEYINPUT5), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT5), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G41), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n262), .A2(G45), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n300), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(new_n231), .ZN(new_n314));
  INV_X1    g0114(.A(G274), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(new_n308), .A3(new_n310), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n307), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G190), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(new_n319), .B2(G200), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n263), .A2(G107), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT25), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n298), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G179), .ZN(new_n329));
  NOR4_X1   g0129(.A1(new_n307), .A2(new_n314), .A3(new_n329), .A4(new_n318), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n298), .B2(new_n324), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT6), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n333), .A2(new_n221), .A3(G107), .ZN(new_n334));
  XNOR2_X1  g0134(.A(G97), .B(G107), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n238), .A2(new_n270), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n336), .A2(new_n238), .B1(new_n219), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT3), .B(G33), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(G20), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n269), .A2(new_n271), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT7), .A3(new_n238), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n230), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n260), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n265), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G97), .ZN(new_n347));
  INV_X1    g0147(.A(new_n263), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n221), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n345), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(G257), .B(new_n300), .C1(new_n311), .C2(new_n312), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT82), .B1(new_n351), .B2(new_n317), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(KEYINPUT82), .A3(new_n317), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT4), .ZN(new_n356));
  INV_X1    g0156(.A(G1698), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n356), .B1(new_n358), .B2(new_n220), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n269), .A2(new_n271), .A3(G250), .A4(G1698), .ZN(new_n360));
  AND2_X1   g0160(.A1(KEYINPUT4), .A2(G244), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n269), .A2(new_n271), .A3(new_n361), .A4(new_n357), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G33), .A2(G283), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n360), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n300), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(G200), .B1(new_n355), .B2(new_n365), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n351), .A2(KEYINPUT82), .A3(new_n317), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(new_n352), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n359), .A2(new_n364), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n237), .B1(G33), .B2(G41), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n368), .A2(new_n371), .A3(G190), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n350), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n327), .B1(new_n355), .B2(new_n365), .ZN(new_n374));
  XOR2_X1   g0174(.A(KEYINPUT71), .B(G179), .Z(new_n375));
  NAND3_X1  g0175(.A1(new_n368), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n345), .A2(new_n347), .A3(new_n349), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n326), .A2(new_n332), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n229), .A2(G1698), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n340), .B(new_n381), .C1(G226), .C2(G1698), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(KEYINPUT74), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT74), .B1(new_n382), .B2(new_n383), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n385), .A2(new_n386), .A3(new_n300), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(new_n315), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n300), .A2(new_n388), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n389), .B1(new_n391), .B2(G238), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT13), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT75), .ZN(new_n395));
  INV_X1    g0195(.A(new_n386), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(new_n370), .A3(new_n384), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT13), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n398), .A3(new_n392), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n394), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(KEYINPUT75), .B(KEYINPUT13), .C1(new_n387), .C2(new_n393), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(G169), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT14), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT14), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n400), .A2(new_n404), .A3(G169), .A4(new_n401), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n394), .A2(G179), .A3(new_n399), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n270), .A2(G20), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n219), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n337), .A2(new_n207), .B1(new_n238), .B2(G68), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n260), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  XOR2_X1   g0212(.A(KEYINPUT76), .B(KEYINPUT11), .Z(new_n413));
  XNOR2_X1  g0213(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n348), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT12), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n263), .B2(G68), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n262), .A2(G20), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n261), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n416), .B(new_n418), .C1(new_n420), .C2(new_n202), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n407), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT8), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G58), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n428), .A2(new_n337), .B1(new_n238), .B2(new_n219), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT15), .B(G87), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n409), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n260), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT73), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n263), .A2(G77), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n420), .A2(new_n219), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n340), .A2(G1698), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n437), .A2(new_n233), .B1(new_n230), .B2(new_n340), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n342), .A2(new_n229), .A3(G1698), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n370), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n389), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n391), .A2(G244), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n436), .B1(new_n375), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(G169), .B2(new_n443), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n424), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n426), .B(KEYINPUT70), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT69), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n427), .B(new_n448), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n263), .ZN(new_n451));
  INV_X1    g0251(.A(new_n450), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n420), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G159), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n337), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(G20), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n289), .A2(KEYINPUT78), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT78), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n302), .A2(new_n461), .A3(new_n286), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT7), .A2(G20), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(G20), .B1(new_n302), .B2(new_n286), .ZN(new_n465));
  OAI21_X1  g0265(.A(G68), .B1(new_n465), .B2(new_n339), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT79), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n289), .A2(new_n238), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n202), .B1(new_n468), .B2(KEYINPUT7), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT79), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n459), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n261), .B1(new_n473), .B2(KEYINPUT16), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT16), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n202), .B1(new_n341), .B2(new_n343), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n459), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n454), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G223), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n357), .ZN(new_n480));
  OR2_X1    g0280(.A1(new_n357), .A2(G226), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n302), .A2(new_n286), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G87), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n300), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n390), .A2(new_n229), .ZN(new_n485));
  NOR4_X1   g0285(.A1(new_n484), .A2(new_n375), .A3(new_n389), .A4(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT80), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n484), .A2(new_n389), .A3(new_n485), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n487), .B(new_n488), .C1(new_n327), .C2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(new_n327), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT80), .B1(new_n491), .B2(new_n486), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT18), .B1(new_n478), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT81), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n482), .A2(new_n483), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n389), .B1(new_n496), .B2(new_n370), .ZN(new_n497));
  INV_X1    g0297(.A(new_n485), .ZN(new_n498));
  AOI21_X1  g0298(.A(G200), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR4_X1   g0299(.A1(new_n484), .A2(G190), .A3(new_n389), .A4(new_n485), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n320), .A3(new_n498), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n502), .B(KEYINPUT81), .C1(G200), .C2(new_n489), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n471), .B1(new_n469), .B2(new_n470), .ZN(new_n506));
  OAI211_X1 g0306(.A(KEYINPUT16), .B(new_n458), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(new_n260), .A3(new_n477), .ZN(new_n508));
  INV_X1    g0308(.A(new_n454), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT17), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n504), .A2(new_n508), .A3(KEYINPUT17), .A4(new_n509), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n490), .A2(new_n492), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n508), .A2(new_n509), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT18), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n494), .A2(new_n512), .A3(new_n513), .A4(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n446), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n208), .A2(G20), .ZN(new_n520));
  INV_X1    g0320(.A(G150), .ZN(new_n521));
  OAI221_X1 g0321(.A(new_n520), .B1(new_n521), .B2(new_n337), .C1(new_n450), .C2(new_n409), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(new_n260), .B1(new_n207), .B2(new_n348), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n207), .B2(new_n420), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n340), .A2(G222), .A3(new_n357), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n525), .B(KEYINPUT68), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n437), .A2(new_n479), .B1(new_n219), .B2(new_n340), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n370), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n391), .A2(G226), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n441), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n375), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n524), .B(new_n532), .C1(G169), .C2(new_n531), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n524), .B(KEYINPUT9), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(G200), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n531), .A2(G190), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT10), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT10), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n535), .A2(new_n540), .A3(new_n536), .A4(new_n537), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n534), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(G200), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n443), .A2(G190), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n544), .A2(KEYINPUT72), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(KEYINPUT72), .ZN(new_n546));
  OAI221_X1 g0346(.A(new_n436), .B1(new_n543), .B2(new_n443), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n400), .A2(G200), .A3(new_n401), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n394), .A2(G190), .A3(new_n399), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n422), .A3(new_n549), .ZN(new_n550));
  AND4_X1   g0350(.A1(new_n519), .A2(new_n542), .A3(new_n547), .A4(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT19), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n408), .A2(new_n552), .A3(G97), .ZN(new_n553));
  NOR2_X1   g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  INV_X1    g0354(.A(G87), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n554), .A2(new_n555), .B1(new_n383), .B2(new_n238), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n553), .B1(new_n556), .B2(new_n552), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n238), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n202), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT83), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n557), .B(KEYINPUT83), .C1(new_n202), .C2(new_n558), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n260), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n430), .A2(new_n348), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n563), .B(new_n564), .C1(new_n265), .C2(new_n430), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n233), .A2(new_n357), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n220), .A2(G1698), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n302), .A2(new_n286), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n300), .B1(new_n568), .B2(new_n280), .ZN(new_n569));
  INV_X1    g0369(.A(new_n312), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n370), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G250), .ZN(new_n572));
  INV_X1    g0372(.A(new_n316), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n327), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n569), .A2(new_n574), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n375), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n565), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(G200), .B1(new_n569), .B2(new_n574), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n346), .A2(G87), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n563), .A2(new_n564), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT84), .ZN(new_n583));
  XNOR2_X1  g0383(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n576), .A2(G190), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n579), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT21), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n317), .B1(new_n313), .B2(new_n226), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n231), .A2(new_n357), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n286), .B(new_n589), .C1(new_n287), .C2(new_n288), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT85), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n302), .A2(G257), .A3(new_n357), .A4(new_n286), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT85), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n302), .A2(new_n593), .A3(new_n286), .A4(new_n589), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n342), .A2(G303), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n591), .A2(new_n592), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n370), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT86), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n596), .A2(KEYINPUT86), .A3(new_n370), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n588), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n346), .A2(G116), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n363), .B(new_n238), .C1(G33), .C2(new_n221), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n603), .B(new_n260), .C1(new_n238), .C2(G116), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT87), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT20), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n348), .A2(new_n225), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n602), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n604), .A2(new_n606), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT87), .B1(new_n604), .B2(new_n606), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(G169), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n587), .B1(new_n601), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n609), .A2(new_n612), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n601), .A2(G179), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n588), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n596), .A2(KEYINPUT86), .A3(new_n370), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT86), .B1(new_n596), .B2(new_n370), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n612), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n602), .A2(new_n607), .A3(new_n608), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n327), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n621), .A2(new_n624), .A3(KEYINPUT21), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n614), .A2(new_n617), .A3(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(G190), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n627), .B(new_n615), .C1(new_n601), .C2(new_n543), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT88), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n616), .B1(new_n621), .B2(G200), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT88), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(new_n627), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n626), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n380), .A2(new_n551), .A3(new_n586), .A4(new_n633), .ZN(G372));
  NAND2_X1  g0434(.A1(new_n626), .A2(KEYINPUT92), .ZN(new_n635));
  INV_X1    g0435(.A(new_n332), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT92), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n614), .A2(new_n617), .A3(new_n637), .A4(new_n625), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT93), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n373), .A2(new_n378), .ZN(new_n642));
  INV_X1    g0442(.A(new_n574), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT91), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n568), .A2(new_n280), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n370), .ZN(new_n646));
  AOI211_X1 g0446(.A(KEYINPUT91), .B(new_n300), .C1(new_n568), .C2(new_n280), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n327), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n565), .A2(new_n649), .A3(new_n577), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n563), .A2(new_n564), .A3(new_n581), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(G200), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n585), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n642), .A2(new_n325), .A3(new_n650), .A4(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n635), .A2(new_n636), .A3(KEYINPUT93), .A4(new_n638), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n641), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n374), .A2(new_n377), .A3(new_n376), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(new_n586), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n650), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n653), .A2(new_n650), .A3(new_n659), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(KEYINPUT26), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n551), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n512), .A2(new_n513), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n446), .A2(new_n667), .A3(new_n550), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n491), .A2(new_n486), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n508), .B2(new_n509), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n539), .A2(new_n541), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n534), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n666), .A2(new_n674), .ZN(G369));
  NAND2_X1  g0475(.A1(new_n635), .A2(new_n638), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n214), .A2(G20), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n262), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n615), .A2(new_n684), .ZN(new_n685));
  MUX2_X1   g0485(.A(new_n633), .B(new_n676), .S(new_n685), .Z(new_n686));
  NAND2_X1  g0486(.A1(new_n332), .A2(new_n683), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT94), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n298), .A2(new_n324), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n636), .B(new_n325), .C1(new_n689), .C2(new_n684), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n686), .A2(G330), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n636), .A2(new_n683), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n626), .A2(new_n684), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n691), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n692), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n216), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n554), .A2(new_n555), .A3(new_n225), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n699), .A2(new_n262), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n240), .B2(new_n699), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT28), .Z(new_n703));
  INV_X1    g0503(.A(G330), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n633), .A2(new_n380), .A3(new_n586), .A4(new_n684), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT31), .ZN(new_n706));
  OAI211_X1 g0506(.A(G179), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n307), .A2(new_n314), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n368), .A2(new_n576), .A3(new_n371), .A4(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT30), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  AND4_X1   g0510(.A1(new_n708), .A2(new_n368), .A3(new_n576), .A4(new_n371), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n601), .A2(new_n711), .A3(new_n712), .A4(G179), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n319), .B1(new_n371), .B2(new_n368), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n621), .A2(new_n715), .A3(new_n375), .A4(new_n648), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n714), .A2(KEYINPUT95), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT95), .B1(new_n714), .B2(new_n716), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n683), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n706), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n714), .A2(new_n716), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n704), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n665), .A2(new_n684), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT96), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT29), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n683), .B1(new_n657), .B2(new_n664), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT96), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n661), .B1(new_n662), .B2(KEYINPUT26), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n651), .A2(new_n583), .A3(new_n580), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n582), .A2(KEYINPUT84), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n585), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n658), .A3(new_n659), .A4(new_n578), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n626), .A2(new_n332), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n732), .B(new_n736), .C1(new_n737), .C2(new_n654), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(KEYINPUT29), .A3(new_n684), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n724), .B1(new_n731), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n703), .B1(new_n740), .B2(G1), .ZN(G364));
  XNOR2_X1  g0541(.A(KEYINPUT71), .B(G179), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n543), .A2(G190), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g0546(.A(KEYINPUT33), .B(G317), .Z(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n743), .A2(new_n320), .A3(new_n543), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G326), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n320), .A2(new_n543), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n238), .A2(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G303), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G190), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G329), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n745), .A2(new_n752), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n340), .B1(new_n761), .B2(G283), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n750), .A2(new_n755), .A3(new_n759), .A4(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n743), .A2(new_n320), .A3(G200), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n748), .B(new_n763), .C1(G322), .C2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G294), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n329), .A2(new_n543), .A3(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G311), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n744), .A2(new_n756), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(KEYINPUT97), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT97), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n744), .A2(new_n773), .A3(new_n756), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n765), .B1(new_n766), .B2(new_n769), .C1(new_n770), .C2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT98), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n769), .A2(new_n221), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n775), .A2(G77), .B1(G87), .B2(new_n754), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT32), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n757), .A2(new_n455), .ZN(new_n782));
  INV_X1    g0582(.A(new_n764), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n780), .B1(new_n781), .B2(new_n782), .C1(new_n201), .C2(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n779), .B(new_n784), .C1(new_n781), .C2(new_n782), .ZN(new_n785));
  INV_X1    g0585(.A(new_n746), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n342), .B1(new_n786), .B2(G68), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n785), .B(new_n787), .C1(new_n230), .C2(new_n760), .ZN(new_n788));
  INV_X1    g0588(.A(new_n749), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n207), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n778), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n791), .A2(KEYINPUT99), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(KEYINPUT99), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n237), .B1(G20), .B2(new_n327), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G13), .A2(G33), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(G20), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n794), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n698), .A2(new_n342), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G355), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n254), .A2(G45), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n460), .A2(new_n462), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n698), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n206), .A2(G45), .A3(new_n207), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n802), .B1(G116), .B2(new_n216), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n796), .B1(new_n800), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n262), .B1(new_n677), .B2(G45), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n699), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n799), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n809), .B(new_n812), .C1(new_n686), .C2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n686), .A2(G330), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n686), .A2(G330), .ZN(new_n816));
  INV_X1    g0616(.A(new_n812), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n814), .B1(new_n815), .B2(new_n818), .ZN(G396));
  INV_X1    g0619(.A(KEYINPUT101), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n436), .B2(new_n684), .ZN(new_n821));
  OR3_X1    g0621(.A1(new_n436), .A2(new_n820), .A3(new_n684), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n547), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n445), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n445), .A2(new_n683), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n727), .A2(new_n730), .A3(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n683), .B(new_n826), .C1(new_n657), .C2(new_n664), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n724), .A2(KEYINPUT102), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n724), .A2(KEYINPUT102), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n827), .A2(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n827), .A2(new_n828), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n831), .B(new_n817), .C1(new_n832), .C2(new_n829), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n794), .A2(new_n797), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n826), .A2(new_n797), .B1(new_n219), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT100), .B(G143), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n786), .A2(G150), .B1(new_n764), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n837), .B1(new_n838), .B2(new_n789), .C1(new_n776), .C2(new_n455), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT34), .Z(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G58), .B2(new_n768), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n761), .A2(G68), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G50), .A2(new_n754), .B1(new_n758), .B2(G132), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n841), .A2(new_n804), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n760), .A2(new_n555), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n783), .A2(new_n766), .B1(new_n770), .B2(new_n757), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(new_n775), .C2(G116), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n754), .A2(G107), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n779), .B1(new_n786), .B2(G283), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n340), .B1(new_n749), .B2(G303), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n847), .A2(new_n848), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n844), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n835), .B(new_n812), .C1(new_n852), .C2(new_n795), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n833), .A2(new_n853), .ZN(G384));
  INV_X1    g0654(.A(KEYINPUT40), .ZN(new_n855));
  INV_X1    g0655(.A(new_n681), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n474), .B1(KEYINPUT16), .B2(new_n473), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n509), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n518), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n857), .A2(new_n509), .B1(new_n669), .B2(new_n681), .ZN(new_n860));
  INV_X1    g0660(.A(new_n510), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT37), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n514), .A2(new_n515), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n515), .A2(new_n856), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n510), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT38), .B1(new_n859), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n424), .A2(new_n683), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n423), .A2(new_n683), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n407), .A2(new_n423), .B1(new_n550), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n826), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n705), .A2(KEYINPUT31), .B1(new_n719), .B2(new_n683), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n855), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n826), .B1(new_n721), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n864), .B1(new_n671), .B2(new_n667), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n864), .A2(new_n865), .A3(new_n510), .ZN(new_n884));
  INV_X1    g0684(.A(new_n670), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(new_n864), .A3(new_n510), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n884), .A2(new_n863), .B1(new_n886), .B2(KEYINPUT37), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n882), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n867), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n881), .A2(new_n890), .A3(KEYINPUT40), .A4(new_n874), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n721), .A2(new_n880), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n879), .A2(new_n891), .A3(new_n551), .A4(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n879), .A2(G330), .A3(new_n891), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n551), .A2(G330), .A3(new_n892), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n893), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT103), .Z(new_n898));
  NAND3_X1  g0698(.A1(new_n731), .A2(new_n551), .A3(new_n739), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n674), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n898), .B(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n890), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n859), .A2(new_n867), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n882), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n903), .A2(new_n871), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n889), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n445), .A2(new_n683), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n908), .B(new_n874), .C1(new_n828), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n671), .A2(new_n856), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n907), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n901), .B(new_n913), .Z(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n262), .B2(new_n677), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT35), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n238), .B(new_n237), .C1(new_n336), .C2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n917), .B(G116), .C1(new_n916), .C2(new_n336), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT36), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n240), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(G50), .B2(new_n202), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(G1), .A3(new_n214), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n915), .A2(new_n919), .A3(new_n922), .ZN(G367));
  NOR2_X1   g0723(.A1(new_n760), .A2(new_n219), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n342), .B(new_n924), .C1(new_n786), .C2(G159), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n925), .B1(new_n201), .B2(new_n753), .C1(new_n838), .C2(new_n757), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n776), .A2(new_n207), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n768), .A2(G68), .ZN(new_n928));
  INV_X1    g0728(.A(new_n836), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n928), .B1(new_n789), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n783), .A2(new_n521), .ZN(new_n931));
  NOR4_X1   g0731(.A1(new_n926), .A2(new_n927), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT46), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n753), .B2(new_n225), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n754), .A2(KEYINPUT46), .A3(G116), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n934), .B(new_n935), .C1(new_n746), .C2(new_n766), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT110), .ZN(new_n937));
  XNOR2_X1  g0737(.A(KEYINPUT111), .B(G317), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n758), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(G303), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n783), .A2(new_n940), .B1(new_n230), .B2(new_n769), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n775), .B2(G283), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n937), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n804), .B(new_n943), .C1(G97), .C2(new_n761), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n749), .A2(G311), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n932), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT47), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n794), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n651), .A2(new_n684), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT104), .Z(new_n950));
  NAND2_X1  g0750(.A1(new_n653), .A2(new_n650), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n661), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(new_n799), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n805), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n800), .B1(new_n216), .B2(new_n430), .C1(new_n955), .C2(new_n250), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n948), .A2(new_n812), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n810), .B(KEYINPUT109), .Z(new_n958));
  INV_X1    g0758(.A(KEYINPUT45), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT107), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n659), .A2(new_n683), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT105), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n642), .B1(new_n350), .B2(new_n684), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n696), .A2(new_n960), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n960), .B1(new_n696), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n959), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n696), .A2(new_n968), .A3(new_n964), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n968), .B1(new_n696), .B2(new_n964), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n691), .A2(new_n695), .ZN(new_n972));
  INV_X1    g0772(.A(new_n693), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n964), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT107), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n696), .A2(new_n960), .A3(new_n964), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n967), .A2(new_n971), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n692), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n967), .A2(new_n971), .A3(new_n692), .A4(new_n977), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n816), .A2(new_n691), .A3(new_n694), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n691), .B1(new_n816), .B2(new_n694), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT108), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(KEYINPUT108), .B2(new_n692), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n740), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n740), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n699), .B(KEYINPUT41), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n958), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n964), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n972), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT42), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n659), .B1(new_n964), .B2(new_n332), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT106), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n993), .B1(new_n683), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n952), .A2(new_n953), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n999), .B1(new_n996), .B2(new_n1000), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n1002), .A2(new_n1003), .B1(new_n692), .B2(new_n991), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1003), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n692), .A2(new_n991), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1005), .A2(new_n1006), .A3(new_n1001), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n957), .B1(new_n990), .B2(new_n1008), .ZN(G387));
  AOI22_X1  g0809(.A1(new_n775), .A2(G303), .B1(new_n764), .B2(new_n938), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n770), .B2(new_n746), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G322), .B2(new_n749), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT48), .Z(new_n1013));
  INV_X1    g0813(.A(G283), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(new_n1014), .B2(new_n769), .C1(new_n766), .C2(new_n753), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(G326), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n760), .A2(new_n225), .B1(new_n757), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n1017), .A2(new_n804), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n804), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n783), .A2(new_n207), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n450), .A2(new_n746), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n769), .A2(new_n430), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n760), .A2(new_n221), .B1(new_n757), .B2(new_n521), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n219), .B2(new_n753), .C1(new_n455), .C2(new_n789), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1021), .B(new_n1027), .C1(G68), .C2(new_n775), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT112), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n794), .B1(new_n1020), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n955), .B1(new_n247), .B2(G45), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n700), .B2(new_n801), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n700), .ZN(new_n1033));
  AOI21_X1  g0833(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n428), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n207), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1033), .B(new_n1034), .C1(new_n1036), .C2(KEYINPUT50), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(KEYINPUT50), .B2(new_n1036), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n1032), .A2(new_n1038), .B1(G107), .B2(new_n216), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n817), .B1(new_n1039), .B2(new_n800), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1030), .B(new_n1040), .C1(new_n691), .C2(new_n813), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n986), .A2(new_n958), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n987), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n699), .B1(new_n740), .B2(new_n986), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1041), .B(new_n1042), .C1(new_n1043), .C2(new_n1044), .ZN(G393));
  NAND3_X1  g0845(.A1(new_n1043), .A2(new_n980), .A3(new_n981), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n982), .A2(new_n987), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n1047), .A3(new_n699), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n980), .A2(new_n981), .A3(new_n958), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n800), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n216), .A2(new_n221), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n805), .C2(new_n257), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n769), .A2(new_n225), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G311), .A2(new_n764), .B1(new_n749), .B2(G317), .ZN(new_n1054));
  XOR2_X1   g0854(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1055));
  XOR2_X1   g0855(.A(new_n1054), .B(new_n1055), .Z(new_n1056));
  OAI221_X1 g0856(.A(new_n342), .B1(new_n940), .B2(new_n746), .C1(new_n776), .C2(new_n766), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n753), .A2(new_n1014), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G322), .B2(new_n758), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n230), .B2(new_n760), .ZN(new_n1060));
  OR4_X1    g0860(.A1(new_n1053), .A2(new_n1056), .A3(new_n1057), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G150), .A2(new_n749), .B1(new_n764), .B2(G159), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT51), .Z(new_n1063));
  NAND2_X1  g0863(.A1(new_n786), .A2(G50), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n769), .A2(new_n219), .B1(new_n929), .B2(new_n757), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n775), .B2(new_n1035), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1063), .A2(new_n804), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n753), .A2(new_n202), .B1(new_n760), .B2(new_n555), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1061), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1052), .B1(new_n1069), .B2(new_n794), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n812), .C1(new_n813), .C2(new_n964), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1049), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1048), .A2(new_n1072), .ZN(G390));
  NAND3_X1  g0873(.A1(new_n724), .A2(new_n875), .A3(new_n874), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n824), .A2(new_n738), .A3(new_n684), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n825), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n874), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n871), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n890), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n665), .A2(new_n684), .A3(new_n875), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n825), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n871), .B1(new_n1082), .B2(new_n874), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT39), .B1(new_n888), .B2(new_n889), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(KEYINPUT39), .B2(new_n870), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1074), .B(new_n1080), .C1(new_n1083), .C2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n909), .B1(new_n729), .B2(new_n875), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n874), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1078), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n903), .A2(new_n906), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1079), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n881), .A2(G330), .A3(new_n874), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1086), .B(new_n958), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1090), .A2(new_n797), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n776), .A2(new_n221), .B1(new_n225), .B2(new_n783), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G283), .B2(new_n749), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n754), .A2(G87), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n786), .A2(G107), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n842), .B1(new_n766), .B2(new_n757), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n340), .B(new_n1099), .C1(G77), .C2(new_n768), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n760), .A2(new_n207), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n754), .A2(G150), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT53), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT54), .B(G143), .Z(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n775), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n764), .A2(G132), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n786), .A2(G137), .ZN(new_n1108));
  INV_X1    g0908(.A(G125), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n340), .B1(new_n757), .B2(new_n1109), .C1(new_n769), .C2(new_n455), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G128), .B2(new_n749), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1101), .B1(new_n1102), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n794), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n450), .A2(new_n834), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1094), .A2(new_n812), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1093), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(KEYINPUT116), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT116), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1093), .A2(new_n1119), .A3(new_n1116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n723), .ZN(new_n1122));
  OAI211_X1 g0922(.A(G330), .B(new_n875), .C1(new_n876), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1088), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1092), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n1082), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1076), .ZN(new_n1127));
  OAI211_X1 g0927(.A(G330), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1088), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1074), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1131), .A2(new_n674), .A3(new_n899), .A4(new_n895), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1086), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n899), .A2(new_n674), .A3(new_n895), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1080), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1092), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1138), .A3(new_n1086), .A4(new_n1131), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1134), .A2(new_n1139), .A3(new_n699), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT115), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT115), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1134), .A2(new_n1139), .A3(new_n1142), .A4(new_n699), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1121), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(G378));
  NAND2_X1  g0945(.A1(new_n834), .A2(new_n207), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n1147));
  NAND2_X1  g0947(.A1(new_n524), .A2(new_n856), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n542), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n542), .A2(new_n1148), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1147), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n673), .A2(new_n533), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1148), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1147), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(new_n1149), .A3(new_n1157), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1152), .A2(new_n1153), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1153), .B1(new_n1152), .B2(new_n1158), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n812), .B(new_n1146), .C1(new_n1161), .C2(new_n798), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n761), .A2(G58), .B1(new_n758), .B2(G283), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n219), .B2(new_n753), .C1(new_n776), .C2(new_n430), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1021), .A2(new_n299), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n928), .B1(new_n789), .B2(new_n225), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1166), .A2(KEYINPUT117), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1166), .A2(KEYINPUT117), .ZN(new_n1168));
  NOR4_X1   g0968(.A1(new_n1164), .A2(new_n1165), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n221), .B2(new_n746), .C1(new_n230), .C2(new_n783), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT58), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1165), .B(new_n207), .C1(G33), .C2(G41), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n786), .A2(G132), .B1(G128), .B2(new_n764), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n754), .A2(new_n1105), .B1(G150), .B2(new_n768), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n1109), .C2(new_n789), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G137), .B2(new_n775), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT59), .Z(new_n1177));
  AOI22_X1  g0977(.A1(new_n761), .A2(G159), .B1(new_n758), .B2(G124), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1178), .A2(new_n270), .A3(new_n299), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1172), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n795), .B1(new_n1171), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1162), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n894), .A2(new_n913), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n879), .A2(G330), .A3(new_n891), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1185), .A2(new_n910), .A3(new_n912), .A4(new_n907), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1184), .A2(new_n1186), .A3(new_n1161), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1161), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1183), .B1(new_n1189), .B2(new_n958), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1161), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1184), .A2(new_n1186), .A3(new_n1161), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(KEYINPUT57), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n899), .A2(new_n674), .A3(new_n895), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1092), .B1(new_n1197), .B2(new_n1080), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1123), .A2(new_n1088), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1199), .B(new_n1079), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1196), .B1(new_n1201), .B2(new_n1131), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n699), .B1(new_n1195), .B2(new_n1202), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1074), .A2(new_n1129), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1204), .A2(new_n1127), .B1(new_n1125), .B2(new_n1082), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1135), .B1(new_n1133), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT57), .B1(new_n1189), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1190), .B1(new_n1203), .B2(new_n1207), .ZN(G375));
  AOI22_X1  g1008(.A1(new_n775), .A2(G150), .B1(G50), .B2(new_n768), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT122), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n786), .A2(new_n1105), .B1(G137), .B2(new_n764), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1021), .B1(G58), .B2(new_n761), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT123), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1213), .B2(new_n1212), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n749), .A2(G132), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G159), .A2(new_n754), .B1(new_n758), .B2(G128), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1210), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n775), .A2(G107), .B1(G116), .B2(new_n786), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1219), .A2(KEYINPUT120), .ZN(new_n1220));
  OAI221_X1 g1020(.A(KEYINPUT120), .B1(new_n225), .B2(new_n746), .C1(new_n776), .C2(new_n230), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n766), .C2(new_n789), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT121), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1222), .B(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1024), .B(new_n1224), .C1(G303), .C2(new_n758), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n754), .A2(G97), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n764), .A2(G283), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1225), .A2(new_n342), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1218), .B1(new_n1228), .B2(new_n924), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n794), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1088), .A2(new_n797), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n834), .A2(new_n202), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1230), .A2(new_n812), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n958), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1236));
  OAI21_X1  g1036(.A(KEYINPUT124), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT124), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1238), .B(new_n1233), .C1(new_n1205), .C2(new_n1235), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1196), .A2(new_n1205), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1132), .A2(new_n1241), .A3(new_n989), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(G381));
  INV_X1    g1044(.A(G375), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1117), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1140), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(G390), .ZN(new_n1250));
  OR2_X1    g1050(.A1(G393), .A2(G396), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(G387), .A2(G384), .A3(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1249), .A2(new_n1250), .A3(new_n1243), .A4(new_n1252), .ZN(G407));
  OAI211_X1 g1053(.A(G407), .B(G213), .C1(G343), .C2(new_n1248), .ZN(G409));
  NAND2_X1  g1054(.A1(G387), .A2(new_n1250), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G390), .B(new_n957), .C1(new_n990), .C2(new_n1008), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT127), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G393), .A2(G396), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1251), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1251), .A2(new_n1258), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1256), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1255), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1189), .A2(new_n989), .A3(new_n1206), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n1269), .A2(new_n1235), .B1(new_n1162), .B2(new_n1182), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1247), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(G375), .B2(new_n1144), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT126), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n833), .A2(new_n1273), .A3(new_n853), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1196), .A2(new_n1205), .A3(KEYINPUT60), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1132), .A3(new_n699), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT60), .B1(new_n1196), .B2(new_n1205), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1240), .B(new_n1274), .C1(new_n1276), .C2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1277), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1282), .A2(new_n699), .A3(new_n1132), .A4(new_n1275), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1283), .A2(new_n1240), .A3(new_n1279), .A4(new_n1274), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n682), .A2(G213), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1272), .A2(new_n1285), .A3(KEYINPUT63), .A4(new_n1286), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1266), .A2(new_n1267), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1272), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1271), .B(KEYINPUT125), .C1(G375), .C2(new_n1144), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1286), .A3(new_n1292), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n682), .A2(G213), .A3(G2897), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1281), .A2(new_n1284), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1281), .B2(new_n1284), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1289), .B1(new_n1293), .B2(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1291), .A2(new_n1285), .A3(new_n1286), .A4(new_n1292), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1288), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1256), .B2(new_n1261), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1264), .B1(new_n1303), .B2(new_n1255), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1299), .A2(KEYINPUT62), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1272), .A2(new_n1286), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT61), .B1(new_n1306), .B2(new_n1297), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1272), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1304), .B1(new_n1305), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1301), .A2(new_n1311), .ZN(G405));
  NOR2_X1   g1112(.A1(G375), .A2(new_n1144), .ZN(new_n1313));
  AND2_X1   g1113(.A1(G375), .A2(new_n1247), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1304), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1313), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1266), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1315), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1285), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1315), .A2(new_n1317), .A3(new_n1281), .A4(new_n1284), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(G402));
endmodule


