//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n540, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n464), .A2(new_n466), .A3(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n474));
  INV_X1    g049(.A(G100), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(new_n462), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT68), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n478), .A2(new_n462), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n477), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT69), .Z(G162));
  NAND3_X1  g061(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n463), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G102), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n462), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n478), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n490), .A2(new_n492), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n507), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n504), .A2(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n502), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  XOR2_X1   g091(.A(KEYINPUT70), .B(G51), .Z(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(G543), .A3(new_n503), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n499), .A2(new_n503), .A3(G89), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n518), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n499), .A2(G63), .ZN(new_n524));
  NAND3_X1  g099(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n501), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G168));
  NAND3_X1  g102(.A1(new_n503), .A2(G52), .A3(G543), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n499), .A2(new_n503), .A3(G90), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n528), .B(new_n529), .C1(new_n530), .C2(new_n501), .ZN(G301));
  INV_X1    g106(.A(G301), .ZN(G171));
  NAND3_X1  g107(.A1(new_n503), .A2(G43), .A3(G543), .ZN(new_n533));
  INV_X1    g108(.A(G81), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  OAI221_X1 g110(.A(new_n533), .B1(new_n534), .B2(new_n512), .C1(new_n535), .C2(new_n501), .ZN(new_n536));
  INV_X1    g111(.A(G860), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT71), .ZN(G153));
  AND3_X1   g114(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G36), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n540), .A2(new_n543), .ZN(G188));
  NAND2_X1  g119(.A1(G78), .A2(G543), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n507), .A2(new_n509), .ZN(new_n546));
  INV_X1    g121(.A(G65), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n512), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n548), .A2(G651), .B1(new_n549), .B2(G91), .ZN(new_n550));
  OAI211_X1 g125(.A(G53), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(new_n552), .ZN(G299));
  INV_X1    g128(.A(G168), .ZN(G286));
  INV_X1    g129(.A(new_n504), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G49), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n549), .A2(G87), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n499), .B2(G74), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(G288));
  NAND2_X1  g134(.A1(G73), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G61), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n546), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n562), .A2(KEYINPUT72), .A3(G651), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n565), .A2(new_n566), .B1(G86), .B2(new_n549), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n555), .A2(G48), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(G305));
  INV_X1    g144(.A(G85), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n512), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n501), .ZN(new_n573));
  AOI211_X1 g148(.A(new_n571), .B(new_n573), .C1(G47), .C2(new_n555), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G301), .A2(G868), .ZN(new_n576));
  NAND2_X1  g151(.A1(G79), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G66), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n546), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n503), .A2(G54), .A3(G543), .ZN(new_n581));
  INV_X1    g156(.A(G92), .ZN(new_n582));
  OAI21_X1  g157(.A(KEYINPUT10), .B1(new_n512), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT10), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n499), .A2(new_n503), .A3(new_n584), .A4(G92), .ZN(new_n585));
  AND4_X1   g160(.A1(new_n580), .A2(new_n581), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(KEYINPUT73), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(KEYINPUT73), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n576), .B1(new_n590), .B2(G868), .ZN(G284));
  OAI21_X1  g166(.A(new_n576), .B1(new_n590), .B2(G868), .ZN(G321));
  NAND2_X1  g167(.A1(G286), .A2(G868), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT9), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n551), .B(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n499), .A2(new_n503), .A3(G91), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n499), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n501), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT74), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G868), .ZN(G297));
  OAI21_X1  g176(.A(new_n593), .B1(new_n600), .B2(G868), .ZN(G280));
  AOI21_X1  g177(.A(new_n589), .B1(G559), .B2(new_n537), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT75), .ZN(G148));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n590), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n535), .A2(new_n501), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n533), .B1(new_n534), .B2(new_n512), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n607), .B1(G868), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g187(.A1(G123), .A2(new_n480), .B1(new_n483), .B2(G135), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(KEYINPUT77), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(KEYINPUT77), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n615), .B(new_n616), .C1(G111), .C2(new_n462), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND2_X1  g194(.A1(new_n478), .A2(new_n491), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT76), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n623), .A2(G2100), .ZN(new_n624));
  AND2_X1   g199(.A1(new_n623), .A2(G2100), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n619), .B(new_n626), .C1(new_n622), .C2(new_n624), .ZN(G156));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  XOR2_X1   g204(.A(G2427), .B(G2430), .Z(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(KEYINPUT78), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n629), .A2(new_n631), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(KEYINPUT78), .ZN(new_n636));
  NAND4_X1  g211(.A1(new_n632), .A2(new_n634), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT16), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(KEYINPUT79), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n642), .A2(new_n644), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n642), .A2(KEYINPUT79), .A3(new_n644), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n646), .A2(new_n647), .A3(G14), .A4(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT17), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  XNOR2_X1  g229(.A(G2084), .B(G2090), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT80), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT81), .Z(new_n658));
  INV_X1    g233(.A(new_n654), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n659), .A3(new_n651), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT18), .Z(new_n661));
  AOI21_X1  g236(.A(new_n656), .B1(new_n659), .B2(new_n652), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n659), .B2(new_n651), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n658), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2096), .B(G2100), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n669), .A2(KEYINPUT82), .ZN(new_n670));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(KEYINPUT82), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n667), .A2(new_n668), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(new_n672), .B2(new_n669), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n672), .A2(KEYINPUT83), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1986), .B(G1996), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  INV_X1    g258(.A(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1991), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n682), .B(new_n686), .ZN(G229));
  NOR2_X1   g262(.A1(G25), .A2(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n480), .A2(G119), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n483), .A2(G131), .ZN(new_n690));
  NOR2_X1   g265(.A1(G95), .A2(G2105), .ZN(new_n691));
  OAI21_X1  g266(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n689), .B(new_n690), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT84), .Z(new_n694));
  AOI21_X1  g269(.A(new_n688), .B1(new_n694), .B2(G29), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT35), .B(G1991), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT85), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G23), .B(G288), .S(G16), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT33), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1976), .ZN(new_n701));
  MUX2_X1   g276(.A(G6), .B(G305), .S(G16), .Z(new_n702));
  XOR2_X1   g277(.A(KEYINPUT32), .B(G1981), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G22), .B(G303), .S(G16), .Z(new_n705));
  XOR2_X1   g280(.A(KEYINPUT87), .B(G1971), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n701), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n698), .B1(new_n708), .B2(KEYINPUT34), .ZN(new_n709));
  MUX2_X1   g284(.A(G24), .B(G290), .S(G16), .Z(new_n710));
  XOR2_X1   g285(.A(KEYINPUT86), .B(G1986), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n709), .B(new_n712), .C1(KEYINPUT34), .C2(new_n708), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT36), .ZN(new_n714));
  NOR2_X1   g289(.A1(G29), .A2(G35), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G162), .B2(G29), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT29), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G2090), .Z(new_n718));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(G27), .ZN(new_n721));
  AOI211_X1 g296(.A(new_n719), .B(new_n721), .C1(new_n497), .C2(G29), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n719), .B2(new_n721), .ZN(new_n723));
  INV_X1    g298(.A(G2078), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G19), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(G16), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n536), .B2(G16), .ZN(new_n728));
  MUX2_X1   g303(.A(new_n727), .B(new_n728), .S(KEYINPUT88), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1341), .ZN(new_n730));
  OR2_X1    g305(.A1(KEYINPUT24), .A2(G34), .ZN(new_n731));
  NAND2_X1  g306(.A1(KEYINPUT24), .A2(G34), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n731), .A2(new_n720), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G160), .B2(new_n720), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(G2084), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT91), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n725), .A2(new_n730), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT28), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n720), .A2(G26), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n480), .A2(G128), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n483), .A2(G140), .ZN(new_n741));
  NOR2_X1   g316(.A1(G104), .A2(G2105), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n740), .B(new_n741), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AOI211_X1 g319(.A(new_n738), .B(new_n739), .C1(new_n744), .C2(G29), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n738), .B2(new_n739), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT89), .B(G2067), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n746), .B(new_n747), .Z(new_n748));
  NOR2_X1   g323(.A1(G29), .A2(G32), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n480), .A2(G129), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n483), .A2(G141), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n491), .A2(G105), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT26), .Z(new_n754));
  NAND4_X1  g329(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n749), .B1(new_n756), .B2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT27), .B(G1996), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT31), .B(G11), .ZN(new_n760));
  NOR2_X1   g335(.A1(G16), .A2(G21), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G168), .B2(G16), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G1966), .ZN(new_n763));
  INV_X1    g338(.A(G28), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n764), .B2(KEYINPUT30), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(KEYINPUT30), .B2(new_n764), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n618), .B2(new_n720), .ZN(new_n767));
  NOR2_X1   g342(.A1(G5), .A2(G16), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G171), .B2(G16), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n767), .B1(new_n769), .B2(G1961), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n759), .A2(new_n760), .A3(new_n763), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n483), .A2(G139), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT25), .Z(new_n774));
  AOI22_X1  g349(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n772), .B(new_n774), .C1(new_n462), .C2(new_n775), .ZN(new_n776));
  MUX2_X1   g351(.A(G33), .B(new_n776), .S(G29), .Z(new_n777));
  AOI22_X1  g352(.A1(new_n777), .A2(G2072), .B1(G2084), .B2(new_n734), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G2072), .B2(new_n777), .ZN(new_n779));
  NOR4_X1   g354(.A1(new_n737), .A2(new_n748), .A3(new_n771), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G1961), .B2(new_n769), .ZN(new_n781));
  INV_X1    g356(.A(G4), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G16), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n589), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1348), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n762), .A2(G1966), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT90), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n784), .A2(new_n785), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G20), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(G16), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G299), .B2(G16), .ZN(new_n793));
  MUX2_X1   g368(.A(new_n792), .B(new_n793), .S(KEYINPUT23), .Z(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT93), .B(G1956), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n781), .A2(new_n790), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n714), .A2(new_n718), .A3(new_n797), .ZN(G150));
  INV_X1    g373(.A(G150), .ZN(G311));
  OAI211_X1 g374(.A(G55), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n800));
  INV_X1    g375(.A(G93), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n512), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n507), .A2(new_n509), .A3(G67), .ZN(new_n803));
  NAND2_X1  g378(.A1(G80), .A2(G543), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n501), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n537), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT37), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n589), .A2(new_n605), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT95), .B1(new_n802), .B2(new_n805), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n813), .A2(new_n536), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n610), .A2(new_n812), .A3(new_n806), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n811), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  AOI21_X1  g396(.A(G860), .B1(new_n821), .B2(KEYINPUT96), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(KEYINPUT96), .B2(new_n821), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n808), .B1(new_n823), .B2(new_n824), .ZN(G145));
  XOR2_X1   g400(.A(new_n618), .B(G160), .Z(new_n826));
  XNOR2_X1  g401(.A(G162), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT97), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n776), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n744), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n755), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n497), .ZN(new_n832));
  INV_X1    g407(.A(G142), .ZN(new_n833));
  NOR2_X1   g408(.A1(G106), .A2(G2105), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n482), .A2(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G130), .B2(new_n480), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n621), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n693), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n827), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n831), .B(G164), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n839), .ZN(new_n843));
  AOI21_X1  g418(.A(G37), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n832), .B1(KEYINPUT98), .B2(new_n839), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n842), .A2(new_n846), .A3(new_n840), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n827), .A2(KEYINPUT99), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n827), .A2(KEYINPUT99), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n845), .A2(new_n847), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g427(.A(new_n606), .B(new_n818), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT41), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n580), .A2(new_n581), .A3(new_n583), .A4(new_n585), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n599), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n599), .A2(new_n855), .A3(KEYINPUT100), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(new_n586), .B2(G299), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n854), .B(new_n856), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT100), .B1(new_n599), .B2(new_n855), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n586), .A2(G299), .A3(new_n858), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n864), .B1(new_n862), .B2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n856), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n861), .B1(new_n867), .B2(KEYINPUT41), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n853), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n856), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT101), .B1(new_n857), .B2(new_n859), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n869), .B1(new_n873), .B2(new_n853), .ZN(new_n874));
  NOR2_X1   g449(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n874), .B(new_n875), .Z(new_n876));
  XNOR2_X1  g451(.A(G303), .B(G288), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(G290), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(G290), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(G305), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n878), .A2(new_n568), .A3(new_n567), .A4(new_n879), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(KEYINPUT102), .B2(KEYINPUT42), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n876), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(G868), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(G868), .B2(new_n806), .ZN(G295));
  OAI21_X1  g462(.A(new_n886), .B1(G868), .B2(new_n806), .ZN(G331));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n860), .B1(new_n873), .B2(new_n854), .ZN(new_n890));
  INV_X1    g465(.A(new_n523), .ZN(new_n891));
  INV_X1    g466(.A(new_n526), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(G301), .A3(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n530), .A2(new_n501), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n529), .A2(new_n528), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n894), .B(new_n896), .C1(new_n526), .C2(new_n523), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n817), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n893), .A2(new_n897), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n816), .A3(new_n815), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(KEYINPUT104), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n818), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n890), .A2(KEYINPUT105), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n902), .A2(new_n904), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(new_n868), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n867), .A2(new_n901), .A3(new_n899), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n910), .A2(KEYINPUT106), .A3(new_n883), .A4(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT105), .B1(new_n890), .B2(new_n905), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n868), .A2(new_n907), .A3(new_n908), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n914), .A2(new_n915), .A3(new_n883), .A4(new_n911), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n873), .A2(new_n854), .B1(new_n901), .B2(new_n899), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n870), .B1(new_n862), .B2(new_n863), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n919), .B1(new_n854), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n873), .B2(new_n908), .ZN(new_n922));
  INV_X1    g497(.A(new_n883), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n912), .A2(new_n913), .A3(new_n918), .A4(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n889), .B1(new_n925), .B2(KEYINPUT43), .ZN(new_n926));
  XNOR2_X1  g501(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n916), .B(KEYINPUT106), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n910), .A2(new_n911), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n923), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n913), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n926), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n928), .A2(new_n913), .A3(new_n927), .A4(new_n930), .ZN(new_n933));
  INV_X1    g508(.A(new_n927), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n925), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n935), .A3(new_n889), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n936), .A2(KEYINPUT107), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(KEYINPUT107), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(G397));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  OR3_X1    g515(.A1(G290), .A2(new_n940), .A3(G1986), .ZN(new_n941));
  XOR2_X1   g516(.A(KEYINPUT108), .B(G1384), .Z(new_n942));
  AOI21_X1  g517(.A(KEYINPUT45), .B1(new_n497), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G40), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n469), .A2(new_n472), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n940), .B1(G290), .B2(G1986), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n941), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(G1986), .A3(G290), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT110), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n744), .B(G2067), .Z(new_n953));
  NAND2_X1  g528(.A1(new_n755), .A2(G1996), .ZN(new_n954));
  INV_X1    g529(.A(G1996), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n756), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n693), .B(new_n696), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n947), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n952), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G288), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(G1976), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  INV_X1    g539(.A(new_n488), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(new_n478), .B2(G126), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n492), .B1(new_n966), .B2(new_n462), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n495), .A2(new_n496), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n470), .A2(new_n471), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n462), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n467), .A2(new_n468), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n971), .B(G40), .C1(new_n462), .C2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n963), .B(G8), .C1(new_n969), .C2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n945), .A2(new_n497), .A3(new_n964), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n963), .B1(new_n976), .B2(G8), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n962), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n979), .A2(KEYINPUT112), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1976), .ZN(new_n983));
  NAND3_X1  g558(.A1(G288), .A2(new_n979), .A3(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n962), .B(new_n980), .C1(new_n975), .C2(new_n977), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n969), .A2(KEYINPUT50), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n497), .A2(new_n988), .A3(new_n964), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n945), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(G2090), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n973), .B1(new_n969), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n994));
  AOI21_X1  g569(.A(G1971), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(G8), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(G303), .A2(G8), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n997), .B(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n975), .A2(new_n977), .ZN(new_n1002));
  NAND2_X1  g577(.A1(G305), .A2(G1981), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n567), .A2(new_n684), .A3(new_n568), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT49), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1005), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1002), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n986), .A2(new_n1001), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n993), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1966), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n990), .A2(G2084), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1013), .A2(KEYINPUT114), .A3(new_n1014), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(G8), .A3(G168), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n999), .B(G8), .C1(new_n991), .C2(new_n995), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT63), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n986), .A2(new_n1008), .A3(new_n1001), .A4(KEYINPUT115), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1011), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT63), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n986), .A2(new_n1008), .A3(new_n1001), .A4(new_n1022), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1028), .B2(new_n1021), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1008), .A2(new_n983), .A3(new_n961), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n1004), .B(KEYINPUT113), .Z(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n986), .A2(new_n1008), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1022), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1033), .A2(new_n1002), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT116), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1030), .A2(new_n1039), .A3(new_n1036), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n1020), .B2(G286), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1043), .B1(new_n1020), .B2(G286), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1042), .A2(KEYINPUT51), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT121), .B1(new_n1013), .B2(G2078), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n993), .A2(new_n1049), .A3(new_n724), .A4(new_n1012), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(KEYINPUT53), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n990), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1961), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n987), .A2(KEYINPUT118), .A3(new_n945), .A4(new_n989), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1057));
  NAND2_X1  g632(.A1(new_n993), .A2(new_n994), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(G2078), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1051), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G171), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT123), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(new_n1063), .A3(G171), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT62), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1028), .B1(new_n1047), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1065), .A2(new_n1068), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1956), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n990), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n993), .A2(new_n994), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT57), .B1(new_n550), .B2(KEYINPUT117), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1076), .B(new_n599), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1077), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1072), .A2(new_n1079), .A3(new_n1074), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1053), .A2(new_n785), .A3(new_n1055), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n976), .A2(G2067), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n590), .A2(KEYINPUT60), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1081), .A2(KEYINPUT61), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT119), .B(G1996), .Z(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1058), .B2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT58), .B(G1341), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n976), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1088), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n993), .A2(KEYINPUT120), .A3(new_n994), .A4(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n610), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT59), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(new_n1097), .A3(new_n610), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT61), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n590), .A2(KEYINPUT60), .ZN(new_n1103));
  OR3_X1    g678(.A1(new_n1084), .A2(new_n1085), .A3(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1086), .A2(new_n1099), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1084), .A2(new_n590), .A3(new_n1080), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1106), .A2(new_n1078), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n943), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1109), .A2(new_n724), .A3(new_n945), .A4(new_n994), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1056), .A2(new_n1059), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(G171), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(KEYINPUT54), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1062), .A2(new_n1064), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1060), .A2(G301), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1115), .B(KEYINPUT54), .C1(G301), .C2(new_n1111), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1105), .A2(new_n1107), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1067), .B1(new_n1070), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n960), .B1(new_n1041), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n946), .B1(new_n953), .B2(new_n756), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n947), .A2(KEYINPUT46), .A3(new_n955), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT46), .B1(new_n947), .B2(new_n955), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n1123), .B(KEYINPUT47), .Z(new_n1124));
  INV_X1    g699(.A(new_n696), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n694), .A2(new_n1125), .ZN(new_n1126));
  OAI22_X1  g701(.A1(new_n957), .A2(new_n1126), .B1(G2067), .B2(new_n744), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n947), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT48), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n949), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n959), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n959), .A2(new_n1131), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n949), .A2(new_n1129), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1124), .B(new_n1128), .C1(new_n1130), .C2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT125), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT126), .B1(new_n1119), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1137), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1069), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1143), .A2(new_n1067), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1139), .B(new_n1140), .C1(new_n1144), .C2(new_n960), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1138), .A2(new_n1145), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g721(.A1(G229), .A2(G227), .ZN(new_n1148));
  AOI21_X1  g722(.A(new_n1148), .B1(new_n844), .B2(new_n850), .ZN(new_n1149));
  AND2_X1   g723(.A1(new_n649), .A2(G319), .ZN(new_n1150));
  NAND4_X1  g724(.A1(new_n933), .A2(new_n935), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n1152));
  XNOR2_X1  g726(.A(new_n1151), .B(new_n1152), .ZN(G308));
  XNOR2_X1  g727(.A(new_n1151), .B(KEYINPUT127), .ZN(G225));
endmodule


