//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT67), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT69), .Z(new_n208));
  NOR3_X1   g007(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n209), .B1(G169gat), .B2(G176gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n208), .A2(new_n210), .B1(G183gat), .B2(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT72), .ZN(new_n213));
  XNOR2_X1  g012(.A(G127gat), .B(G134gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT70), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G127gat), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT70), .B1(new_n217), .B2(G134gat), .ZN(new_n218));
  INV_X1    g017(.A(G120gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G113gat), .ZN(new_n220));
  INV_X1    g019(.A(G113gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G120gat), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI22_X1  g022(.A1(new_n216), .A2(new_n218), .B1(KEYINPUT1), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT71), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT1), .B1(new_n220), .B2(new_n222), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n214), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G134gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G127gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n217), .A2(G134gat), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT70), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n218), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n226), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n226), .A2(new_n214), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT71), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n213), .B1(new_n228), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239));
  INV_X1    g038(.A(G169gat), .ZN(new_n240));
  INV_X1    g039(.A(G176gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(KEYINPUT23), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT23), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(G169gat), .B2(G176gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G183gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(new_n203), .A3(KEYINPUT64), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(G183gat), .B2(G190gat), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT24), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT24), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(G183gat), .A3(G190gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n246), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT65), .B1(new_n257), .B2(KEYINPUT25), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n247), .A2(KEYINPUT24), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n261), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n252), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n248), .A2(new_n250), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n259), .B(new_n260), .C1(new_n264), .C2(new_n246), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n256), .A2(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT25), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n239), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n271), .ZN(new_n273));
  AOI211_X1 g072(.A(KEYINPUT66), .B(new_n273), .C1(new_n258), .C2(new_n265), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n212), .B(new_n238), .C1(new_n272), .C2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G227gat), .A2(G233gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n212), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n256), .A2(new_n250), .A3(new_n248), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n270), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n259), .B1(new_n279), .B2(new_n260), .ZN(new_n280));
  AOI211_X1 g079(.A(KEYINPUT65), .B(KEYINPUT25), .C1(new_n278), .C2(new_n270), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n271), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT66), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n239), .A3(new_n271), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n277), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n228), .A2(new_n236), .A3(new_n213), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n238), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n275), .B(new_n276), .C1(new_n285), .C2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT34), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT32), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n275), .B1(new_n285), .B2(new_n287), .ZN(new_n291));
  INV_X1    g090(.A(new_n276), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT33), .B1(new_n291), .B2(new_n292), .ZN(new_n294));
  XOR2_X1   g093(.A(G15gat), .B(G43gat), .Z(new_n295));
  XNOR2_X1  g094(.A(G71gat), .B(G99gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n293), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  AOI221_X4 g098(.A(new_n290), .B1(KEYINPUT33), .B2(new_n297), .C1(new_n291), .C2(new_n292), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n289), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g102(.A(KEYINPUT73), .B(new_n289), .C1(new_n299), .C2(new_n300), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n294), .A2(new_n298), .ZN(new_n305));
  INV_X1    g104(.A(new_n293), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n289), .ZN(new_n308));
  INV_X1    g107(.A(new_n300), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G228gat), .A2(G233gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n311), .B(KEYINPUT82), .Z(new_n312));
  INV_X1    g111(.A(G148gat), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT76), .B1(new_n313), .B2(G141gat), .ZN(new_n314));
  INV_X1    g113(.A(G141gat), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT77), .B1(new_n315), .B2(G148gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(new_n315), .A3(G148gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(new_n313), .A3(G141gat), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n314), .A2(new_n316), .A3(new_n318), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  OR2_X1    g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(KEYINPUT2), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n313), .A2(G141gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n315), .A2(G148gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(new_n322), .A3(new_n323), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  XNOR2_X1  g131(.A(G197gat), .B(G204gat), .ZN(new_n333));
  INV_X1    g132(.A(G211gat), .ZN(new_n334));
  INV_X1    g133(.A(G218gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n333), .B1(KEYINPUT22), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT83), .ZN(new_n338));
  XOR2_X1   g137(.A(G211gat), .B(G218gat), .Z(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n337), .A2(new_n339), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n339), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n332), .B(new_n340), .C1(new_n343), .C2(new_n338), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n331), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n345), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n343), .B1(new_n347), .B2(new_n332), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n312), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G22gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n311), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT29), .B1(new_n331), .B2(new_n345), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT3), .B1(new_n343), .B2(new_n332), .ZN(new_n353));
  OAI221_X1 g152(.A(new_n351), .B1(new_n352), .B2(new_n343), .C1(new_n331), .C2(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n349), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n350), .B1(new_n349), .B2(new_n354), .ZN(new_n356));
  OAI21_X1  g155(.A(G78gat), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n354), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G22gat), .ZN(new_n359));
  INV_X1    g158(.A(G78gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n349), .A2(new_n350), .A3(new_n354), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT31), .B(G50gat), .ZN(new_n363));
  INV_X1    g162(.A(G106gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n357), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n357), .B2(new_n362), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n303), .A2(new_n304), .A3(new_n310), .A4(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G1gat), .B(G29gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT0), .ZN(new_n371));
  XNOR2_X1  g170(.A(G57gat), .B(G85gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n371), .B(new_n372), .Z(new_n373));
  NAND2_X1  g172(.A1(new_n325), .A2(new_n330), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n374), .A2(KEYINPUT3), .B1(new_n224), .B2(new_n227), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n347), .ZN(new_n376));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT5), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n228), .A2(new_n236), .A3(new_n331), .ZN(new_n382));
  XOR2_X1   g181(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n224), .A2(new_n227), .A3(new_n325), .A4(new_n330), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n385), .A2(KEYINPUT79), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n382), .A2(new_n390), .A3(new_n384), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n381), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(G127gat), .B(G134gat), .Z(new_n393));
  AOI21_X1  g192(.A(new_n218), .B1(new_n393), .B2(KEYINPUT70), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n227), .B1(new_n394), .B2(new_n226), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n374), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n387), .A3(KEYINPUT80), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n374), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n379), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n228), .A2(new_n236), .A3(new_n331), .A4(new_n383), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n387), .A2(KEYINPUT4), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n401), .A2(new_n402), .B1(new_n347), .B2(new_n375), .ZN(new_n403));
  OAI22_X1  g202(.A1(new_n377), .A2(new_n400), .B1(new_n403), .B2(KEYINPUT5), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n373), .B1(new_n392), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT81), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n385), .A2(KEYINPUT79), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n388), .A2(new_n386), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n391), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(new_n376), .A3(new_n380), .ZN(new_n412));
  INV_X1    g211(.A(new_n400), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n401), .A2(new_n402), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n376), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n413), .A2(new_n378), .B1(new_n415), .B2(new_n379), .ZN(new_n416));
  INV_X1    g215(.A(new_n373), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n407), .B1(new_n408), .B2(new_n418), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n392), .A2(new_n404), .A3(new_n373), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT81), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(KEYINPUT6), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n343), .ZN(new_n425));
  AND2_X1   g224(.A1(G226gat), .A2(G233gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n282), .A2(new_n212), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(KEYINPUT29), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n425), .B(new_n427), .C1(new_n285), .C2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G8gat), .B(G36gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT74), .ZN(new_n432));
  XNOR2_X1  g231(.A(G64gat), .B(G92gat), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n432), .B(new_n433), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n282), .A2(new_n212), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n285), .A2(new_n426), .B1(new_n428), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n430), .B(new_n435), .C1(new_n437), .C2(new_n425), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT75), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT30), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT30), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n438), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n430), .B1(new_n437), .B2(new_n425), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n434), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n424), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT35), .B1(new_n369), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n310), .A2(new_n301), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n357), .A2(new_n362), .ZN(new_n451));
  INV_X1    g250(.A(new_n365), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n357), .A2(new_n362), .A3(new_n365), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT84), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n446), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n441), .A2(KEYINPUT84), .A3(new_n443), .A4(new_n445), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n418), .A2(new_n405), .A3(new_n406), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT35), .B1(new_n461), .B2(new_n423), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n456), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n449), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n403), .A2(new_n377), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT39), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n378), .B1(new_n397), .B2(new_n399), .ZN(new_n467));
  OR3_X1    g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n417), .B1(new_n465), .B2(new_n466), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT85), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT40), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n418), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n471), .B2(new_n470), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n459), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n461), .A2(new_n423), .A3(new_n438), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n444), .A2(KEYINPUT37), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT37), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n430), .B(new_n477), .C1(new_n437), .C2(new_n425), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n434), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n475), .B1(KEYINPUT38), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n481));
  INV_X1    g280(.A(new_n427), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n212), .B1(new_n272), .B2(new_n274), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n482), .B1(new_n483), .B2(new_n428), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n481), .B1(new_n484), .B2(new_n425), .ZN(new_n485));
  INV_X1    g284(.A(new_n437), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n485), .B1(new_n343), .B2(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n484), .A2(new_n481), .A3(new_n425), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT37), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n478), .A2(new_n434), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(KEYINPUT38), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n455), .B1(new_n480), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n304), .A2(new_n310), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n307), .A2(new_n309), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT73), .B1(new_n496), .B2(new_n289), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT36), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n450), .A2(KEYINPUT36), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n448), .A2(new_n455), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n494), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n464), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G15gat), .B(G22gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G1gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n506), .A2(KEYINPUT16), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(new_n505), .ZN(new_n509));
  INV_X1    g308(.A(G8gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G43gat), .B(G50gat), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n512), .A2(KEYINPUT15), .ZN(new_n513));
  XOR2_X1   g312(.A(KEYINPUT90), .B(G29gat), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G36gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(G29gat), .A2(G36gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT14), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n513), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n513), .A2(new_n517), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n522), .B(new_n515), .C1(KEYINPUT15), .C2(new_n512), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT17), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n521), .A2(new_n523), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n509), .B(G8gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n526), .ZN(new_n531));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n529), .A2(new_n531), .A3(KEYINPUT18), .A4(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n532), .A3(new_n531), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT18), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n509), .A2(G8gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n509), .A2(G8gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n524), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n531), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n532), .B(KEYINPUT13), .Z(new_n541));
  AOI21_X1  g340(.A(KEYINPUT92), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n543));
  INV_X1    g342(.A(new_n541), .ZN(new_n544));
  AOI211_X1 g343(.A(new_n543), .B(new_n544), .C1(new_n531), .C2(new_n539), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n533), .B(new_n536), .C1(new_n542), .C2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT88), .ZN(new_n548));
  XOR2_X1   g347(.A(G113gat), .B(G141gat), .Z(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G169gat), .B(G197gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT12), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n546), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n539), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n524), .B1(new_n537), .B2(new_n538), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n541), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n543), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n540), .A2(KEYINPUT92), .A3(new_n541), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n561), .A2(new_n553), .A3(new_n533), .A4(new_n536), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT93), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n555), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n546), .A2(KEYINPUT93), .A3(new_n554), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G85gat), .A2(G92gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT7), .ZN(new_n569));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  INV_X1    g369(.A(G85gat), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G99gat), .B(G106gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT96), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n569), .A2(new_n573), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n579), .A2(new_n575), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n575), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n525), .A2(new_n528), .A3(new_n577), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n577), .ZN(new_n584));
  AND2_X1   g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n584), .A2(new_n526), .B1(KEYINPUT41), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G190gat), .B(G218gat), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n585), .A2(KEYINPUT41), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT95), .ZN(new_n591));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n588), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n583), .A2(new_n594), .A3(new_n586), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n589), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n593), .B1(new_n589), .B2(new_n595), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT97), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n601));
  INV_X1    g400(.A(G155gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(G57gat), .B(G64gat), .ZN(new_n608));
  XOR2_X1   g407(.A(G71gat), .B(G78gat), .Z(new_n609));
  INV_X1    g408(.A(KEYINPUT94), .ZN(new_n610));
  AOI211_X1 g409(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n610), .B2(new_n609), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n608), .A2(new_n607), .ZN(new_n613));
  OR3_X1    g412(.A1(new_n613), .A2(new_n610), .A3(new_n609), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n612), .A2(new_n614), .ZN(new_n619));
  OAI211_X1 g418(.A(G231gat), .B(G233gat), .C1(new_n619), .C2(KEYINPUT21), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n620), .A3(new_n217), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n615), .A2(new_n616), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n530), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n217), .B1(new_n618), .B2(new_n620), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n511), .B1(new_n616), .B2(new_n615), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n618), .A2(new_n620), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(G127gat), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n627), .B1(new_n629), .B2(new_n621), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n606), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n624), .B1(new_n622), .B2(new_n625), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(new_n627), .A3(new_n621), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(new_n633), .A3(new_n605), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n599), .A2(new_n600), .A3(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n631), .A2(new_n634), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n597), .A2(new_n598), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT97), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n579), .B(new_n575), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n619), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n576), .A2(new_n612), .A3(new_n614), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n612), .B2(new_n614), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n643), .A2(new_n644), .B1(new_n584), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT98), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n643), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n648), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n584), .A2(new_n645), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT10), .B1(new_n641), .B2(new_n642), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n655), .B(new_n647), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n649), .A2(new_n651), .A3(new_n654), .A4(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n654), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n646), .A2(new_n648), .ZN(new_n661));
  INV_X1    g460(.A(new_n651), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n636), .A2(new_n639), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT99), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n636), .A2(new_n639), .A3(KEYINPUT99), .A4(new_n665), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n502), .A2(new_n567), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n424), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(new_n506), .ZN(G1324gat));
  NOR2_X1   g471(.A1(new_n670), .A2(new_n460), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(new_n510), .B2(new_n673), .ZN(new_n676));
  MUX2_X1   g475(.A(new_n675), .B(new_n676), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g476(.A(G15gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n670), .B2(new_n450), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT100), .Z(new_n680));
  AND2_X1   g479(.A1(new_n498), .A2(new_n499), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n670), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(new_n682), .ZN(G1326gat));
  NOR2_X1   g482(.A1(new_n670), .A2(new_n368), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT43), .B(G22gat), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  NAND2_X1  g485(.A1(new_n502), .A2(new_n638), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(KEYINPUT101), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n599), .B1(new_n464), .B2(new_n501), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n566), .A2(new_n635), .A3(new_n664), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n514), .B1(new_n695), .B2(new_n424), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n690), .A2(new_n694), .ZN(new_n697));
  INV_X1    g496(.A(new_n424), .ZN(new_n698));
  INV_X1    g497(.A(new_n514), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT102), .ZN(G1328gat));
  INV_X1    g502(.A(G36gat), .ZN(new_n704));
  INV_X1    g503(.A(new_n460), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n697), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT46), .Z(new_n707));
  OAI21_X1  g506(.A(G36gat), .B1(new_n695), .B2(new_n460), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1329gat));
  INV_X1    g508(.A(new_n681), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n689), .A2(new_n710), .A3(new_n692), .A4(new_n694), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G43gat), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n450), .A2(G43gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n713), .B1(new_n712), .B2(new_n715), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n712), .A2(KEYINPUT103), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(KEYINPUT47), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OAI22_X1  g520(.A1(new_n716), .A2(new_n717), .B1(new_n719), .B2(KEYINPUT47), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1330gat));
  OAI21_X1  g522(.A(G50gat), .B1(new_n695), .B2(new_n368), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT48), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(G50gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n697), .A2(new_n727), .A3(new_n455), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n724), .B(new_n728), .C1(new_n725), .C2(KEYINPUT48), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1331gat));
  NAND3_X1  g531(.A1(new_n566), .A2(new_n639), .A3(new_n636), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n665), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n502), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n698), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g537(.A1(new_n735), .A2(new_n460), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  NAND3_X1  g542(.A1(new_n736), .A2(G71gat), .A3(new_n710), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT106), .B1(new_n735), .B2(new_n450), .ZN(new_n745));
  INV_X1    g544(.A(G71gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n735), .A2(KEYINPUT106), .A3(new_n450), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n744), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n368), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT107), .B(G78gat), .Z(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1335gat));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n754), .B1(new_n566), .B2(new_n637), .ZN(new_n755));
  AOI211_X1 g554(.A(KEYINPUT108), .B(new_n635), .C1(new_n564), .C2(new_n565), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n665), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n693), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n424), .ZN(new_n760));
  INV_X1    g559(.A(new_n757), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT51), .B1(new_n690), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT110), .Z(new_n763));
  NAND4_X1  g562(.A1(new_n502), .A2(KEYINPUT51), .A3(new_n638), .A4(new_n761), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n690), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n761), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n698), .A2(new_n571), .A3(new_n664), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n760), .B1(new_n768), .B2(new_n769), .ZN(G1336gat));
  OAI21_X1  g569(.A(G92gat), .B1(new_n759), .B2(new_n460), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n705), .A2(new_n572), .A3(new_n664), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n771), .B(new_n772), .C1(new_n768), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n771), .B1(new_n775), .B2(new_n773), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT52), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n759), .B2(new_n681), .ZN(new_n779));
  OR3_X1    g578(.A1(new_n450), .A2(G99gat), .A3(new_n665), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n768), .B2(new_n780), .ZN(G1338gat));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n689), .A2(new_n455), .A3(new_n692), .A4(new_n758), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G106gat), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n368), .A2(G106gat), .A3(new_n665), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n782), .B(new_n784), .C1(new_n768), .C2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n762), .ZN(new_n788));
  AOI211_X1 g587(.A(new_n599), .B(new_n757), .C1(new_n464), .C2(new_n501), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT109), .B1(new_n789), .B2(KEYINPUT51), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n764), .A2(new_n765), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n793), .A3(new_n785), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT111), .B1(new_n775), .B2(new_n786), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n784), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n796), .A2(new_n797), .A3(KEYINPUT53), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n797), .B1(new_n796), .B2(KEYINPUT53), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n787), .B1(new_n798), .B2(new_n799), .ZN(G1339gat));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n646), .B2(new_n648), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n649), .A2(new_n802), .A3(new_n658), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n654), .B1(new_n661), .B2(new_n801), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT55), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n659), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT113), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n808), .A3(new_n659), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n803), .A2(new_n804), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n807), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n540), .A2(new_n541), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n532), .B1(new_n529), .B2(new_n531), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n552), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n562), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n813), .A2(new_n599), .A3(new_n817), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n813), .A2(new_n566), .B1(new_n665), .B2(new_n817), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n599), .B2(new_n819), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n820), .A2(new_n635), .B1(new_n664), .B2(new_n733), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n705), .A2(new_n424), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n369), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n567), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n456), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(new_n221), .A3(new_n566), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n826), .A2(new_n828), .ZN(G1340gat));
  AOI21_X1  g628(.A(G120gat), .B1(new_n825), .B2(new_n664), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n827), .A2(new_n219), .A3(new_n665), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(G1341gat));
  NAND3_X1  g631(.A1(new_n825), .A2(new_n217), .A3(new_n635), .ZN(new_n833));
  OAI21_X1  g632(.A(G127gat), .B1(new_n827), .B2(new_n637), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1342gat));
  NAND3_X1  g634(.A1(new_n825), .A2(new_n229), .A3(new_n638), .ZN(new_n836));
  XNOR2_X1  g635(.A(KEYINPUT114), .B(KEYINPUT56), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  OAI21_X1  g638(.A(G134gat), .B1(new_n827), .B2(new_n599), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(G1343gat));
  NAND2_X1  g640(.A1(new_n681), .A2(new_n822), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n821), .A2(new_n455), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n806), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n564), .A2(new_n565), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n810), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT115), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n811), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n849), .A2(new_n853), .A3(new_n811), .A4(new_n850), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n847), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n817), .A2(new_n665), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n599), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n818), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n635), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n733), .A2(new_n664), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n455), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT57), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n567), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n863), .A2(KEYINPUT117), .A3(G141gat), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT117), .B1(new_n863), .B2(G141gat), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n710), .A2(new_n368), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n823), .A2(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n867), .A2(G141gat), .A3(new_n566), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n868), .A2(KEYINPUT58), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n863), .A2(G141gat), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT118), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT118), .B1(new_n871), .B2(new_n872), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n869), .A2(new_n870), .B1(new_n873), .B2(new_n874), .ZN(G1344gat));
  INV_X1    g674(.A(new_n867), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n313), .A3(new_n664), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n845), .A2(new_n862), .ZN(new_n878));
  AOI211_X1 g677(.A(KEYINPUT59), .B(new_n313), .C1(new_n878), .C2(new_n664), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n819), .A2(new_n599), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n635), .B1(new_n881), .B2(new_n858), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT57), .B(new_n455), .C1(new_n882), .C2(new_n860), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT119), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n668), .A2(new_n566), .A3(new_n669), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n852), .A2(new_n854), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n564), .A2(new_n565), .A3(new_n846), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n856), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n858), .B1(new_n888), .B2(new_n638), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n885), .B1(new_n889), .B2(new_n637), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n844), .B1(new_n890), .B2(new_n368), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n821), .A2(new_n892), .A3(KEYINPUT57), .A4(new_n455), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n884), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n894), .A2(new_n681), .A3(new_n664), .A4(new_n822), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n880), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n877), .B1(new_n879), .B2(new_n896), .ZN(G1345gat));
  NAND3_X1  g696(.A1(new_n876), .A2(new_n602), .A3(new_n635), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n878), .A2(new_n635), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n602), .ZN(G1346gat));
  NOR3_X1   g699(.A1(new_n867), .A2(G162gat), .A3(new_n599), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT120), .Z(new_n902));
  NAND2_X1  g701(.A1(new_n878), .A2(new_n638), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G162gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1347gat));
  NOR2_X1   g704(.A1(new_n460), .A2(new_n698), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n821), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(new_n824), .ZN(new_n908));
  AOI21_X1  g707(.A(G169gat), .B1(new_n908), .B2(new_n567), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n456), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n910), .A2(new_n240), .A3(new_n566), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n909), .A2(new_n911), .ZN(G1348gat));
  NOR3_X1   g711(.A1(new_n910), .A2(new_n241), .A3(new_n665), .ZN(new_n913));
  XOR2_X1   g712(.A(new_n913), .B(KEYINPUT122), .Z(new_n914));
  AOI21_X1  g713(.A(G176gat), .B1(new_n908), .B2(new_n664), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(G1349gat));
  NAND3_X1  g718(.A1(new_n908), .A2(new_n202), .A3(new_n635), .ZN(new_n920));
  OAI21_X1  g719(.A(G183gat), .B1(new_n910), .B2(new_n637), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g721(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(G1350gat));
  OAI21_X1  g723(.A(G190gat), .B1(new_n910), .B2(new_n599), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT61), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n908), .A2(new_n203), .A3(new_n638), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1351gat));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n884), .A2(new_n891), .A3(new_n929), .A4(new_n893), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n681), .A2(new_n906), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n455), .B1(new_n859), .B2(new_n885), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n933), .A2(new_n844), .B1(new_n883), .B2(KEYINPUT119), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n929), .B1(new_n934), .B2(new_n893), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n567), .A2(G197gat), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n932), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n843), .A2(new_n931), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(G197gat), .B1(new_n939), .B2(new_n567), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n937), .A2(new_n940), .ZN(G1352gat));
  NAND2_X1  g740(.A1(new_n894), .A2(KEYINPUT124), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n942), .A2(new_n664), .A3(new_n931), .A4(new_n930), .ZN(new_n943));
  XOR2_X1   g742(.A(KEYINPUT125), .B(G204gat), .Z(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  AND4_X1   g745(.A1(new_n664), .A2(new_n843), .A3(new_n931), .A4(new_n944), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT126), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n946), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1353gat));
  AND2_X1   g752(.A1(new_n931), .A2(new_n635), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n334), .B1(new_n894), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT63), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n334), .A3(new_n635), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1354gat));
  OAI21_X1  g757(.A(KEYINPUT127), .B1(new_n932), .B2(new_n935), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(new_n638), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n932), .A2(new_n935), .A3(KEYINPUT127), .ZN(new_n961));
  OAI21_X1  g760(.A(G218gat), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n939), .A2(new_n335), .A3(new_n638), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1355gat));
endmodule


