

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U323 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U324 ( .A(KEYINPUT46), .B(KEYINPUT116), .ZN(n387) );
  XNOR2_X1 U325 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U326 ( .A(G120GAT), .B(G71GAT), .Z(n439) );
  XNOR2_X1 U327 ( .A(n366), .B(n365), .ZN(n369) );
  AND2_X1 U328 ( .A1(n493), .A2(n580), .ZN(n494) );
  XNOR2_X1 U329 ( .A(n464), .B(KEYINPUT26), .ZN(n570) );
  XNOR2_X1 U330 ( .A(n494), .B(KEYINPUT37), .ZN(n518) );
  XNOR2_X1 U331 ( .A(n455), .B(n454), .ZN(n531) );
  XNOR2_X1 U332 ( .A(KEYINPUT109), .B(n497), .ZN(n504) );
  XNOR2_X1 U333 ( .A(n457), .B(KEYINPUT124), .ZN(n458) );
  XNOR2_X1 U334 ( .A(n459), .B(n458), .ZN(G1350GAT) );
  XOR2_X1 U335 ( .A(G211GAT), .B(G78GAT), .Z(n292) );
  XNOR2_X1 U336 ( .A(G127GAT), .B(G71GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U338 ( .A(G57GAT), .B(KEYINPUT13), .Z(n367) );
  XOR2_X1 U339 ( .A(n293), .B(n367), .Z(n295) );
  XNOR2_X1 U340 ( .A(G183GAT), .B(G155GAT), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n301) );
  XOR2_X1 U342 ( .A(KEYINPUT68), .B(G1GAT), .Z(n297) );
  XNOR2_X1 U343 ( .A(G22GAT), .B(G15GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n370) );
  XOR2_X1 U345 ( .A(n370), .B(KEYINPUT12), .Z(n299) );
  NAND2_X1 U346 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U348 ( .A(n301), .B(n300), .Z(n309) );
  XOR2_X1 U349 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n303) );
  XNOR2_X1 U350 ( .A(G8GAT), .B(G64GAT), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U352 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n305) );
  XNOR2_X1 U353 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n580) );
  XOR2_X1 U357 ( .A(KEYINPUT0), .B(KEYINPUT83), .Z(n311) );
  XNOR2_X1 U358 ( .A(KEYINPUT82), .B(G127GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U360 ( .A(G113GAT), .B(n312), .Z(n443) );
  XOR2_X1 U361 ( .A(G134GAT), .B(KEYINPUT74), .Z(n393) );
  XOR2_X1 U362 ( .A(G85GAT), .B(G162GAT), .Z(n314) );
  XNOR2_X1 U363 ( .A(G29GAT), .B(G148GAT), .ZN(n313) );
  XNOR2_X1 U364 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U365 ( .A(n393), .B(n315), .Z(n317) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n443), .B(n318), .ZN(n334) );
  XOR2_X1 U369 ( .A(KEYINPUT95), .B(KEYINPUT4), .Z(n323) );
  XOR2_X1 U370 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n320) );
  XNOR2_X1 U371 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U373 ( .A(G141GAT), .B(n321), .Z(n435) );
  XNOR2_X1 U374 ( .A(n435), .B(KEYINPUT5), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U376 ( .A(KEYINPUT6), .B(KEYINPUT91), .Z(n325) );
  XNOR2_X1 U377 ( .A(G120GAT), .B(KEYINPUT1), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U379 ( .A(n327), .B(n326), .Z(n332) );
  XOR2_X1 U380 ( .A(G57GAT), .B(KEYINPUT92), .Z(n329) );
  XNOR2_X1 U381 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U383 ( .A(G1GAT), .B(n330), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n334), .B(n333), .ZN(n519) );
  XOR2_X1 U386 ( .A(G169GAT), .B(G8GAT), .Z(n371) );
  XOR2_X1 U387 ( .A(G36GAT), .B(G190GAT), .Z(n391) );
  XNOR2_X1 U388 ( .A(n371), .B(n391), .ZN(n338) );
  XNOR2_X1 U389 ( .A(G64GAT), .B(G92GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(G176GAT), .B(G204GAT), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n354) );
  INV_X1 U392 ( .A(n354), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n344) );
  XOR2_X1 U394 ( .A(G211GAT), .B(KEYINPUT21), .Z(n340) );
  XNOR2_X1 U395 ( .A(G197GAT), .B(G218GAT), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n423) );
  XOR2_X1 U397 ( .A(KEYINPUT100), .B(n423), .Z(n342) );
  NAND2_X1 U398 ( .A1(G226GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U400 ( .A(n344), .B(n343), .Z(n352) );
  XOR2_X1 U401 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n346) );
  XNOR2_X1 U402 ( .A(KEYINPUT86), .B(G183GAT), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U404 ( .A(KEYINPUT17), .B(n347), .Z(n453) );
  XOR2_X1 U405 ( .A(KEYINPUT99), .B(KEYINPUT97), .Z(n349) );
  XNOR2_X1 U406 ( .A(KEYINPUT98), .B(KEYINPUT96), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n453), .B(n350), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n466) );
  XOR2_X1 U410 ( .A(G99GAT), .B(G85GAT), .Z(n392) );
  NAND2_X1 U411 ( .A1(n392), .A2(n337), .ZN(n356) );
  INV_X1 U412 ( .A(n392), .ZN(n353) );
  NAND2_X1 U413 ( .A1(n354), .A2(n353), .ZN(n355) );
  NAND2_X1 U414 ( .A1(n356), .A2(n355), .ZN(n358) );
  AND2_X1 U415 ( .A1(G230GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U417 ( .A(KEYINPUT70), .B(n359), .Z(n366) );
  XNOR2_X1 U418 ( .A(G106GAT), .B(G78GAT), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n360), .B(G148GAT), .ZN(n427) );
  XNOR2_X1 U420 ( .A(n427), .B(KEYINPUT71), .ZN(n364) );
  XOR2_X1 U421 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n362) );
  XNOR2_X1 U422 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n361) );
  XOR2_X1 U423 ( .A(n362), .B(n361), .Z(n363) );
  XNOR2_X1 U424 ( .A(n439), .B(n367), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n412) );
  XNOR2_X1 U426 ( .A(n412), .B(KEYINPUT41), .ZN(n548) );
  XOR2_X1 U427 ( .A(n371), .B(n370), .Z(n373) );
  NAND2_X1 U428 ( .A1(G229GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U430 ( .A(n374), .B(KEYINPUT69), .Z(n378) );
  XOR2_X1 U431 ( .A(G29GAT), .B(G43GAT), .Z(n376) );
  XNOR2_X1 U432 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n396) );
  XNOR2_X1 U434 ( .A(n396), .B(KEYINPUT29), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n386) );
  XOR2_X1 U436 ( .A(G141GAT), .B(G197GAT), .Z(n380) );
  XNOR2_X1 U437 ( .A(G36GAT), .B(G50GAT), .ZN(n379) );
  XNOR2_X1 U438 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U439 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n382) );
  XNOR2_X1 U440 ( .A(G113GAT), .B(KEYINPUT30), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U442 ( .A(n384), .B(n383), .Z(n385) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n572) );
  INV_X1 U444 ( .A(n572), .ZN(n533) );
  NAND2_X1 U445 ( .A1(n548), .A2(n533), .ZN(n388) );
  NAND2_X1 U446 ( .A1(n389), .A2(n580), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n390), .B(KEYINPUT117), .ZN(n409) );
  XOR2_X1 U448 ( .A(n392), .B(n391), .Z(n395) );
  XOR2_X1 U449 ( .A(G50GAT), .B(G162GAT), .Z(n424) );
  XNOR2_X1 U450 ( .A(n424), .B(n393), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n400) );
  XOR2_X1 U452 ( .A(G92GAT), .B(n396), .Z(n398) );
  NAND2_X1 U453 ( .A1(G232GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U455 ( .A(n400), .B(n399), .Z(n408) );
  XOR2_X1 U456 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n402) );
  XNOR2_X1 U457 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U459 ( .A(KEYINPUT65), .B(KEYINPUT11), .Z(n404) );
  XNOR2_X1 U460 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n408), .B(n407), .ZN(n566) );
  NAND2_X1 U464 ( .A1(n409), .A2(n566), .ZN(n411) );
  XNOR2_X1 U465 ( .A(KEYINPUT47), .B(KEYINPUT118), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n419) );
  XNOR2_X1 U467 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n415) );
  INV_X1 U468 ( .A(n566), .ZN(n557) );
  XOR2_X1 U469 ( .A(KEYINPUT36), .B(KEYINPUT108), .Z(n413) );
  XNOR2_X1 U470 ( .A(n557), .B(n413), .ZN(n583) );
  NOR2_X1 U471 ( .A1(n583), .A2(n580), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n416) );
  NAND2_X1 U473 ( .A1(n412), .A2(n416), .ZN(n417) );
  NOR2_X1 U474 ( .A1(n533), .A2(n417), .ZN(n418) );
  NOR2_X1 U475 ( .A1(n419), .A2(n418), .ZN(n420) );
  XNOR2_X1 U476 ( .A(KEYINPUT48), .B(n420), .ZN(n529) );
  NOR2_X1 U477 ( .A1(n466), .A2(n529), .ZN(n421) );
  XOR2_X1 U478 ( .A(KEYINPUT54), .B(n421), .Z(n422) );
  NOR2_X1 U479 ( .A1(n519), .A2(n422), .ZN(n571) );
  XOR2_X1 U480 ( .A(KEYINPUT23), .B(n423), .Z(n426) );
  XNOR2_X1 U481 ( .A(G22GAT), .B(n424), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n431) );
  XOR2_X1 U483 ( .A(n427), .B(KEYINPUT90), .Z(n429) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U486 ( .A(n431), .B(n430), .Z(n437) );
  XOR2_X1 U487 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n433) );
  XNOR2_X1 U488 ( .A(G204GAT), .B(KEYINPUT88), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n468) );
  NAND2_X1 U492 ( .A1(n571), .A2(n468), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n438), .B(KEYINPUT55), .ZN(n456) );
  XOR2_X1 U494 ( .A(n439), .B(KEYINPUT87), .Z(n441) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U497 ( .A(n442), .B(G99GAT), .Z(n445) );
  XNOR2_X1 U498 ( .A(G43GAT), .B(n443), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U500 ( .A(G134GAT), .B(G190GAT), .Z(n447) );
  XNOR2_X1 U501 ( .A(G169GAT), .B(G15GAT), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(n449), .B(n448), .Z(n455) );
  XOR2_X1 U504 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n451) );
  XNOR2_X1 U505 ( .A(G176GAT), .B(KEYINPUT20), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n454) );
  NAND2_X1 U508 ( .A1(n456), .A2(n531), .ZN(n565) );
  NOR2_X1 U509 ( .A1(n580), .A2(n565), .ZN(n459) );
  INV_X1 U510 ( .A(G183GAT), .ZN(n457) );
  NAND2_X1 U511 ( .A1(n533), .A2(n412), .ZN(n495) );
  NOR2_X1 U512 ( .A1(n580), .A2(n557), .ZN(n461) );
  XNOR2_X1 U513 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U515 ( .A(KEYINPUT16), .B(n462), .Z(n479) );
  XOR2_X1 U516 ( .A(n468), .B(KEYINPUT28), .Z(n524) );
  XOR2_X1 U517 ( .A(n466), .B(KEYINPUT27), .Z(n465) );
  NAND2_X1 U518 ( .A1(n519), .A2(n465), .ZN(n544) );
  NOR2_X1 U519 ( .A1(n524), .A2(n544), .ZN(n530) );
  XNOR2_X1 U520 ( .A(KEYINPUT101), .B(n530), .ZN(n463) );
  NOR2_X1 U521 ( .A1(n531), .A2(n463), .ZN(n477) );
  NOR2_X1 U522 ( .A1(n468), .A2(n531), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n570), .A2(n465), .ZN(n471) );
  INV_X1 U524 ( .A(n466), .ZN(n521) );
  NAND2_X1 U525 ( .A1(n531), .A2(n521), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n469) );
  XOR2_X1 U527 ( .A(KEYINPUT25), .B(n469), .Z(n470) );
  NAND2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n473) );
  INV_X1 U529 ( .A(n519), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U531 ( .A(KEYINPUT102), .B(n474), .ZN(n475) );
  INV_X1 U532 ( .A(n475), .ZN(n476) );
  NOR2_X1 U533 ( .A1(n477), .A2(n476), .ZN(n492) );
  INV_X1 U534 ( .A(n492), .ZN(n478) );
  NAND2_X1 U535 ( .A1(n479), .A2(n478), .ZN(n507) );
  NOR2_X1 U536 ( .A1(n495), .A2(n507), .ZN(n489) );
  NAND2_X1 U537 ( .A1(n489), .A2(n519), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n483) );
  NAND2_X1 U541 ( .A1(n489), .A2(n521), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(n484), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT35), .B(KEYINPUT106), .Z(n486) );
  NAND2_X1 U545 ( .A1(n489), .A2(n531), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n488) );
  XOR2_X1 U547 ( .A(G15GAT), .B(KEYINPUT105), .Z(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  XOR2_X1 U549 ( .A(G22GAT), .B(KEYINPUT107), .Z(n491) );
  NAND2_X1 U550 ( .A1(n489), .A2(n524), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(G1327GAT) );
  XOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT110), .Z(n499) );
  NOR2_X1 U553 ( .A1(n583), .A2(n492), .ZN(n493) );
  NOR2_X1 U554 ( .A1(n518), .A2(n495), .ZN(n496) );
  XOR2_X1 U555 ( .A(KEYINPUT38), .B(n496), .Z(n497) );
  NAND2_X1 U556 ( .A1(n519), .A2(n504), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U558 ( .A(KEYINPUT39), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n504), .A2(n521), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n501), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U561 ( .A1(n504), .A2(n531), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n504), .A2(n524), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n505), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n509) );
  XOR2_X1 U567 ( .A(KEYINPUT112), .B(n548), .Z(n561) );
  NOR2_X1 U568 ( .A1(n561), .A2(n533), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n506), .B(KEYINPUT113), .ZN(n517) );
  NOR2_X1 U570 ( .A1(n517), .A2(n507), .ZN(n513) );
  NAND2_X1 U571 ( .A1(n513), .A2(n519), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n521), .A2(n513), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n531), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT114), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U579 ( .A1(n513), .A2(n524), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(n516), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n519), .A2(n525), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n525), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n522), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n525), .A2(n531), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT115), .Z(n527) );
  NAND2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  XOR2_X1 U593 ( .A(G113GAT), .B(KEYINPUT119), .Z(n535) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U595 ( .A1(n529), .A2(n532), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n541), .A2(n533), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n535), .B(n534), .ZN(G1340GAT) );
  INV_X1 U598 ( .A(n541), .ZN(n538) );
  NOR2_X1 U599 ( .A1(n561), .A2(n538), .ZN(n537) );
  XNOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  NOR2_X1 U602 ( .A1(n580), .A2(n538), .ZN(n539) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(n539), .Z(n540) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U606 ( .A1(n541), .A2(n557), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NOR2_X1 U608 ( .A1(n529), .A2(n544), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n545), .A2(n570), .ZN(n554) );
  NOR2_X1 U610 ( .A1(n572), .A2(n554), .ZN(n546) );
  XOR2_X1 U611 ( .A(KEYINPUT120), .B(n546), .Z(n547) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n550) );
  INV_X1 U614 ( .A(n554), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n556), .A2(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U617 ( .A(n551), .B(KEYINPUT121), .Z(n553) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n580), .A2(n554), .ZN(n555) );
  XOR2_X1 U621 ( .A(G155GAT), .B(n555), .Z(G1346GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U624 ( .A1(n572), .A2(n565), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1348GAT) );
  NOR2_X1 U627 ( .A1(n565), .A2(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(n564), .ZN(G1349GAT) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(n569), .ZN(G1351GAT) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n582) );
  NOR2_X1 U636 ( .A1(n572), .A2(n582), .ZN(n577) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n574) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(KEYINPUT126), .B(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  NOR2_X1 U642 ( .A1(n412), .A2(n582), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n582), .ZN(n581) );
  XOR2_X1 U646 ( .A(G211GAT), .B(n581), .Z(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

