//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1076, new_n1077, new_n1078;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XOR2_X1   g002(.A(G78gat), .B(G106gat), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT2), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT75), .ZN(new_n210));
  XNOR2_X1  g009(.A(G155gat), .B(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n212), .B(KEYINPUT2), .C1(new_n207), .C2(new_n208), .ZN(new_n213));
  INV_X1    g012(.A(G148gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G141gat), .ZN(new_n215));
  INV_X1    g014(.A(G141gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G148gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n210), .A2(new_n211), .A3(new_n213), .A4(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n216), .A2(G148gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n214), .A2(G141gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n211), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT74), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT2), .B1(new_n215), .B2(new_n217), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT74), .ZN(new_n227));
  NOR3_X1   g026(.A1(new_n226), .A2(new_n227), .A3(new_n211), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n206), .B(new_n219), .C1(new_n225), .C2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT29), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G197gat), .A2(G204gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(G197gat), .A2(G204gat), .ZN(new_n234));
  AND2_X1   g033(.A1(G211gat), .A2(G218gat), .ZN(new_n235));
  OAI22_X1  g034(.A1(new_n233), .A2(new_n234), .B1(new_n235), .B2(KEYINPUT22), .ZN(new_n236));
  NOR2_X1   g035(.A1(G211gat), .A2(G218gat), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n235), .A2(new_n237), .A3(KEYINPUT72), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G197gat), .ZN(new_n240));
  INV_X1    g039(.A(G204gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT22), .ZN(new_n243));
  NAND2_X1  g042(.A1(G211gat), .A2(G218gat), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n242), .A2(new_n232), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(G211gat), .A2(G218gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT72), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n244), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n239), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n219), .B1(new_n225), .B2(new_n228), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n245), .B1(new_n244), .B2(new_n246), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n246), .A2(new_n244), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n230), .B1(new_n236), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n206), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G228gat), .ZN(new_n259));
  INV_X1    g058(.A(G233gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT79), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n262), .B1(new_n231), .B2(new_n250), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n236), .A2(new_n238), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n245), .A2(new_n248), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT29), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n252), .B1(KEYINPUT3), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n264), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n250), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(new_n229), .B2(new_n230), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n230), .B1(new_n239), .B2(new_n249), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT74), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n227), .B1(new_n226), .B2(new_n211), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n273), .A2(new_n206), .B1(new_n276), .B2(new_n219), .ZN(new_n277));
  NOR4_X1   g076(.A1(new_n272), .A2(new_n277), .A3(KEYINPUT79), .A4(new_n262), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n263), .B1(new_n270), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G22gat), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n218), .A2(new_n211), .A3(new_n213), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n275), .A2(new_n274), .B1(new_n281), .B2(new_n210), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT29), .B1(new_n282), .B2(new_n206), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n261), .B(new_n269), .C1(new_n283), .C2(new_n271), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT79), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n264), .A3(new_n269), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G22gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(new_n288), .A3(new_n263), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n205), .B1(new_n290), .B2(KEYINPUT78), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT78), .ZN(new_n292));
  AOI211_X1 g091(.A(new_n292), .B(new_n204), .C1(new_n280), .C2(new_n289), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n203), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n261), .B1(new_n251), .B2(new_n257), .ZN(new_n295));
  AOI211_X1 g094(.A(G22gat), .B(new_n295), .C1(new_n285), .C2(new_n286), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n288), .B1(new_n287), .B2(new_n263), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT78), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n204), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n290), .A2(KEYINPUT78), .A3(new_n205), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n202), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT0), .B(G57gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(G85gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G1gat), .B(G29gat), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n304), .B(new_n305), .Z(new_n306));
  NAND2_X1  g105(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n307));
  INV_X1    g106(.A(G127gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G134gat), .ZN(new_n309));
  INV_X1    g108(.A(G134gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G127gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G120gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G113gat), .ZN(new_n314));
  INV_X1    g113(.A(G113gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G120gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n312), .B1(KEYINPUT69), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G113gat), .B(G120gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT69), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT1), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT68), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT68), .B1(new_n314), .B2(new_n316), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT1), .ZN(new_n326));
  INV_X1    g125(.A(new_n309), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT67), .B(G134gat), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(G127gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n322), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n307), .A2(new_n330), .A3(new_n229), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT68), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(new_n323), .ZN(new_n335));
  XOR2_X1   g134(.A(KEYINPUT67), .B(G134gat), .Z(new_n336));
  OAI21_X1  g135(.A(new_n309), .B1(new_n336), .B2(new_n308), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n335), .A2(new_n337), .B1(new_n318), .B2(new_n321), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n282), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n282), .B2(new_n338), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n282), .A2(new_n338), .A3(new_n343), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n331), .B(new_n342), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT5), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n252), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n339), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n347), .B1(new_n349), .B2(new_n341), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n341), .A2(KEYINPUT5), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n331), .B(new_n352), .C1(new_n344), .C2(new_n345), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n306), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT6), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n351), .A2(new_n306), .A3(new_n353), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n354), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n339), .A2(KEYINPUT4), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n282), .A2(new_n338), .A3(new_n343), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n338), .B1(new_n206), .B2(new_n282), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n362), .A2(new_n363), .B1(new_n364), .B2(new_n307), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n346), .A2(new_n350), .B1(new_n365), .B2(new_n352), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT6), .B1(new_n366), .B2(new_n306), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT76), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n356), .B1(new_n361), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G226gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(new_n260), .ZN(new_n371));
  NAND2_X1  g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372));
  INV_X1    g171(.A(G169gat), .ZN(new_n373));
  INV_X1    g172(.A(G176gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT26), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT26), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(G169gat), .B2(G176gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n372), .B(new_n375), .C1(new_n377), .C2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G183gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(KEYINPUT27), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT66), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(KEYINPUT65), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT65), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(KEYINPUT27), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT27), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G183gat), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n386), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n386), .B1(new_n388), .B2(G183gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT66), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n385), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G190gat), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT28), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n388), .A2(G183gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(new_n383), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(KEYINPUT28), .A3(new_n394), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n381), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT23), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(new_n373), .A3(new_n374), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n379), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT25), .B1(new_n404), .B2(KEYINPUT64), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n372), .A2(KEYINPUT24), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n382), .A2(new_n394), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT24), .A3(new_n372), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n405), .B(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n400), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n371), .B1(new_n411), .B2(new_n230), .ZN(new_n412));
  AOI211_X1 g211(.A(new_n370), .B(new_n260), .C1(new_n400), .C2(new_n410), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n250), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n371), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n400), .B2(new_n410), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n415), .B(new_n271), .C1(new_n371), .C2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418));
  INV_X1    g217(.A(G64gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G92gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n414), .A2(new_n417), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT73), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT30), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n423), .B1(new_n414), .B2(new_n417), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT30), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(KEYINPUT73), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT77), .B1(new_n369), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n354), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(new_n367), .B2(KEYINPUT76), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n359), .A2(new_n360), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n355), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n424), .A2(KEYINPUT73), .A3(new_n429), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n429), .B1(new_n424), .B2(KEYINPUT73), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n437), .A2(new_n438), .A3(new_n427), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT77), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n436), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT28), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n389), .A2(new_n386), .A3(KEYINPUT66), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT65), .B1(new_n396), .B2(new_n383), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n384), .B1(new_n387), .B2(new_n386), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n442), .B1(new_n446), .B2(G190gat), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n380), .B1(new_n447), .B2(new_n398), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n405), .A2(new_n409), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n405), .A2(new_n409), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT70), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT70), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n400), .A2(new_n410), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n330), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G227gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(new_n260), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n411), .A2(KEYINPUT70), .A3(new_n338), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT32), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT33), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G15gat), .B(G43gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(G71gat), .B(G99gat), .ZN(new_n464));
  XOR2_X1   g263(.A(new_n463), .B(new_n464), .Z(new_n465));
  NAND3_X1  g264(.A1(new_n460), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n465), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n459), .B(KEYINPUT32), .C1(new_n461), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n455), .A2(new_n458), .ZN(new_n470));
  INV_X1    g269(.A(new_n457), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT34), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT34), .ZN(new_n473));
  AOI211_X1 g272(.A(new_n473), .B(new_n457), .C1(new_n455), .C2(new_n458), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT71), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n470), .A2(new_n471), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n473), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n470), .A2(KEYINPUT34), .A3(new_n471), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT71), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(new_n468), .A3(new_n466), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n302), .A2(new_n432), .A3(new_n441), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n472), .A2(new_n474), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(new_n466), .A3(new_n468), .ZN(new_n487));
  INV_X1    g286(.A(new_n486), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n294), .A2(new_n301), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n492));
  INV_X1    g291(.A(new_n306), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT80), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n366), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n351), .A2(new_n494), .A3(new_n353), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n367), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT82), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n355), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n354), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n492), .B1(new_n501), .B2(new_n431), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n439), .A2(new_n503), .A3(KEYINPUT83), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n490), .A2(new_n491), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT81), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n414), .A2(new_n417), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT37), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n414), .A2(new_n417), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n422), .A3(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n512), .A2(KEYINPUT38), .ZN(new_n513));
  INV_X1    g312(.A(new_n424), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(new_n512), .B2(KEYINPUT38), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n501), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n331), .B1(new_n345), .B2(new_n344), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n341), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n518), .B(KEYINPUT39), .C1(new_n341), .C2(new_n349), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n519), .B(new_n306), .C1(KEYINPUT39), .C2(new_n518), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT40), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n495), .A2(new_n496), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n521), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n431), .A2(new_n522), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n516), .A2(new_n302), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n477), .A2(new_n482), .A3(KEYINPUT36), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n489), .A2(new_n487), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(KEYINPUT36), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n432), .A2(new_n441), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n526), .B(new_n529), .C1(new_n530), .C2(new_n302), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n506), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G57gat), .B(G64gat), .Z(new_n533));
  NAND2_X1  g332(.A1(G71gat), .A2(G78gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(KEYINPUT92), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G71gat), .B(G78gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n533), .A2(KEYINPUT92), .A3(new_n538), .A4(new_n536), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT93), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT93), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT21), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G127gat), .B(G155gat), .Z(new_n548));
  XOR2_X1   g347(.A(new_n547), .B(new_n548), .Z(new_n549));
  NOR2_X1   g348(.A1(new_n545), .A2(new_n546), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT88), .ZN(new_n551));
  AND2_X1   g350(.A1(G15gat), .A2(G22gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(G15gat), .A2(G22gat), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT87), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G15gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n288), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT87), .ZN(new_n557));
  NAND2_X1  g356(.A1(G15gat), .A2(G22gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G1gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT16), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n554), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(G1gat), .B1(new_n554), .B2(new_n559), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n562), .A2(new_n563), .A3(G8gat), .ZN(new_n564));
  INV_X1    g363(.A(G8gat), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT87), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n557), .B1(new_n556), .B2(new_n558), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n560), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n554), .A2(new_n559), .A3(new_n561), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n551), .B1(new_n564), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(G8gat), .B1(new_n562), .B2(new_n563), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n565), .A3(new_n569), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT88), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  OR3_X1    g374(.A1(new_n550), .A2(KEYINPUT94), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT94), .B1(new_n550), .B2(new_n575), .ZN(new_n577));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n579), .B1(new_n576), .B2(new_n577), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n549), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n582), .ZN(new_n584));
  INV_X1    g383(.A(new_n549), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n588));
  XNOR2_X1  g387(.A(G183gat), .B(G211gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n583), .A2(new_n586), .A3(new_n590), .ZN(new_n593));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n595), .A2(new_n596), .B1(new_n597), .B2(KEYINPUT8), .ZN(new_n598));
  INV_X1    g397(.A(G85gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n421), .ZN(new_n600));
  INV_X1    g399(.A(new_n595), .ZN(new_n601));
  NAND2_X1  g400(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n598), .B(new_n600), .C1(new_n603), .C2(new_n596), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  OR2_X1    g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT97), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT17), .ZN(new_n610));
  INV_X1    g409(.A(G43gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT85), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT85), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(G43gat), .ZN(new_n614));
  INV_X1    g413(.A(G50gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(KEYINPUT86), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT86), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(G50gat), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n617), .A2(new_n619), .A3(new_n611), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT15), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT15), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n611), .A2(new_n615), .ZN(new_n623));
  NAND2_X1  g422(.A1(G43gat), .A2(G50gat), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(G29gat), .ZN(new_n626));
  INV_X1    g425(.A(G36gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n627), .A3(KEYINPUT14), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT14), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(G29gat), .B2(G36gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n626), .A2(new_n627), .ZN(new_n632));
  NOR4_X1   g431(.A1(new_n621), .A2(new_n625), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n625), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT84), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n628), .A2(new_n630), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n632), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n631), .A2(KEYINPUT84), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n634), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n610), .B1(new_n633), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n621), .ZN(new_n643));
  INV_X1    g442(.A(new_n631), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n643), .A2(new_n634), .A3(new_n644), .A4(new_n637), .ZN(new_n645));
  INV_X1    g444(.A(new_n640), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n625), .B1(new_n646), .B2(new_n638), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n647), .A3(KEYINPUT17), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n609), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n608), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n645), .A2(new_n647), .ZN(new_n653));
  NAND2_X1  g452(.A1(G232gat), .A2(G233gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT95), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n652), .A2(new_n653), .B1(KEYINPUT41), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n649), .A2(new_n651), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n651), .B1(new_n649), .B2(new_n657), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n594), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  INV_X1    g461(.A(new_n594), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n663), .A3(new_n658), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n656), .A2(KEYINPUT41), .ZN(new_n665));
  XNOR2_X1  g464(.A(G134gat), .B(G162gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n661), .A2(new_n664), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n661), .A2(new_n664), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n592), .A2(new_n593), .A3(new_n670), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(G229gat), .A2(G233gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n564), .A2(new_n570), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n642), .A2(new_n677), .A3(new_n648), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n572), .A2(KEYINPUT88), .A3(new_n573), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT88), .B1(new_n572), .B2(new_n573), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n653), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT89), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n575), .A2(KEYINPUT89), .A3(new_n653), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n676), .B(new_n678), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT90), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT18), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n575), .B2(new_n653), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n675), .B(KEYINPUT91), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT13), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n678), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n688), .A2(new_n675), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT18), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(KEYINPUT90), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n687), .A2(new_n692), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT11), .B(G169gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G197gat), .ZN(new_n699));
  XOR2_X1   g498(.A(G113gat), .B(G141gat), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT12), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n687), .A2(new_n702), .A3(new_n696), .A4(new_n692), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT101), .B(KEYINPUT10), .Z(new_n707));
  NAND2_X1  g506(.A1(new_n540), .A2(new_n541), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT93), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n710), .A2(new_n542), .B1(new_n606), .B2(new_n607), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n606), .A2(new_n708), .A3(new_n607), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n707), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n542), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(new_n652), .A3(KEYINPUT10), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(G230gat), .A2(G233gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n711), .A2(new_n717), .A3(new_n712), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(G120gat), .B(G148gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(new_n374), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(new_n241), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n726));
  INV_X1    g525(.A(new_n717), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n713), .B2(new_n715), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n719), .ZN(new_n729));
  INV_X1    g528(.A(new_n724), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n726), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR4_X1   g530(.A1(new_n728), .A2(new_n719), .A3(KEYINPUT102), .A4(new_n724), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n725), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n706), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n674), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n532), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n436), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n560), .ZN(G1324gat));
  NOR2_X1   g538(.A1(new_n737), .A2(new_n439), .ZN(new_n740));
  OR2_X1    g539(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n743), .A2(KEYINPUT42), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(KEYINPUT42), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n744), .B(new_n745), .C1(new_n565), .C2(new_n740), .ZN(G1325gat));
  OAI21_X1  g545(.A(G15gat), .B1(new_n737), .B2(new_n529), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n532), .A2(new_n555), .A3(new_n528), .A4(new_n736), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT103), .Z(G1326gat));
  NOR2_X1   g549(.A1(new_n737), .A2(new_n302), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT43), .B(G22gat), .Z(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1327gat));
  NAND2_X1  g552(.A1(new_n673), .A2(new_n670), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n532), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n592), .A2(new_n593), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n735), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n626), .A3(new_n369), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n761), .A2(KEYINPUT104), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(KEYINPUT104), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n754), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(KEYINPUT44), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n506), .A2(KEYINPUT105), .A3(new_n531), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT105), .B1(new_n506), .B2(new_n531), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n755), .A2(KEYINPUT44), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n759), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G29gat), .B1(new_n774), .B2(new_n436), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n762), .A2(KEYINPUT45), .A3(new_n763), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n766), .A2(new_n775), .A3(new_n776), .ZN(G1328gat));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n627), .A3(new_n431), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT46), .Z(new_n779));
  OAI21_X1  g578(.A(G36gat), .B1(new_n774), .B2(new_n439), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(G1329gat));
  NAND2_X1  g580(.A1(new_n612), .A2(new_n614), .ZN(new_n782));
  INV_X1    g581(.A(new_n529), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n773), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n767), .B1(new_n506), .B2(new_n531), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n785), .A2(new_n528), .A3(new_n782), .A4(new_n758), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(KEYINPUT106), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI211_X1 g591(.A(KEYINPUT107), .B(KEYINPUT47), .C1(new_n786), .C2(KEYINPUT106), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n784), .A2(new_n787), .B1(new_n793), .B2(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1330gat));
  INV_X1    g596(.A(new_n302), .ZN(new_n798));
  INV_X1    g597(.A(new_n768), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT105), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n490), .A2(new_n502), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n504), .A2(new_n491), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n801), .A2(new_n802), .B1(KEYINPUT35), .B2(new_n484), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n526), .A2(new_n529), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n302), .B1(new_n432), .B2(new_n441), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n800), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n506), .A2(KEYINPUT105), .A3(new_n531), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n799), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n785), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n798), .B(new_n758), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n617), .A2(new_n619), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n771), .A2(new_n772), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n817), .A2(KEYINPUT108), .A3(new_n798), .A4(new_n758), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n814), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  NOR4_X1   g618(.A1(new_n755), .A2(new_n302), .A3(new_n816), .A4(new_n759), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(KEYINPUT48), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT48), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n815), .B1(new_n773), .B2(new_n798), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n820), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(G1331gat));
  NAND2_X1  g625(.A1(new_n807), .A2(new_n808), .ZN(new_n827));
  INV_X1    g626(.A(new_n674), .ZN(new_n828));
  INV_X1    g627(.A(new_n706), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n733), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n369), .B(KEYINPUT109), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(G57gat), .Z(G1332gat));
  AOI21_X1  g632(.A(new_n439), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT110), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n674), .B(new_n706), .C1(new_n807), .C2(new_n808), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT110), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n837), .A2(new_n838), .A3(new_n733), .A4(new_n834), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n840), .B(new_n841), .ZN(G1333gat));
  OAI21_X1  g641(.A(G71gat), .B1(new_n830), .B2(new_n529), .ZN(new_n843));
  INV_X1    g642(.A(G71gat), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n837), .A2(new_n844), .A3(new_n528), .A4(new_n733), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT50), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n846), .B(new_n847), .ZN(G1334gat));
  NOR2_X1   g647(.A1(new_n830), .A2(new_n302), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g649(.A1(new_n757), .A2(new_n706), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n733), .B(new_n851), .C1(new_n809), .C2(new_n811), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n852), .A2(new_n599), .A3(new_n436), .ZN(new_n853));
  INV_X1    g652(.A(new_n851), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n755), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n785), .A2(KEYINPUT111), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT51), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n851), .B1(new_n785), .B2(KEYINPUT111), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n860));
  AOI211_X1 g659(.A(new_n855), .B(new_n767), .C1(new_n506), .C2(new_n531), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n369), .B(new_n733), .C1(new_n858), .C2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n853), .B1(new_n599), .B2(new_n863), .ZN(G1336gat));
  AOI211_X1 g663(.A(new_n734), .B(new_n854), .C1(new_n771), .C2(new_n772), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n421), .B1(new_n865), .B2(new_n431), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n439), .A2(G92gat), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n860), .B1(new_n859), .B2(new_n861), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n526), .A2(new_n529), .ZN(new_n870));
  INV_X1    g669(.A(new_n805), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n870), .A2(new_n871), .B1(new_n485), .B2(new_n505), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n855), .B1(new_n872), .B2(new_n767), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n873), .A2(new_n857), .A3(KEYINPUT51), .A4(new_n851), .ZN(new_n874));
  AOI211_X1 g673(.A(new_n734), .B(new_n868), .C1(new_n869), .C2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT52), .B1(new_n866), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n733), .B(new_n867), .C1(new_n858), .C2(new_n862), .ZN(new_n877));
  OAI21_X1  g676(.A(G92gat), .B1(new_n852), .B2(new_n439), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT52), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n876), .A2(new_n880), .ZN(G1337gat));
  AOI21_X1  g680(.A(G99gat), .B1(new_n489), .B2(new_n487), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n733), .B(new_n882), .C1(new_n858), .C2(new_n862), .ZN(new_n883));
  OAI21_X1  g682(.A(G99gat), .B1(new_n852), .B2(new_n529), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1338gat));
  OAI21_X1  g684(.A(G106gat), .B1(new_n852), .B2(new_n302), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n302), .A2(G106gat), .A3(new_n734), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT112), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n858), .B2(new_n862), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT53), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n886), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(G1339gat));
  NOR3_X1   g693(.A1(new_n674), .A2(new_n706), .A3(new_n733), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n713), .A2(new_n727), .A3(new_n715), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n718), .A2(new_n897), .A3(KEYINPUT54), .ZN(new_n898));
  XOR2_X1   g697(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n899));
  NAND2_X1  g698(.A1(new_n728), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n898), .A2(new_n724), .A3(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT55), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT102), .B1(new_n721), .B2(new_n724), .ZN(new_n904));
  INV_X1    g703(.A(new_n732), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n898), .A2(KEYINPUT55), .A3(new_n724), .A4(new_n900), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n689), .A2(new_n691), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n675), .B1(new_n688), .B2(new_n693), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n701), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n705), .A2(new_n911), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n754), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n706), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n733), .A2(new_n705), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT114), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT114), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n733), .A2(new_n705), .A3(new_n917), .A4(new_n911), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n914), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n913), .B1(new_n919), .B2(new_n767), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n896), .B1(new_n920), .B2(new_n757), .ZN(new_n921));
  INV_X1    g720(.A(new_n831), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n302), .A2(new_n483), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n439), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT116), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n315), .A3(new_n706), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n921), .A2(new_n490), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n436), .A2(new_n431), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  AOI211_X1 g731(.A(KEYINPUT115), .B(new_n315), .C1(new_n932), .C2(new_n706), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT115), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n706), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(G113gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n928), .B1(new_n933), .B2(new_n936), .ZN(G1340gat));
  NAND3_X1  g736(.A1(new_n927), .A2(new_n313), .A3(new_n733), .ZN(new_n938));
  OAI21_X1  g737(.A(G120gat), .B1(new_n931), .B2(new_n734), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1341gat));
  NOR3_X1   g739(.A1(new_n931), .A2(new_n308), .A3(new_n756), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT117), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n308), .B1(new_n925), .B2(new_n756), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(G1342gat));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT118), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n925), .A2(new_n336), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n754), .ZN(new_n950));
  NOR4_X1   g749(.A1(new_n925), .A2(KEYINPUT118), .A3(new_n336), .A4(new_n767), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n923), .A2(new_n439), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n953), .A2(new_n328), .A3(new_n924), .A4(new_n754), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT118), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n949), .A2(new_n948), .A3(new_n754), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT56), .ZN(new_n957));
  OAI21_X1  g756(.A(G134gat), .B1(new_n931), .B2(new_n767), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n952), .A2(new_n957), .A3(new_n958), .ZN(G1343gat));
  NAND2_X1  g758(.A1(new_n529), .A2(new_n930), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n906), .A2(new_n907), .ZN(new_n961));
  XOR2_X1   g760(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n962));
  NAND2_X1  g761(.A1(new_n901), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n706), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n754), .B1(new_n964), .B2(new_n915), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n756), .B1(new_n965), .B2(new_n913), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n798), .B1(new_n967), .B2(new_n895), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n960), .B1(new_n968), .B2(KEYINPUT57), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT57), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n921), .A2(new_n970), .A3(new_n798), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n969), .A2(new_n706), .A3(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT120), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n969), .A2(KEYINPUT120), .A3(new_n706), .A4(new_n971), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n974), .A2(G141gat), .A3(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT58), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n783), .A2(new_n302), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n923), .A2(new_n439), .A3(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n980), .A2(new_n216), .A3(new_n706), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n976), .A2(new_n977), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n972), .A2(G141gat), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(new_n981), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(KEYINPUT58), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n982), .A2(new_n985), .ZN(G1344gat));
  NAND3_X1  g785(.A1(new_n980), .A2(new_n214), .A3(new_n733), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT59), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n916), .A2(new_n918), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n990), .B1(new_n704), .B2(new_n705), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n767), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n754), .A2(new_n908), .A3(new_n912), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n757), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g793(.A(KEYINPUT57), .B(new_n798), .C1(new_n994), .C2(new_n895), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n995), .A2(KEYINPUT121), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT121), .ZN(new_n997));
  NAND4_X1  g796(.A1(new_n921), .A2(new_n997), .A3(KEYINPUT57), .A4(new_n798), .ZN(new_n998));
  AND3_X1   g797(.A1(new_n733), .A2(new_n705), .A3(new_n911), .ZN(new_n999));
  AOI22_X1  g798(.A1(new_n704), .A2(new_n705), .B1(new_n901), .B2(new_n962), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n999), .B1(new_n1000), .B2(new_n961), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n993), .B1(new_n1001), .B2(new_n754), .ZN(new_n1002));
  AOI211_X1 g801(.A(KEYINPUT122), .B(new_n895), .C1(new_n1002), .C2(new_n756), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT122), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1004), .B1(new_n966), .B2(new_n896), .ZN(new_n1005));
  NOR3_X1   g804(.A1(new_n1003), .A2(new_n1005), .A3(new_n302), .ZN(new_n1006));
  OAI211_X1 g805(.A(new_n996), .B(new_n998), .C1(new_n1006), .C2(KEYINPUT57), .ZN(new_n1007));
  INV_X1    g806(.A(new_n960), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1007), .A2(new_n733), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n988), .B1(new_n1009), .B2(G148gat), .ZN(new_n1010));
  AND2_X1   g809(.A1(new_n969), .A2(new_n971), .ZN(new_n1011));
  AOI211_X1 g810(.A(KEYINPUT59), .B(new_n214), .C1(new_n1011), .C2(new_n733), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n987), .B1(new_n1010), .B2(new_n1012), .ZN(G1345gat));
  NAND3_X1  g812(.A1(new_n1011), .A2(G155gat), .A3(new_n757), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n207), .B1(new_n979), .B2(new_n756), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g815(.A(new_n1016), .ZN(G1346gat));
  NAND3_X1  g816(.A1(new_n1011), .A2(G162gat), .A3(new_n754), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n208), .B1(new_n979), .B2(new_n767), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g819(.A(new_n1020), .ZN(G1347gat));
  NOR2_X1   g820(.A1(new_n922), .A2(new_n439), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n929), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g822(.A(G169gat), .B1(new_n1023), .B2(new_n829), .ZN(new_n1024));
  AND3_X1   g823(.A1(new_n921), .A2(new_n436), .A3(new_n431), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n1025), .A2(new_n373), .A3(new_n924), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1024), .B1(new_n829), .B2(new_n1026), .ZN(G1348gat));
  NOR3_X1   g826(.A1(new_n1023), .A2(new_n374), .A3(new_n734), .ZN(new_n1028));
  INV_X1    g827(.A(KEYINPUT123), .ZN(new_n1029));
  OR2_X1    g828(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1025), .A2(new_n924), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n374), .B1(new_n1031), .B2(new_n734), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1033));
  AND3_X1   g832(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .ZN(G1349gat));
  OAI21_X1  g833(.A(G183gat), .B1(new_n1023), .B2(new_n756), .ZN(new_n1035));
  NAND2_X1  g834(.A1(new_n757), .A2(new_n397), .ZN(new_n1036));
  OAI21_X1  g835(.A(new_n1035), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g836(.A(new_n1037), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g837(.A(KEYINPUT61), .ZN(new_n1039));
  NAND4_X1  g838(.A1(new_n921), .A2(new_n490), .A3(new_n754), .A4(new_n1022), .ZN(new_n1040));
  AOI21_X1  g839(.A(new_n1039), .B1(new_n1040), .B2(G190gat), .ZN(new_n1041));
  OR2_X1    g840(.A1(new_n1041), .A2(KEYINPUT124), .ZN(new_n1042));
  NAND3_X1  g841(.A1(new_n1040), .A2(new_n1039), .A3(G190gat), .ZN(new_n1043));
  INV_X1    g842(.A(KEYINPUT125), .ZN(new_n1044));
  OR2_X1    g843(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g844(.A1(new_n1041), .A2(KEYINPUT124), .ZN(new_n1046));
  NAND2_X1  g845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1047));
  NAND4_X1  g846(.A1(new_n1042), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  NAND3_X1  g847(.A1(new_n1025), .A2(new_n924), .A3(new_n754), .ZN(new_n1049));
  OAI21_X1  g848(.A(new_n1048), .B1(G190gat), .B2(new_n1049), .ZN(G1351gat));
  NOR3_X1   g849(.A1(new_n922), .A2(new_n783), .A3(new_n439), .ZN(new_n1051));
  NOR2_X1   g850(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1052));
  AOI21_X1  g851(.A(KEYINPUT57), .B1(new_n1052), .B2(new_n798), .ZN(new_n1053));
  NAND2_X1  g852(.A1(new_n996), .A2(new_n998), .ZN(new_n1054));
  OAI211_X1 g853(.A(new_n706), .B(new_n1051), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g854(.A1(new_n1055), .A2(KEYINPUT126), .ZN(new_n1056));
  INV_X1    g855(.A(KEYINPUT126), .ZN(new_n1057));
  NAND4_X1  g856(.A1(new_n1007), .A2(new_n1057), .A3(new_n706), .A4(new_n1051), .ZN(new_n1058));
  NAND3_X1  g857(.A1(new_n1056), .A2(new_n1058), .A3(G197gat), .ZN(new_n1059));
  NAND4_X1  g858(.A1(new_n1025), .A2(new_n240), .A3(new_n706), .A4(new_n978), .ZN(new_n1060));
  NAND2_X1  g859(.A1(new_n1059), .A2(new_n1060), .ZN(G1352gat));
  NAND3_X1  g860(.A1(new_n1007), .A2(new_n733), .A3(new_n1051), .ZN(new_n1062));
  XOR2_X1   g861(.A(KEYINPUT127), .B(G204gat), .Z(new_n1063));
  NAND2_X1  g862(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g863(.A1(new_n1025), .A2(new_n978), .ZN(new_n1065));
  NOR2_X1   g864(.A1(new_n734), .A2(new_n1063), .ZN(new_n1066));
  INV_X1    g865(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g866(.A(KEYINPUT62), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  OR3_X1    g867(.A1(new_n1065), .A2(KEYINPUT62), .A3(new_n1067), .ZN(new_n1069));
  NAND3_X1  g868(.A1(new_n1064), .A2(new_n1068), .A3(new_n1069), .ZN(G1353gat));
  OR3_X1    g869(.A1(new_n1065), .A2(G211gat), .A3(new_n756), .ZN(new_n1071));
  OAI211_X1 g870(.A(new_n757), .B(new_n1051), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1072));
  AND3_X1   g871(.A1(new_n1072), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1073));
  AOI21_X1  g872(.A(KEYINPUT63), .B1(new_n1072), .B2(G211gat), .ZN(new_n1074));
  OAI21_X1  g873(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(G1354gat));
  NAND3_X1  g874(.A1(new_n1007), .A2(new_n754), .A3(new_n1051), .ZN(new_n1076));
  NAND2_X1  g875(.A1(new_n1076), .A2(G218gat), .ZN(new_n1077));
  OR2_X1    g876(.A1(new_n767), .A2(G218gat), .ZN(new_n1078));
  OAI21_X1  g877(.A(new_n1077), .B1(new_n1065), .B2(new_n1078), .ZN(G1355gat));
endmodule


