//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1142, new_n1143;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT67), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT68), .B(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(G137), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n461), .A2(G101), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  XOR2_X1   g044(.A(KEYINPUT3), .B(G2104), .Z(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT69), .Z(G160));
  NAND2_X1  g052(.A1(new_n463), .A2(new_n465), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n474), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OR3_X1    g057(.A1(KEYINPUT70), .A2(G100), .A3(G2105), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n474), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT70), .B1(G100), .B2(G2105), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n483), .A2(new_n484), .A3(G2104), .A4(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n480), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI21_X1  g063(.A(KEYINPUT71), .B1(new_n474), .B2(G114), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(new_n491), .A3(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n489), .A2(new_n492), .A3(G2104), .A4(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n463), .A2(G126), .A3(G2105), .A4(new_n465), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT3), .B(G2104), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(G138), .A3(new_n474), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT4), .A2(G138), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n463), .A2(new_n474), .A3(new_n465), .A4(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n496), .A2(new_n497), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT75), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT74), .A3(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT73), .B(G651), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n509), .B(new_n511), .C1(new_n512), .C2(new_n510), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n506), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n508), .A2(KEYINPUT73), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT6), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n509), .A2(new_n511), .ZN(new_n525));
  INV_X1    g100(.A(new_n518), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT75), .A4(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G88), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n510), .B1(new_n520), .B2(new_n522), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n509), .A2(new_n511), .ZN(new_n531));
  NOR3_X1   g106(.A1(new_n530), .A2(new_n531), .A3(new_n514), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G50), .ZN(new_n533));
  NAND2_X1  g108(.A1(G75), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G62), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n518), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(new_n512), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT76), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n529), .A2(new_n533), .A3(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  XNOR2_X1  g115(.A(KEYINPUT77), .B(G89), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n528), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n532), .B2(G51), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n542), .A2(new_n544), .A3(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  NAND2_X1  g123(.A1(new_n528), .A2(G90), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT78), .B(G52), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n518), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n532), .A2(new_n550), .B1(new_n512), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n549), .A2(new_n554), .ZN(G171));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n518), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(new_n512), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT79), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n519), .A2(G81), .A3(new_n527), .ZN(new_n561));
  XNOR2_X1  g136(.A(KEYINPUT80), .B(G43), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n532), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT81), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(G188));
  INV_X1    g147(.A(KEYINPUT82), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT9), .B1(new_n532), .B2(G53), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n524), .A2(new_n525), .A3(G53), .A4(G543), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n573), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  XNOR2_X1  g154(.A(KEYINPUT83), .B(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n518), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n519), .A2(G91), .A3(new_n527), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n532), .A2(KEYINPUT9), .A3(G53), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n575), .A2(new_n576), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT82), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n578), .A2(new_n582), .A3(new_n583), .A4(new_n586), .ZN(G299));
  NAND2_X1  g162(.A1(new_n549), .A2(new_n554), .ZN(G301));
  INV_X1    g163(.A(G74), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n508), .B1(new_n518), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n532), .B2(G49), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n519), .A2(new_n527), .ZN(new_n592));
  INV_X1    g167(.A(G87), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(G288));
  AND3_X1   g169(.A1(new_n526), .A2(G61), .A3(new_n512), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n512), .A2(G73), .ZN(new_n596));
  INV_X1    g171(.A(G48), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n513), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n595), .B1(new_n598), .B2(G543), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n519), .A2(G86), .A3(new_n527), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(new_n532), .A2(G47), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  OAI221_X1 g179(.A(new_n602), .B1(new_n523), .B2(new_n603), .C1(new_n592), .C2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n519), .A2(G92), .A3(new_n527), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n519), .A2(KEYINPUT10), .A3(G92), .A4(new_n527), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n532), .A2(G54), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n526), .A2(G66), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n508), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n606), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n606), .B1(new_n618), .B2(G868), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  INV_X1    g196(.A(new_n586), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n583), .A2(new_n582), .ZN(new_n623));
  AOI21_X1  g198(.A(KEYINPUT82), .B1(new_n584), .B2(new_n585), .ZN(new_n624));
  NOR3_X1   g199(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n621), .B1(G868), .B2(new_n625), .ZN(G280));
  XNOR2_X1  g201(.A(G280), .B(KEYINPUT84), .ZN(G297));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n618), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n618), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n479), .A2(G123), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n481), .A2(G135), .ZN(new_n635));
  NOR2_X1   g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(new_n474), .B2(G111), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT85), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n498), .A2(new_n461), .A3(new_n474), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT15), .B(G2435), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2443), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n656), .B(new_n657), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G14), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(new_n666), .A3(KEYINPUT17), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2072), .B(G2078), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n670), .C1(new_n668), .C2(new_n664), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n670), .B2(new_n669), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n676), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  AOI22_X1  g257(.A1(new_n680), .A2(KEYINPUT20), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n682), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n684), .A2(new_n676), .A3(new_n679), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n683), .B(new_n685), .C1(KEYINPUT20), .C2(new_n680), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1986), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1991), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(G229));
  NOR2_X1   g267(.A1(G16), .A2(G24), .ZN(new_n693));
  XNOR2_X1  g268(.A(G290), .B(KEYINPUT88), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1986), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G25), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n479), .A2(G119), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n481), .A2(G131), .ZN(new_n701));
  OR2_X1    g276(.A1(G95), .A2(G2105), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n702), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(new_n698), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT87), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT35), .B(G1991), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n710), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(G1971), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(G6), .ZN(new_n714));
  INV_X1    g289(.A(G305), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n710), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT32), .B(G1981), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n710), .A2(G23), .ZN(new_n719));
  INV_X1    g294(.A(G288), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n710), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT33), .B(G1976), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT90), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n721), .B(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n713), .A2(new_n718), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n709), .B1(new_n725), .B2(KEYINPUT34), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n697), .B(new_n726), .C1(KEYINPUT34), .C2(new_n725), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n728), .A2(KEYINPUT91), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n727), .B(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n698), .A2(G35), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n731), .B(new_n732), .C1(new_n487), .C2(G29), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n731), .B2(new_n732), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT97), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n734), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G2090), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT98), .ZN(new_n739));
  NAND2_X1  g314(.A1(G171), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G5), .B2(G16), .ZN(new_n741));
  INV_X1    g316(.A(G1961), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(KEYINPUT24), .A2(G34), .ZN(new_n744));
  NAND2_X1  g319(.A1(KEYINPUT24), .A2(G34), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n744), .A2(new_n698), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G160), .B2(new_n698), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n481), .A2(G141), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  AND2_X1   g327(.A1(new_n474), .A2(G105), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n479), .A2(G129), .B1(new_n461), .B2(new_n753), .ZN(new_n754));
  AND3_X1   g329(.A1(new_n750), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G29), .B2(G32), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT27), .B(G1996), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n743), .B1(G2084), .B2(new_n747), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT94), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT99), .B(G1956), .Z(new_n761));
  OAI21_X1  g336(.A(KEYINPUT23), .B1(new_n625), .B2(new_n710), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n710), .A2(G20), .ZN(new_n763));
  MUX2_X1   g338(.A(KEYINPUT23), .B(new_n762), .S(new_n763), .Z(new_n764));
  OAI21_X1  g339(.A(new_n760), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n481), .A2(G139), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n498), .A2(G127), .ZN(new_n767));
  AND2_X1   g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(G2105), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT25), .Z(new_n771));
  NAND3_X1  g346(.A1(new_n766), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G33), .B(new_n772), .S(G29), .Z(new_n773));
  AOI22_X1  g348(.A1(new_n757), .A2(new_n758), .B1(G2072), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n747), .A2(G2084), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n774), .B(new_n775), .C1(G2072), .C2(new_n773), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT93), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n710), .A2(G4), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n618), .B2(new_n710), .ZN(new_n779));
  OAI22_X1  g354(.A1(new_n737), .A2(G2090), .B1(G1348), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(G1348), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n742), .B2(new_n741), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n764), .A2(new_n761), .ZN(new_n784));
  NOR2_X1   g359(.A1(G16), .A2(G21), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G168), .B2(G16), .ZN(new_n786));
  INV_X1    g361(.A(G1966), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n698), .A2(G26), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n479), .A2(G128), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n481), .A2(G140), .ZN(new_n791));
  OR2_X1    g366(.A1(G104), .A2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n789), .B1(new_n794), .B2(G29), .ZN(new_n795));
  MUX2_X1   g370(.A(new_n789), .B(new_n795), .S(KEYINPUT28), .Z(new_n796));
  INV_X1    g371(.A(G2067), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G28), .ZN(new_n799));
  AOI21_X1  g374(.A(G29), .B1(new_n799), .B2(KEYINPUT30), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(KEYINPUT30), .B2(new_n799), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n639), .B2(new_n698), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n698), .A2(G27), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G164), .B2(new_n698), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2078), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT31), .B(G11), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n710), .A2(G19), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n565), .B2(new_n710), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1341), .ZN(new_n810));
  NOR4_X1   g385(.A1(new_n798), .A2(new_n806), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n783), .A2(new_n784), .A3(new_n788), .A4(new_n811), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n765), .A2(new_n777), .A3(new_n812), .ZN(new_n813));
  AND3_X1   g388(.A1(new_n730), .A2(new_n739), .A3(new_n813), .ZN(G311));
  NAND3_X1  g389(.A1(new_n730), .A2(new_n739), .A3(new_n813), .ZN(G150));
  NAND2_X1  g390(.A1(G80), .A2(G543), .ZN(new_n816));
  INV_X1    g391(.A(G67), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n518), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(new_n512), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT101), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n519), .A2(G93), .A3(new_n527), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n532), .A2(G55), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n821), .A2(KEYINPUT102), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(KEYINPUT102), .B1(new_n821), .B2(new_n822), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT103), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n618), .A2(G559), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT39), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n825), .A2(new_n565), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n564), .B(new_n820), .C1(new_n823), .C2(new_n824), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n830), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n828), .B1(new_n836), .B2(G860), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT104), .ZN(G145));
  XNOR2_X1  g413(.A(new_n794), .B(new_n504), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(new_n772), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n772), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n755), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n479), .A2(G130), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n481), .A2(G142), .ZN(new_n846));
  NOR2_X1   g421(.A1(G106), .A2(G2105), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(new_n474), .B2(G118), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n845), .B(new_n846), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(new_n642), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n704), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n840), .A2(new_n755), .A3(new_n841), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n844), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(KEYINPUT105), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n639), .B(G160), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n487), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n844), .A2(new_n852), .ZN(new_n858));
  INV_X1    g433(.A(new_n851), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(KEYINPUT105), .A3(new_n853), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n858), .A2(KEYINPUT106), .A3(new_n859), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT106), .B1(new_n858), .B2(new_n859), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n856), .B(new_n853), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(G395));
  INV_X1    g444(.A(KEYINPUT110), .ZN(new_n870));
  XNOR2_X1  g445(.A(G290), .B(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(G288), .B(G305), .Z(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(G166), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n875), .ZN(new_n877));
  OAI21_X1  g452(.A(G303), .B1(new_n877), .B2(new_n873), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT42), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n833), .B(new_n630), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n617), .A2(new_n625), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n615), .B1(new_n609), .B2(new_n610), .ZN(new_n884));
  NAND3_X1  g459(.A1(G299), .A2(new_n884), .A3(new_n612), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(KEYINPUT108), .A3(new_n885), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n618), .A2(new_n888), .A3(G299), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(KEYINPUT41), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n881), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n889), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n881), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT109), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT109), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n880), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n880), .B1(new_n894), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g473(.A(G868), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n825), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n899), .B1(G868), .B2(new_n900), .ZN(G295));
  OAI21_X1  g476(.A(new_n899), .B1(G868), .B2(new_n900), .ZN(G331));
  NAND3_X1  g477(.A1(new_n549), .A2(KEYINPUT111), .A3(new_n554), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n903), .A2(new_n544), .A3(new_n542), .A4(new_n546), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n831), .A2(new_n832), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n831), .B2(new_n832), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT112), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT111), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(G301), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(G301), .A2(new_n908), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n905), .A2(new_n906), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n911), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n914), .A2(new_n909), .ZN(new_n915));
  AOI21_X1  g490(.A(G286), .B1(G171), .B2(KEYINPUT111), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n821), .A2(new_n822), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n821), .A2(KEYINPUT102), .A3(new_n822), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n564), .B1(new_n921), .B2(new_n820), .ZN(new_n922));
  INV_X1    g497(.A(new_n832), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n916), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n831), .A2(new_n832), .A3(new_n904), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n892), .B1(new_n913), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n876), .A2(new_n878), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n890), .A2(new_n886), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n912), .B1(new_n905), .B2(new_n906), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n915), .A3(new_n925), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n866), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT113), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n930), .A2(new_n931), .B1(new_n889), .B2(new_n887), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n879), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n933), .A2(KEYINPUT113), .A3(new_n866), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n936), .A2(new_n937), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n930), .A2(KEYINPUT41), .A3(new_n931), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n892), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n882), .A2(new_n885), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n930), .A2(KEYINPUT41), .A3(new_n931), .A4(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n928), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(new_n940), .A3(new_n866), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n943), .B1(new_n949), .B2(KEYINPUT43), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n942), .A2(new_n950), .A3(KEYINPUT114), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT114), .B1(new_n942), .B2(new_n950), .ZN(new_n952));
  AND4_X1   g527(.A1(new_n937), .A2(new_n948), .A3(new_n940), .A4(new_n866), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n936), .A2(new_n940), .A3(new_n941), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(KEYINPUT43), .ZN(new_n955));
  OAI22_X1  g530(.A1(new_n951), .A2(new_n952), .B1(KEYINPUT44), .B2(new_n955), .ZN(G397));
  XNOR2_X1  g531(.A(new_n755), .B(G1996), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n794), .B(new_n797), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n704), .B(new_n708), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT115), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(G290), .B(G1986), .Z(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n504), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G40), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n468), .A2(new_n475), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n964), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G8), .ZN(new_n974));
  INV_X1    g549(.A(new_n475), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n468), .A2(new_n969), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n968), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n787), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n966), .A2(KEYINPUT50), .ZN(new_n980));
  INV_X1    g555(.A(G2084), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n504), .A2(new_n982), .A3(new_n965), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n980), .A2(new_n970), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n974), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(KEYINPUT118), .B(G8), .Z(new_n986));
  NAND2_X1  g561(.A1(G286), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT51), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n990));
  INV_X1    g565(.A(new_n986), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n979), .B2(new_n984), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n990), .B1(new_n992), .B2(KEYINPUT125), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n468), .A2(new_n969), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n966), .B2(new_n967), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n977), .A2(new_n975), .ZN(new_n996));
  AOI21_X1  g571(.A(G1966), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n984), .ZN(new_n998));
  OAI211_X1 g573(.A(KEYINPUT125), .B(new_n986), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n987), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n989), .B1(new_n993), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT62), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n988), .B1(new_n997), .B2(new_n998), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G303), .A2(G8), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n977), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n504), .A2(KEYINPUT116), .A3(KEYINPUT45), .A4(new_n965), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n995), .A2(new_n1009), .A3(new_n975), .A4(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT117), .B(G1971), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n980), .A2(new_n970), .A3(new_n983), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(G2090), .ZN(new_n1015));
  OAI211_X1 g590(.A(G8), .B(new_n1007), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1007), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1014), .ZN(new_n1018));
  INV_X1    g593(.A(G2090), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1011), .A2(new_n1012), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1017), .B1(new_n1020), .B2(new_n991), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n986), .B1(new_n971), .B2(new_n966), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT49), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G305), .A2(G1981), .ZN(new_n1024));
  INV_X1    g599(.A(G1981), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n599), .B2(new_n600), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1023), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT119), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1029), .B(new_n1023), .C1(new_n1024), .C2(new_n1026), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1022), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  OR3_X1    g606(.A1(new_n1024), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1032));
  INV_X1    g607(.A(G1976), .ZN(new_n1033));
  OAI221_X1 g608(.A(new_n986), .B1(G288), .B2(new_n1033), .C1(new_n971), .C2(new_n966), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1031), .A2(new_n1032), .B1(KEYINPUT52), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n720), .A2(G1976), .ZN(new_n1036));
  OR3_X1    g611(.A1(new_n1034), .A2(KEYINPUT52), .A3(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1016), .A2(new_n1021), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G2078), .ZN(new_n1040));
  AND4_X1   g615(.A1(new_n1040), .A2(new_n995), .A3(new_n1010), .A4(new_n1009), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT53), .B1(new_n1041), .B2(new_n975), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(new_n742), .B2(new_n1014), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n995), .A2(new_n996), .A3(KEYINPUT53), .A4(new_n1040), .ZN(new_n1044));
  AOI21_X1  g619(.A(G301), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1004), .A2(new_n1039), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT127), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT62), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT127), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1004), .A2(new_n1039), .A3(new_n1050), .A4(new_n1045), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1047), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1020), .A2(new_n974), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1007), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n1033), .A3(new_n720), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1024), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1022), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT120), .B(KEYINPUT63), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n992), .A2(G168), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1038), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT63), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1017), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1063), .B1(new_n1065), .B2(new_n1054), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1061), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1017), .B(new_n1064), .C1(new_n1020), .C2(new_n974), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1053), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1059), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT56), .B(G2072), .Z(new_n1071));
  OAI22_X1  g646(.A1(new_n1011), .A2(new_n1071), .B1(new_n1018), .B2(G1956), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n584), .A2(new_n585), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(new_n623), .B2(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1075), .A2(KEYINPUT122), .ZN(new_n1076));
  NOR2_X1   g651(.A1(G299), .A2(new_n1073), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1075), .A2(KEYINPUT122), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1072), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1348), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n970), .A2(new_n965), .A3(new_n504), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1014), .A2(new_n1081), .B1(new_n1082), .B2(new_n797), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n617), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n1085));
  OR3_X1    g660(.A1(new_n1072), .A2(new_n1079), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1085), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1083), .A2(new_n617), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1083), .A2(new_n617), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT60), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1083), .A2(new_n1092), .A3(new_n618), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT58), .B(G1341), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n1011), .A2(G1996), .B1(new_n1082), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(KEYINPUT124), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1095), .A2(new_n565), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1095), .B2(new_n565), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1091), .B(new_n1093), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT61), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1086), .A2(new_n1080), .A3(new_n1087), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1088), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1109));
  XNOR2_X1  g684(.A(G171), .B(KEYINPUT54), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n472), .A2(KEYINPUT126), .ZN(new_n1113));
  OAI21_X1  g688(.A(G2105), .B1(new_n472), .B2(KEYINPUT126), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1041), .B(KEYINPUT53), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1043), .A2(new_n1110), .A3(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1112), .A2(new_n1039), .A3(new_n1048), .A4(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1055), .B(new_n1070), .C1(new_n1108), .C2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n973), .B1(new_n1052), .B2(new_n1118), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n959), .A2(new_n708), .A3(new_n704), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n794), .A2(G2067), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n972), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n972), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1123), .A2(G1986), .A3(G290), .ZN(new_n1124));
  XOR2_X1   g699(.A(new_n1124), .B(KEYINPUT48), .Z(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n962), .B2(new_n1123), .ZN(new_n1126));
  INV_X1    g701(.A(new_n958), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n972), .B1(new_n843), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT46), .ZN(new_n1129));
  OR3_X1    g704(.A1(new_n1123), .A2(new_n1129), .A3(G1996), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1123), .B2(G1996), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT47), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1122), .A2(new_n1126), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1119), .A2(new_n1134), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g710(.A1(G401), .A2(G227), .ZN(new_n1137));
  NAND2_X1  g711(.A1(new_n867), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g712(.A1(G229), .A2(new_n459), .ZN(new_n1139));
  INV_X1    g713(.A(new_n1139), .ZN(new_n1140));
  NOR3_X1   g714(.A1(new_n955), .A2(new_n1138), .A3(new_n1140), .ZN(G308));
  AND2_X1   g715(.A1(new_n867), .A2(new_n1137), .ZN(new_n1142));
  AND2_X1   g716(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n1143));
  OAI211_X1 g717(.A(new_n1142), .B(new_n1139), .C1(new_n1143), .C2(new_n953), .ZN(G225));
endmodule


