//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  XOR2_X1   g000(.A(G155gat), .B(G162gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT77), .B(G148gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G141gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n202), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n209), .B1(G155gat), .B2(G162gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT78), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G141gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G148gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n209), .B1(new_n206), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n202), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n208), .A2(new_n211), .B1(new_n202), .B2(new_n215), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(G127gat), .B(G134gat), .Z(new_n222));
  XNOR2_X1  g021(.A(G113gat), .B(G120gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G113gat), .B(G120gat), .Z(new_n225));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n226));
  XNOR2_X1  g025(.A(G127gat), .B(G134gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n228), .A3(KEYINPUT79), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT79), .B1(new_n224), .B2(new_n228), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n218), .A2(new_n221), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G225gat), .A2(G233gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n224), .A2(new_n228), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n219), .A2(new_n236), .A3(KEYINPUT4), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n233), .A2(new_n234), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT5), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT79), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n229), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n237), .B1(new_n245), .B2(new_n219), .ZN(new_n246));
  INV_X1    g045(.A(new_n234), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n242), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n245), .B1(KEYINPUT3), .B2(new_n217), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n249), .B2(new_n221), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n237), .A2(new_n238), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT4), .B1(new_n219), .B2(new_n236), .ZN(new_n252));
  NOR3_X1   g051(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT5), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n241), .A2(new_n248), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G1gat), .B(G29gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT0), .ZN(new_n256));
  XNOR2_X1  g055(.A(G57gat), .B(G85gat), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n256), .B(new_n257), .Z(new_n258));
  AOI21_X1  g057(.A(KEYINPUT6), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT85), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n259), .B(new_n260), .C1(new_n258), .C2(new_n254), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n248), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n250), .A2(new_n253), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n263), .A3(new_n258), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT6), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n254), .A2(new_n258), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT85), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(KEYINPUT6), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n261), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(G226gat), .A2(G233gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(G183gat), .A2(G190gat), .ZN(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(KEYINPUT26), .ZN(new_n278));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT26), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OR2_X1    g081(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n287), .A2(KEYINPUT27), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT27), .B(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT70), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT28), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n291), .A2(new_n285), .A3(new_n294), .ZN(new_n295));
  OAI221_X1 g094(.A(new_n274), .B1(new_n278), .B2(new_n282), .C1(new_n293), .C2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n297));
  AND2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n280), .A2(KEYINPUT23), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT67), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n300), .A2(new_n301), .A3(new_n305), .A4(new_n302), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT25), .B1(new_n280), .B2(KEYINPUT23), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n283), .A2(new_n287), .A3(new_n284), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n274), .A2(KEYINPUT24), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT24), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(G183gat), .A3(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n308), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT25), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n298), .B1(new_n277), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(G169gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n276), .A2(KEYINPUT64), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT64), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G176gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n324), .B1(new_n310), .B2(new_n312), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n315), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT65), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(KEYINPUT65), .B(new_n315), .C1(new_n323), .C2(new_n325), .ZN(new_n329));
  AOI221_X4 g128(.A(new_n297), .B1(new_n307), .B2(new_n314), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n329), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n307), .A2(new_n314), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT69), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n273), .B(new_n296), .C1(new_n330), .C2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n329), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n287), .A2(KEYINPUT24), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n336), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n274), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n322), .B(new_n317), .C1(new_n337), .C2(new_n324), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT65), .B1(new_n338), .B2(new_n315), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n332), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n296), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n273), .A2(KEYINPUT29), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n334), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G197gat), .B(G204gat), .ZN(new_n345));
  INV_X1    g144(.A(G211gat), .ZN(new_n346));
  INV_X1    g145(.A(G218gat), .ZN(new_n347));
  OAI22_X1  g146(.A1(new_n346), .A2(new_n347), .B1(KEYINPUT73), .B2(KEYINPUT22), .ZN(new_n348));
  AND2_X1   g147(.A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G211gat), .B(G218gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT74), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n344), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n353), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n296), .A3(new_n273), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n293), .A2(new_n295), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n274), .B1(new_n278), .B2(new_n282), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n297), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n331), .A2(KEYINPUT69), .A3(new_n332), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n342), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n355), .B(new_n356), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n365));
  NAND3_X1  g164(.A1(new_n354), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT37), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n372), .B1(new_n354), .B2(new_n364), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n272), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n362), .A2(new_n273), .B1(new_n342), .B2(new_n341), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n364), .B(new_n369), .C1(new_n375), .C2(new_n355), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT75), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT75), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n354), .A2(new_n378), .A3(new_n364), .A4(new_n369), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n353), .B(new_n356), .C1(new_n362), .C2(new_n363), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n381), .B(KEYINPUT37), .C1(new_n375), .C2(new_n353), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n366), .A2(new_n382), .A3(new_n370), .A4(new_n271), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n270), .A2(new_n374), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n220), .B1(new_n352), .B2(KEYINPUT29), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n217), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n219), .B2(new_n220), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n386), .B1(new_n353), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT83), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n388), .B(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G228gat), .A2(G233gat), .ZN(new_n392));
  INV_X1    g191(.A(G22gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT31), .B(G50gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n391), .B(new_n396), .Z(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(KEYINPUT76), .B(KEYINPUT30), .Z(new_n399));
  NAND3_X1  g198(.A1(new_n377), .A2(new_n379), .A3(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n340), .A2(new_n296), .A3(new_n273), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n296), .B1(new_n330), .B2(new_n333), .ZN(new_n402));
  AOI211_X1 g201(.A(new_n353), .B(new_n401), .C1(new_n402), .C2(new_n342), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n355), .B1(new_n334), .B2(new_n343), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n370), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n354), .A2(KEYINPUT30), .A3(new_n364), .A4(new_n369), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT84), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n400), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n251), .A2(new_n252), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n233), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n247), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n415), .B(KEYINPUT39), .C1(new_n247), .C2(new_n246), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n416), .B(new_n258), .C1(KEYINPUT39), .C2(new_n415), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT40), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n267), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n418), .B2(new_n417), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n384), .B(new_n398), .C1(new_n412), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n402), .A2(new_n235), .ZN(new_n422));
  NAND2_X1  g221(.A1(G227gat), .A2(G233gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n360), .A2(new_n361), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(new_n296), .A3(new_n236), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT34), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT34), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n422), .A2(new_n425), .A3(new_n428), .A4(new_n423), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G71gat), .B(G99gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT71), .ZN(new_n432));
  INV_X1    g231(.A(G15gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G43gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n423), .B1(new_n422), .B2(new_n425), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(KEYINPUT33), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT32), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n423), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n236), .B1(new_n424), .B2(new_n296), .ZN(new_n443));
  AOI211_X1 g242(.A(new_n359), .B(new_n235), .C1(new_n360), .C2(new_n361), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446));
  INV_X1    g245(.A(new_n436), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n445), .B(KEYINPUT32), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n430), .B1(new_n441), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT72), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n427), .A2(new_n429), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n445), .A2(KEYINPUT32), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n445), .A2(new_n446), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n436), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n456), .B2(new_n448), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT72), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n453), .A3(new_n448), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n452), .A2(new_n458), .A3(KEYINPUT36), .A4(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT36), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n456), .A2(new_n453), .A3(new_n448), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n461), .B1(new_n462), .B2(new_n457), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT81), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(new_n254), .B2(new_n258), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n262), .A2(new_n263), .ZN(new_n467));
  INV_X1    g266(.A(new_n258), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(KEYINPUT81), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n266), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n269), .B1(new_n470), .B2(KEYINPUT82), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n254), .A2(new_n465), .A3(new_n258), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT81), .B1(new_n467), .B2(new_n468), .ZN(new_n473));
  OAI211_X1 g272(.A(KEYINPUT82), .B(new_n259), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n397), .B1(new_n476), .B2(new_n408), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n421), .A2(new_n464), .A3(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n270), .A2(new_n397), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n450), .A2(KEYINPUT88), .A3(new_n459), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT88), .B1(new_n450), .B2(new_n459), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n412), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT35), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI211_X1 g283(.A(new_n451), .B(new_n453), .C1(new_n456), .C2(new_n448), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n456), .A2(new_n448), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT72), .B1(new_n486), .B2(new_n430), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n459), .A2(new_n398), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n476), .A2(new_n483), .A3(new_n408), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n478), .A2(new_n484), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G29gat), .A2(G36gat), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NOR3_X1   g294(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(KEYINPUT15), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(KEYINPUT15), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT15), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n435), .A2(G50gat), .ZN(new_n502));
  INV_X1    g301(.A(G50gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(G43gat), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n501), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n500), .A2(new_n505), .A3(new_n493), .ZN(new_n506));
  NOR2_X1   g305(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n507));
  INV_X1    g306(.A(G36gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT90), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n495), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n499), .B(KEYINPUT17), .C1(new_n506), .C2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT92), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n433), .A2(new_n393), .ZN(new_n516));
  NAND2_X1  g315(.A1(G15gat), .A2(G22gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(G1gat), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G8gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT92), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G1gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT16), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n516), .B2(new_n517), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n515), .B(G8gat), .C1(new_n521), .C2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n524), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n515), .A2(G8gat), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n526), .A2(new_n527), .A3(new_n520), .A4(new_n518), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n514), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n499), .B1(new_n506), .B2(new_n513), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n531), .A2(KEYINPUT91), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT91), .B1(new_n531), .B2(new_n532), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n525), .A2(new_n528), .A3(KEYINPUT93), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT93), .B1(new_n525), .B2(new_n528), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n531), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n535), .A2(KEYINPUT18), .A3(new_n536), .A4(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n535), .A2(new_n536), .A3(new_n540), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT18), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n536), .B(KEYINPUT13), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT93), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n531), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n549), .A3(new_n537), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n546), .B1(new_n540), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT89), .B(G197gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT11), .B(G169gat), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT12), .ZN(new_n558));
  AND4_X1   g357(.A1(new_n541), .A2(new_n544), .A3(new_n552), .A4(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n551), .B1(new_n542), .B2(new_n543), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n558), .B1(new_n560), .B2(new_n541), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n492), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n565));
  INV_X1    g364(.A(G57gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(G64gat), .ZN(new_n567));
  INV_X1    g366(.A(G64gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G57gat), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n565), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT94), .ZN(new_n571));
  AND2_X1   g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(KEYINPUT94), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n570), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n576), .ZN(new_n579));
  XNOR2_X1  g378(.A(G57gat), .B(G64gat), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n579), .B(new_n571), .C1(new_n580), .C2(new_n565), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  OR2_X1    g384(.A1(new_n585), .A2(G127gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(G127gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n578), .A2(new_n581), .ZN(new_n589));
  AOI211_X1 g388(.A(new_n539), .B(new_n538), .C1(KEYINPUT21), .C2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n588), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n593));
  INV_X1    g392(.A(G155gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n592), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n601));
  AND2_X1   g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT96), .ZN(new_n604));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n606), .B(KEYINPUT97), .Z(new_n607));
  XNOR2_X1  g406(.A(G99gat), .B(G106gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(G85gat), .A2(G92gat), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT7), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT8), .ZN(new_n615));
  INV_X1    g414(.A(G85gat), .ZN(new_n616));
  INV_X1    g415(.A(G92gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n608), .B1(new_n613), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n615), .A2(new_n611), .A3(new_n618), .A4(new_n612), .ZN(new_n621));
  INV_X1    g420(.A(new_n608), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n531), .A2(new_n624), .B1(KEYINPUT41), .B2(new_n602), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT99), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT98), .B1(new_n620), .B2(new_n623), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n619), .A2(new_n613), .A3(new_n608), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n621), .A2(new_n622), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n514), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n533), .B2(new_n534), .ZN(new_n634));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT100), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n626), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n626), .B2(new_n634), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n601), .B(new_n607), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n636), .ZN(new_n640));
  INV_X1    g439(.A(new_n634), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n625), .B(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n640), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n626), .A2(new_n634), .A3(new_n636), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n645), .A3(new_n606), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n601), .B1(new_n648), .B2(new_n607), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n600), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n581), .B(new_n578), .C1(new_n620), .C2(new_n623), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n589), .A2(new_n628), .A3(new_n630), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT10), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n589), .A2(KEYINPUT10), .A3(new_n628), .A4(new_n630), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n624), .A2(KEYINPUT102), .A3(KEYINPUT10), .A4(new_n589), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n659), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(G230gat), .A2(G233gat), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n665), .B1(new_n656), .B2(new_n657), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT103), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n655), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI211_X1 g471(.A(KEYINPUT104), .B(new_n654), .C1(new_n667), .C2(new_n669), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n651), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n564), .A2(new_n476), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  INV_X1    g477(.A(new_n412), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n564), .A2(new_n679), .A3(new_n676), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  AND2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(new_n519), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(KEYINPUT42), .B2(new_n682), .ZN(G1325gat));
  NOR2_X1   g484(.A1(new_n480), .A2(new_n481), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n564), .A2(new_n433), .A3(new_n687), .A4(new_n676), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n564), .A2(new_n676), .ZN(new_n689));
  INV_X1    g488(.A(new_n464), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n688), .B1(new_n691), .B2(new_n433), .ZN(G1326gat));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n397), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT43), .B(G22gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  NOR2_X1   g494(.A1(new_n600), .A2(new_n650), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n674), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n564), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n476), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n699), .A2(G29gat), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT45), .Z(new_n702));
  AND3_X1   g501(.A1(new_n598), .A2(KEYINPUT105), .A3(new_n599), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT105), .B1(new_n598), .B2(new_n599), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n675), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n563), .ZN(new_n708));
  AOI221_X4 g507(.A(KEYINPUT106), .B1(new_n489), .B2(new_n490), .C1(new_n482), .C2(new_n483), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n484), .B2(new_n491), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n478), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n713));
  NOR2_X1   g512(.A1(new_n650), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n648), .A2(new_n607), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT101), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n646), .A3(new_n639), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n716), .B1(new_n492), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n708), .B1(new_n715), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n700), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n702), .A2(new_n724), .ZN(G1328gat));
  NOR3_X1   g524(.A1(new_n699), .A2(G36gat), .A3(new_n412), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT46), .ZN(new_n727));
  OAI21_X1  g526(.A(G36gat), .B1(new_n723), .B2(new_n412), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1329gat));
  INV_X1    g528(.A(new_n708), .ZN(new_n730));
  INV_X1    g529(.A(new_n714), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT88), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n462), .B2(new_n457), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n450), .A2(KEYINPUT88), .A3(new_n459), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n733), .A2(new_n734), .B1(new_n409), .B2(new_n411), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT35), .B1(new_n735), .B2(new_n479), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n489), .A2(new_n490), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT106), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n484), .A2(new_n710), .A3(new_n491), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n731), .B1(new_n740), .B2(new_n478), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n690), .B(new_n730), .C1(new_n741), .C2(new_n720), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G43gat), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT47), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n564), .A2(new_n435), .A3(new_n687), .A4(new_n698), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n743), .B(new_n746), .C1(new_n744), .C2(KEYINPUT47), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1330gat));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n503), .B1(new_n722), .B2(new_n397), .ZN(new_n752));
  AND4_X1   g551(.A1(new_n503), .A2(new_n564), .A3(new_n397), .A4(new_n698), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n751), .B(KEYINPUT48), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n397), .B(new_n730), .C1(new_n741), .C2(new_n720), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n753), .B1(new_n756), .B2(G50gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n757), .B2(KEYINPUT109), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n754), .A2(new_n758), .ZN(G1331gat));
  AOI21_X1  g558(.A(new_n563), .B1(new_n740), .B2(new_n478), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n651), .A2(new_n674), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n700), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(new_n566), .ZN(G1332gat));
  INV_X1    g563(.A(new_n762), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n679), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT49), .B(G64gat), .Z(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(G1333gat));
  NAND3_X1  g568(.A1(new_n765), .A2(G71gat), .A3(new_n690), .ZN(new_n770));
  INV_X1    g569(.A(G71gat), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n687), .A2(KEYINPUT110), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n686), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n771), .B1(new_n762), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n770), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n770), .B2(new_n776), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(G1334gat));
  NOR2_X1   g579(.A1(new_n762), .A2(new_n398), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT112), .B(G78gat), .Z(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1335gat));
  NAND2_X1  g582(.A1(new_n715), .A2(new_n721), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n600), .A2(new_n563), .A3(new_n674), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT113), .B1(new_n786), .B2(new_n700), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G85gat), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n786), .A2(KEYINPUT113), .A3(new_n700), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n712), .A2(new_n562), .A3(new_n696), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT51), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n760), .A2(new_n792), .A3(new_n696), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(new_n793), .A3(new_n675), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n476), .A2(new_n616), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n788), .A2(new_n789), .B1(new_n794), .B2(new_n795), .ZN(G1336gat));
  OAI211_X1 g595(.A(new_n679), .B(new_n785), .C1(new_n741), .C2(new_n720), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G92gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n679), .A2(new_n617), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT52), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n798), .B(new_n802), .C1(new_n794), .C2(new_n799), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(G1337gat));
  OAI21_X1  g603(.A(G99gat), .B1(new_n786), .B2(new_n464), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n686), .A2(G99gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n794), .B2(new_n806), .ZN(G1338gat));
  OAI211_X1 g606(.A(new_n397), .B(new_n785), .C1(new_n741), .C2(new_n720), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G106gat), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n398), .A2(G106gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n794), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT53), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n809), .B(new_n813), .C1(new_n794), .C2(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1339gat));
  NAND2_X1  g614(.A1(new_n676), .A2(new_n562), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n560), .A2(new_n541), .A3(new_n558), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n536), .B1(new_n535), .B2(new_n540), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n540), .A2(new_n550), .A3(new_n546), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n557), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n665), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n659), .A2(new_n662), .A3(new_n663), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n666), .A2(KEYINPUT54), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n664), .A2(new_n825), .A3(new_n665), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n655), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n670), .A2(new_n654), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n655), .A4(new_n826), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n650), .A2(new_n821), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n672), .A2(new_n817), .A3(new_n673), .A4(new_n820), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n562), .B2(new_n832), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n719), .B1(new_n835), .B2(KEYINPUT114), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n837), .B(new_n834), .C1(new_n562), .C2(new_n832), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n833), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n705), .B1(new_n839), .B2(KEYINPUT115), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n841));
  AOI211_X1 g640(.A(new_n841), .B(new_n833), .C1(new_n836), .C2(new_n838), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n816), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n489), .ZN(new_n845));
  NOR4_X1   g644(.A1(new_n844), .A2(new_n679), .A3(new_n700), .A4(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n563), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n735), .A2(new_n476), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n844), .B2(new_n397), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n843), .A2(new_n850), .A3(new_n398), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n848), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n563), .A2(G113gat), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n847), .B1(new_n852), .B2(new_n853), .ZN(G1340gat));
  AOI21_X1  g653(.A(G120gat), .B1(new_n846), .B2(new_n675), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n675), .A2(G120gat), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n852), .B2(new_n856), .ZN(G1341gat));
  AND2_X1   g656(.A1(new_n846), .A2(new_n600), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n858), .A2(KEYINPUT117), .ZN(new_n859));
  AOI21_X1  g658(.A(G127gat), .B1(new_n858), .B2(KEYINPUT117), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n706), .A2(G127gat), .ZN(new_n861));
  AOI22_X1  g660(.A1(new_n859), .A2(new_n860), .B1(new_n852), .B2(new_n861), .ZN(G1342gat));
  NOR2_X1   g661(.A1(new_n844), .A2(new_n700), .ZN(new_n863));
  INV_X1    g662(.A(G134gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n412), .A2(new_n719), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT118), .Z(new_n866));
  NAND4_X1  g665(.A1(new_n863), .A2(new_n864), .A3(new_n489), .A4(new_n866), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT56), .Z(new_n868));
  AND2_X1   g667(.A1(new_n852), .A2(new_n719), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n864), .B2(new_n869), .ZN(G1343gat));
  NOR3_X1   g669(.A1(new_n690), .A2(new_n679), .A3(new_n700), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n562), .A2(new_n213), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT57), .B1(new_n843), .B2(new_n397), .ZN(new_n873));
  INV_X1    g672(.A(new_n827), .ZN(new_n874));
  XNOR2_X1  g673(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n830), .B(new_n831), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n834), .B1(new_n876), .B2(new_n562), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n719), .B1(new_n877), .B2(KEYINPUT120), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n878), .B1(KEYINPUT120), .B2(new_n877), .ZN(new_n879));
  INV_X1    g678(.A(new_n833), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n600), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n881), .A2(new_n882), .B1(new_n562), .B2(new_n676), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n397), .A2(KEYINPUT57), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n871), .B(new_n872), .C1(new_n873), .C2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n398), .B1(new_n460), .B2(new_n463), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n843), .A2(new_n412), .A3(new_n476), .A4(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n213), .B1(new_n889), .B2(new_n562), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n887), .A2(KEYINPUT58), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n887), .A2(new_n890), .A3(KEYINPUT121), .A4(KEYINPUT58), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n887), .A2(new_n890), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI211_X1 g698(.A(KEYINPUT122), .B(KEYINPUT58), .C1(new_n887), .C2(new_n890), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n893), .A2(new_n895), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n891), .A2(new_n892), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n894), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n905), .B(KEYINPUT123), .C1(new_n899), .C2(new_n900), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(new_n906), .ZN(G1344gat));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n883), .A2(new_n398), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(KEYINPUT57), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n844), .A2(new_n885), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n871), .A2(new_n675), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n912), .A2(KEYINPUT124), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(new_n205), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT124), .B1(new_n912), .B2(new_n913), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n908), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n873), .A2(new_n886), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(new_n871), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT59), .B(new_n203), .C1(new_n919), .C2(new_n675), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n675), .A2(new_n203), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n917), .A2(new_n920), .B1(new_n889), .B2(new_n921), .ZN(G1345gat));
  AOI21_X1  g721(.A(new_n594), .B1(new_n919), .B2(new_n706), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n889), .A2(G155gat), .A3(new_n882), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n923), .A2(new_n924), .ZN(G1346gat));
  INV_X1    g724(.A(G162gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n926), .B1(new_n919), .B2(new_n719), .ZN(new_n927));
  AND4_X1   g726(.A1(new_n926), .A2(new_n863), .A3(new_n866), .A4(new_n888), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n927), .A2(new_n928), .ZN(G1347gat));
  NOR2_X1   g728(.A1(new_n412), .A2(new_n476), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n844), .A2(new_n845), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n563), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n930), .B1(new_n772), .B2(new_n774), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n934), .A2(KEYINPUT125), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(KEYINPUT125), .ZN(new_n936));
  AOI22_X1  g735(.A1(new_n935), .A2(new_n936), .B1(new_n851), .B2(new_n849), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n562), .A2(new_n275), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n933), .B1(new_n937), .B2(new_n938), .ZN(G1348gat));
  AOI21_X1  g738(.A(G176gat), .B1(new_n932), .B2(new_n675), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n674), .B1(new_n319), .B2(new_n321), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n937), .B2(new_n941), .ZN(G1349gat));
  AOI21_X1  g741(.A(new_n287), .B1(new_n937), .B2(new_n706), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n932), .A2(new_n290), .A3(new_n600), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  OR3_X1    g746(.A1(new_n943), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n943), .B2(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1350gat));
  NAND2_X1  g749(.A1(new_n937), .A2(new_n719), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G190gat), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n951), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n932), .A2(new_n283), .A3(new_n284), .A4(new_n719), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n956), .B(KEYINPUT127), .Z(new_n957));
  NAND3_X1  g756(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(G1351gat));
  NOR2_X1   g757(.A1(new_n690), .A2(new_n931), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n960), .A2(new_n844), .A3(new_n398), .ZN(new_n961));
  AOI21_X1  g760(.A(G197gat), .B1(new_n961), .B2(new_n563), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n912), .A2(new_n960), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n563), .A2(G197gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(G1352gat));
  INV_X1    g764(.A(new_n963), .ZN(new_n966));
  OAI21_X1  g765(.A(G204gat), .B1(new_n966), .B2(new_n674), .ZN(new_n967));
  INV_X1    g766(.A(G204gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n961), .A2(new_n968), .A3(new_n675), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT62), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n969), .A2(KEYINPUT62), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n967), .A2(new_n970), .A3(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n961), .A2(new_n346), .A3(new_n600), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n963), .A2(new_n600), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n974), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  OAI21_X1  g776(.A(G218gat), .B1(new_n966), .B2(new_n650), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n961), .A2(new_n347), .A3(new_n719), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1355gat));
endmodule


