//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT64), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n206), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT0), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n203), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(new_n216), .A2(new_n217), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n223), .B1(new_n217), .B2(new_n216), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n214), .A2(new_n224), .ZN(G361));
  XOR2_X1   g0025(.A(G226), .B(G232), .Z(new_n226));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(G50), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G68), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n202), .A2(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n237), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G1), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G20), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n220), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n245), .A2(G13), .A3(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n247), .A2(new_n252), .A3(new_n238), .ZN(new_n253));
  INV_X1    g0053(.A(new_n251), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n253), .B1(new_n238), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT66), .B1(new_n201), .B2(KEYINPUT8), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT66), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(new_n257), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n221), .A2(G33), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT67), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n264));
  INV_X1    g0064(.A(G150), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n249), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n255), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT71), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(KEYINPUT9), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(KEYINPUT9), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n272), .B(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n245), .B1(G41), .B2(G45), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(G1), .B(G13), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n280), .A2(new_n275), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n281), .A2(G226), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n288), .A2(G223), .B1(G77), .B2(new_n286), .ZN(new_n289));
  INV_X1    g0089(.A(G222), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT3), .B(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n287), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n277), .B(new_n282), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G200), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(G190), .B2(new_n295), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n274), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n270), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(new_n295), .B2(G169), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n295), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n288), .A2(G226), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n286), .A2(G1698), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G223), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G87), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT74), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT74), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n307), .A2(new_n309), .A3(new_n313), .A4(new_n310), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(new_n314), .A3(new_n294), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n277), .B1(new_n281), .B2(G232), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G200), .ZN(new_n318));
  XNOR2_X1  g0118(.A(G58), .B(G68), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(G20), .B1(G159), .B2(new_n266), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT7), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(new_n291), .B2(G20), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n320), .B1(new_n324), .B2(new_n202), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT16), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n250), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n326), .B2(new_n325), .ZN(new_n328));
  INV_X1    g0128(.A(new_n260), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n329), .A2(new_n252), .A3(new_n247), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n254), .B2(new_n329), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n315), .A2(G190), .A3(new_n316), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n318), .A2(new_n328), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT17), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n317), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n315), .A2(new_n304), .A3(new_n316), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(KEYINPUT75), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT75), .ZN(new_n340));
  INV_X1    g0140(.A(new_n316), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n280), .B1(new_n311), .B2(KEYINPUT74), .ZN(new_n342));
  AOI211_X1 g0142(.A(G179), .B(new_n341), .C1(new_n342), .C2(new_n314), .ZN(new_n343));
  AOI21_X1  g0143(.A(G169), .B1(new_n315), .B2(new_n316), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n328), .A2(new_n331), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT18), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n347), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n339), .B2(new_n345), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT18), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n335), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n277), .B1(new_n281), .B2(G238), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n308), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n288), .A2(G232), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n355), .B1(new_n358), .B2(new_n280), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT13), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n359), .B(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT14), .B1(new_n361), .B2(new_n336), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n359), .B(KEYINPUT13), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(G169), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(G179), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n262), .A2(G77), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n266), .A2(G50), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(KEYINPUT72), .B1(G20), .B2(new_n202), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(KEYINPUT72), .B2(new_n369), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n249), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT11), .ZN(new_n373));
  XOR2_X1   g0173(.A(KEYINPUT73), .B(KEYINPUT12), .Z(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n251), .B(KEYINPUT70), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(KEYINPUT12), .B2(new_n251), .ZN(new_n378));
  INV_X1    g0178(.A(new_n376), .ZN(new_n379));
  OR3_X1    g0179(.A1(new_n379), .A2(new_n249), .A3(new_n247), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n375), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G68), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n373), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n367), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n383), .B1(new_n361), .B2(G190), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n363), .A2(G200), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G20), .A2(G77), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT15), .B(G87), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT8), .B(G58), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n389), .B1(new_n390), .B2(new_n261), .C1(new_n267), .C2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G77), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n392), .A2(new_n249), .B1(new_n379), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n380), .B2(new_n393), .ZN(new_n395));
  AND2_X1   g0195(.A1(KEYINPUT69), .A2(G107), .ZN(new_n396));
  NOR2_X1   g0196(.A1(KEYINPUT69), .A2(G107), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n286), .A2(new_n399), .B1(new_n288), .B2(G238), .ZN(new_n400));
  INV_X1    g0200(.A(G232), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(new_n292), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n294), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n277), .B1(new_n281), .B2(G244), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G190), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI211_X1 g0207(.A(new_n395), .B(new_n407), .C1(G200), .C2(new_n405), .ZN(new_n408));
  INV_X1    g0208(.A(new_n405), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n395), .B1(new_n409), .B2(G169), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n405), .A2(G179), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n306), .A2(new_n354), .A3(new_n388), .A4(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G116), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n278), .A2(new_n415), .A3(G20), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n221), .A2(KEYINPUT23), .A3(G107), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n398), .A2(G20), .ZN(new_n418));
  AOI211_X1 g0218(.A(new_n416), .B(new_n417), .C1(new_n418), .C2(KEYINPUT23), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n291), .A2(new_n221), .A3(G87), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT22), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT24), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n250), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n423), .B2(new_n422), .ZN(new_n425));
  XOR2_X1   g0225(.A(KEYINPUT84), .B(KEYINPUT25), .Z(new_n426));
  NOR2_X1   g0226(.A1(new_n251), .A2(G107), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n245), .A2(G33), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n251), .A2(new_n429), .A3(new_n220), .A4(new_n248), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n428), .B1(G107), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n291), .A2(G257), .A3(G1698), .ZN(new_n435));
  INV_X1    g0235(.A(G294), .ZN(new_n436));
  INV_X1    g0236(.A(G250), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n435), .B1(new_n278), .B2(new_n436), .C1(new_n292), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n294), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT5), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n440), .A2(KEYINPUT78), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(KEYINPUT78), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n279), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G45), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(G1), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT76), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n440), .A2(G41), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n245), .B(G45), .C1(new_n279), .C2(KEYINPUT5), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT76), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n443), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(G264), .A3(new_n280), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n439), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT85), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n455));
  OAI211_X1 g0255(.A(G274), .B(new_n280), .C1(new_n455), .C2(G41), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n450), .A2(KEYINPUT77), .A3(new_n448), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT77), .B1(new_n450), .B2(new_n448), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT85), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n439), .A2(new_n461), .A3(new_n452), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n454), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT86), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n296), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT77), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n449), .A2(KEYINPUT76), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n446), .B1(new_n445), .B2(new_n447), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n450), .A2(KEYINPUT77), .A3(new_n448), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n456), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n453), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n406), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n464), .B1(new_n463), .B2(new_n296), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n434), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT6), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n477), .A2(new_n478), .A3(G107), .ZN(new_n479));
  XNOR2_X1  g0279(.A(G97), .B(G107), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  OAI22_X1  g0281(.A1(new_n481), .A2(new_n221), .B1(new_n393), .B2(new_n267), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n398), .B1(new_n322), .B2(new_n323), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n249), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n251), .A2(G97), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n485), .B1(new_n431), .B2(G97), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n283), .A2(new_n285), .A3(G244), .A4(new_n287), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n291), .A2(KEYINPUT4), .A3(G244), .A4(new_n287), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G283), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n291), .A2(G250), .A3(G1698), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n294), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n451), .A2(G257), .A3(new_n280), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n460), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n487), .B1(G200), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n406), .B2(new_n497), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n261), .A2(KEYINPUT19), .A3(new_n478), .ZN(new_n500));
  INV_X1    g0300(.A(G87), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(new_n478), .C1(new_n396), .C2(new_n397), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n221), .B1(new_n278), .B2(new_n478), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n500), .B1(new_n504), .B2(KEYINPUT19), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n283), .A2(new_n285), .A3(new_n221), .A4(G68), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT79), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n291), .A2(KEYINPUT79), .A3(new_n221), .A4(G68), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n249), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n379), .A2(new_n390), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n431), .A2(G87), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n445), .A2(G274), .ZN(new_n515));
  OAI21_X1  g0315(.A(G250), .B1(new_n444), .B2(G1), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n294), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n283), .A2(new_n285), .A3(G244), .A4(G1698), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n283), .A2(new_n285), .A3(G238), .A4(new_n287), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n519), .C1(new_n278), .C2(new_n415), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n517), .B1(new_n520), .B2(new_n294), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n521), .A2(new_n296), .ZN(new_n522));
  AOI211_X1 g0322(.A(new_n406), .B(new_n517), .C1(new_n520), .C2(new_n294), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n520), .A2(new_n294), .ZN(new_n525));
  INV_X1    g0325(.A(new_n517), .ZN(new_n526));
  AOI21_X1  g0326(.A(G169), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI211_X1 g0327(.A(G179), .B(new_n517), .C1(new_n520), .C2(new_n294), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n390), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT80), .B1(new_n431), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT80), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n430), .A2(new_n532), .A3(new_n390), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n511), .A2(new_n534), .A3(new_n512), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n514), .A2(new_n524), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n497), .A2(new_n336), .B1(new_n484), .B2(new_n486), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n495), .A2(new_n460), .A3(new_n304), .A4(new_n496), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n499), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n492), .B(new_n221), .C1(G33), .C2(new_n478), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n541), .B(new_n249), .C1(new_n221), .C2(G116), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT20), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n379), .A2(new_n415), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n376), .A2(G116), .A3(new_n250), .A4(new_n429), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n288), .A2(G264), .B1(G303), .B2(new_n286), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n308), .A2(G257), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n280), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT81), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n451), .A2(G270), .A3(new_n280), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n460), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n552), .B1(new_n460), .B2(new_n553), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n551), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n547), .B1(new_n557), .B2(G200), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n406), .B2(new_n557), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n476), .A2(new_n540), .A3(new_n559), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n463), .A2(new_n304), .B1(new_n336), .B2(new_n472), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n433), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n451), .A2(G270), .A3(new_n280), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT81), .B1(new_n563), .B2(new_n471), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n550), .B1(new_n564), .B2(new_n554), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n547), .A2(G169), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT82), .ZN(new_n569));
  INV_X1    g0369(.A(new_n567), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n557), .A2(KEYINPUT21), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT82), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT83), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n565), .A2(G179), .A3(new_n547), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n569), .A2(new_n573), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT21), .B1(new_n557), .B2(new_n570), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n569), .A2(new_n573), .A3(new_n575), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n577), .B1(new_n578), .B2(KEYINPUT83), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n560), .A2(new_n562), .A3(new_n576), .A4(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n414), .A2(new_n580), .ZN(G372));
  INV_X1    g0381(.A(new_n384), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n582), .A2(new_n412), .ZN(new_n583));
  XNOR2_X1  g0383(.A(new_n333), .B(KEYINPUT17), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n387), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT18), .B1(new_n346), .B2(new_n347), .ZN(new_n586));
  AOI211_X1 g0386(.A(new_n349), .B(new_n351), .C1(new_n345), .C2(new_n339), .ZN(new_n587));
  OAI22_X1  g0387(.A1(new_n583), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n299), .B(KEYINPUT10), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n305), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n529), .A2(new_n535), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n497), .A2(new_n336), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n592), .A2(new_n538), .A3(new_n487), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n536), .A3(KEYINPUT26), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT26), .B1(new_n593), .B2(new_n536), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n578), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT87), .ZN(new_n599));
  INV_X1    g0399(.A(new_n577), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT87), .B1(new_n578), .B2(new_n577), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(new_n562), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n476), .A2(new_n540), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n597), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n590), .B1(new_n414), .B2(new_n605), .ZN(G369));
  NAND2_X1  g0406(.A1(new_n579), .A2(new_n576), .ZN(new_n607));
  INV_X1    g0407(.A(new_n547), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n221), .A2(G13), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n245), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n610), .A2(KEYINPUT27), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(KEYINPUT27), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(G213), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(G343), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n607), .B1(new_n608), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n601), .A2(new_n602), .A3(new_n547), .A4(new_n615), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n559), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(G330), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n433), .A2(new_n615), .ZN(new_n622));
  XOR2_X1   g0422(.A(new_n622), .B(KEYINPUT88), .Z(new_n623));
  AND3_X1   g0423(.A1(new_n623), .A2(new_n562), .A3(new_n476), .ZN(new_n624));
  INV_X1    g0424(.A(new_n562), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n624), .B1(new_n625), .B2(new_n615), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n615), .B1(new_n579), .B2(new_n576), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n624), .A2(new_n629), .B1(new_n625), .B2(new_n616), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(G399));
  INV_X1    g0431(.A(new_n502), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n415), .ZN(new_n633));
  INV_X1    g0433(.A(new_n215), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(G41), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n633), .A2(new_n245), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n219), .B2(new_n635), .ZN(new_n637));
  XOR2_X1   g0437(.A(new_n637), .B(KEYINPUT28), .Z(new_n638));
  NOR3_X1   g0438(.A1(new_n605), .A2(KEYINPUT29), .A3(new_n615), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n575), .B1(new_n568), .B2(KEYINPUT82), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n571), .A2(new_n572), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT83), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n642), .A2(new_n562), .A3(new_n576), .A4(new_n600), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n604), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT91), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT91), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n643), .A2(new_n646), .A3(new_n604), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n594), .B1(new_n596), .B2(KEYINPUT89), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n593), .A2(new_n536), .A3(new_n649), .A4(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT90), .B1(new_n651), .B2(new_n591), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT90), .ZN(new_n653));
  INV_X1    g0453(.A(new_n591), .ZN(new_n654));
  AOI211_X1 g0454(.A(new_n653), .B(new_n654), .C1(new_n648), .C2(new_n650), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n645), .A2(new_n647), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n616), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n639), .B1(new_n658), .B2(KEYINPUT29), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT31), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n565), .A2(G179), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n454), .A2(new_n462), .ZN(new_n663));
  INV_X1    g0463(.A(new_n521), .ZN(new_n664));
  NOR4_X1   g0464(.A1(new_n662), .A2(new_n663), .A3(new_n664), .A4(new_n497), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT30), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT30), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n521), .A2(G179), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n463), .A2(new_n557), .A3(new_n497), .A4(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n661), .B1(new_n670), .B2(new_n615), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n580), .B2(new_n615), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(new_n661), .A3(new_n615), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n620), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n660), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n638), .B1(new_n676), .B2(G1), .ZN(G364));
  NOR2_X1   g0477(.A1(new_n634), .A2(new_n291), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n243), .A2(new_n444), .ZN(new_n680));
  AOI211_X1 g0480(.A(new_n679), .B(new_n680), .C1(new_n444), .C2(new_n219), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT92), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n634), .A2(new_n286), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G355), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(G116), .B2(new_n215), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n681), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n682), .B2(new_n685), .ZN(new_n687));
  NOR2_X1   g0487(.A1(G13), .A2(G33), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OR3_X1    g0489(.A1(new_n689), .A2(KEYINPUT93), .A3(G20), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT93), .B1(new_n689), .B2(G20), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n220), .B1(G20), .B2(new_n336), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n245), .B1(new_n609), .B2(G45), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n635), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n221), .A2(new_n406), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n304), .A2(G200), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n221), .A2(G190), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n700), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI22_X1  g0505(.A1(G58), .A2(new_n702), .B1(new_n705), .B2(G77), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(KEYINPUT94), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(KEYINPUT94), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n304), .A2(new_n296), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n699), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n296), .A2(G179), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n699), .A2(new_n711), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n710), .A2(new_n238), .B1(new_n712), .B2(new_n501), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n709), .A2(new_n703), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n713), .B1(G68), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n707), .A2(new_n708), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n703), .A2(new_n711), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n286), .B1(new_n719), .B2(G107), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G179), .A2(G200), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n703), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G159), .ZN(new_n723));
  OR3_X1    g0523(.A1(new_n722), .A2(KEYINPUT32), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT32), .B1(new_n722), .B2(new_n723), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n221), .B1(new_n721), .B2(G190), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n478), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n720), .A2(new_n724), .A3(new_n725), .A4(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n722), .ZN(new_n730));
  AOI22_X1  g0530(.A1(G322), .A2(new_n702), .B1(new_n730), .B2(G329), .ZN(new_n731));
  INV_X1    g0531(.A(new_n712), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G303), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G326), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n710), .A2(new_n735), .B1(new_n726), .B2(new_n436), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT95), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n291), .B1(new_n719), .B2(G283), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT33), .B(G317), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n715), .A2(new_n740), .B1(new_n705), .B2(G311), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n734), .A2(new_n738), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n736), .A2(new_n737), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n717), .A2(new_n729), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n693), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n695), .A2(new_n698), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n619), .B2(new_n692), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n621), .A2(new_n698), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n619), .A2(new_n620), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(G396));
  AND2_X1   g0551(.A1(new_n395), .A2(new_n615), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n408), .A2(new_n752), .B1(new_n411), .B2(new_n410), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n412), .A2(new_n616), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(new_n605), .B2(new_n615), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n675), .B(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n605), .A2(new_n615), .A3(new_n755), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(KEYINPUT97), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n698), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(new_n759), .B2(new_n757), .ZN(new_n761));
  INV_X1    g0561(.A(new_n698), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n693), .A2(new_n688), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n762), .B1(new_n393), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n693), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n718), .A2(new_n501), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n291), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n767), .B1(new_n768), .B2(new_n714), .C1(new_n436), .C2(new_n701), .ZN(new_n769));
  INV_X1    g0569(.A(G303), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n710), .A2(new_n770), .B1(new_n722), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G107), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n712), .A2(new_n773), .B1(new_n704), .B2(new_n415), .ZN(new_n774));
  NOR4_X1   g0574(.A1(new_n769), .A2(new_n727), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n710), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G137), .A2(new_n776), .B1(new_n705), .B2(G159), .ZN(new_n777));
  INV_X1    g0577(.A(G143), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n777), .B1(new_n778), .B2(new_n701), .C1(new_n265), .C2(new_n714), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT34), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n719), .A2(G68), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n238), .B2(new_n712), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n782), .A2(KEYINPUT96), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(KEYINPUT96), .ZN(new_n784));
  INV_X1    g0584(.A(G132), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n291), .B1(new_n726), .B2(new_n201), .C1(new_n785), .C2(new_n722), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n775), .B1(new_n780), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n755), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n764), .B1(new_n765), .B2(new_n788), .C1(new_n789), .C2(new_n689), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n761), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G384));
  INV_X1    g0592(.A(new_n481), .ZN(new_n793));
  OAI211_X1 g0593(.A(G116), .B(new_n222), .C1(new_n793), .C2(KEYINPUT35), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(KEYINPUT35), .B2(new_n793), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT36), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n219), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n245), .B(G13), .C1(new_n797), .C2(new_n239), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT98), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n383), .A2(new_n615), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI221_X4 g0602(.A(new_n802), .B1(new_n386), .B2(new_n385), .C1(new_n367), .C2(new_n383), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n384), .A2(new_n616), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n384), .A2(new_n387), .A3(new_n801), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n806), .B(KEYINPUT98), .C1(new_n384), .C2(new_n616), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n808), .A2(new_n672), .A3(new_n673), .A4(new_n789), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT38), .ZN(new_n811));
  INV_X1    g0611(.A(new_n613), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n347), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n333), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n348), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT37), .B1(new_n352), .B2(new_n814), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n584), .B1(new_n587), .B2(new_n586), .ZN(new_n819));
  INV_X1    g0619(.A(new_n813), .ZN(new_n820));
  AOI221_X4 g0620(.A(new_n811), .B1(new_n817), .B2(new_n818), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n817), .A2(new_n818), .ZN(new_n823));
  AOI21_X1  g0623(.A(KEYINPUT38), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT40), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(KEYINPUT100), .A2(KEYINPUT40), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n810), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n822), .A2(KEYINPUT38), .A3(new_n823), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n817), .A2(new_n818), .A3(KEYINPUT99), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT99), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n832), .B(KEYINPUT37), .C1(new_n352), .C2(new_n814), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n831), .B(new_n833), .C1(new_n354), .C2(new_n813), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n811), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n809), .A2(KEYINPUT100), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n829), .B1(new_n836), .B2(new_n826), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n674), .A2(new_n414), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(G330), .A3(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n754), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n808), .B1(new_n758), .B2(new_n842), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n843), .A2(new_n825), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n350), .A2(new_n353), .A3(new_n613), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT39), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n835), .A2(new_n846), .A3(new_n830), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT39), .B1(new_n821), .B2(new_n824), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n384), .A2(new_n615), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n844), .A2(new_n845), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n841), .B(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n590), .ZN(new_n855));
  INV_X1    g0655(.A(new_n414), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n660), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n245), .B2(new_n609), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n854), .A2(new_n857), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n799), .B1(new_n859), .B2(new_n860), .ZN(G367));
  OAI221_X1 g0661(.A(new_n694), .B1(new_n215), .B2(new_n390), .C1(new_n233), .C2(new_n679), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT104), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n762), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n863), .B2(new_n862), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n478), .A2(new_n718), .B1(new_n704), .B2(new_n768), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n291), .B(new_n866), .C1(G303), .C2(new_n702), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n732), .A2(KEYINPUT46), .A3(G116), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT46), .B1(new_n732), .B2(G116), .ZN(new_n869));
  INV_X1    g0669(.A(new_n726), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n869), .B1(new_n399), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(G317), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n710), .A2(new_n771), .B1(new_n722), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(G294), .B2(new_n715), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n867), .A2(new_n868), .A3(new_n871), .A4(new_n874), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n714), .A2(new_n723), .B1(new_n704), .B2(new_n238), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT105), .ZN(new_n877));
  AOI22_X1  g0677(.A1(G58), .A2(new_n732), .B1(new_n702), .B2(G150), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n718), .A2(new_n393), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(G143), .B2(new_n776), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n726), .A2(new_n202), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n286), .B(new_n881), .C1(G137), .C2(new_n730), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n877), .A2(new_n878), .A3(new_n880), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT47), .B1(new_n875), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(new_n765), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n875), .A2(KEYINPUT47), .A3(new_n883), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n865), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n514), .A2(new_n616), .ZN(new_n888));
  MUX2_X1   g0688(.A(new_n536), .B(new_n654), .S(new_n888), .Z(new_n889));
  INV_X1    g0689(.A(new_n692), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n487), .A2(new_n615), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n499), .A2(new_n539), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n593), .A2(new_n615), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n630), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g0696(.A1(KEYINPUT102), .A2(KEYINPUT44), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(KEYINPUT102), .B2(KEYINPUT44), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n897), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n630), .A2(new_n895), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n902), .B(KEYINPUT45), .Z(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n628), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT103), .ZN(new_n907));
  INV_X1    g0707(.A(new_n621), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n624), .A2(new_n629), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n627), .B2(new_n629), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n905), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n676), .A2(new_n911), .ZN(new_n912));
  OR3_X1    g0712(.A1(new_n906), .A2(new_n907), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n676), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n635), .B(KEYINPUT41), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n697), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n624), .A2(new_n629), .A3(new_n895), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n539), .B1(new_n562), .B2(new_n893), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n917), .A2(KEYINPUT42), .B1(new_n616), .B2(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n918), .A2(new_n920), .B1(KEYINPUT43), .B2(new_n889), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n921), .B(new_n922), .Z(new_n923));
  NAND2_X1  g0723(.A1(new_n905), .A2(new_n895), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n926), .A2(KEYINPUT101), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(KEYINPUT101), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n891), .B1(new_n916), .B2(new_n930), .ZN(G387));
  NAND2_X1  g0731(.A1(new_n911), .A2(new_n697), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT106), .ZN(new_n933));
  XNOR2_X1  g0733(.A(KEYINPUT107), .B(G150), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n712), .A2(new_n393), .B1(new_n722), .B2(new_n934), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n286), .B(new_n935), .C1(G97), .C2(new_n719), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n726), .A2(new_n390), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n260), .A2(new_n715), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n701), .A2(new_n238), .B1(new_n704), .B2(new_n202), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G159), .B2(new_n776), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n936), .A2(new_n938), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n291), .B1(new_n730), .B2(G326), .ZN(new_n943));
  AOI22_X1  g0743(.A1(G322), .A2(new_n776), .B1(new_n705), .B2(G303), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n944), .B1(new_n771), .B2(new_n714), .C1(new_n872), .C2(new_n701), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT48), .Z(new_n946));
  OAI22_X1  g0746(.A1(new_n712), .A2(new_n436), .B1(new_n726), .B2(new_n768), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n943), .B1(new_n415), .B2(new_n718), .C1(new_n948), .C2(KEYINPUT49), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n948), .A2(KEYINPUT49), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n942), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n693), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n230), .A2(new_n444), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n953), .A2(new_n678), .B1(new_n633), .B2(new_n683), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n391), .A2(G50), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT50), .Z(new_n956));
  OAI21_X1  g0756(.A(new_n444), .B1(new_n202), .B2(new_n393), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n956), .A2(new_n633), .A3(new_n957), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n954), .A2(new_n958), .B1(G107), .B2(new_n215), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n762), .B1(new_n959), .B2(new_n694), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n952), .B(new_n960), .C1(new_n627), .C2(new_n890), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n676), .A2(new_n911), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n912), .A2(new_n635), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n933), .B(new_n961), .C1(new_n962), .C2(new_n963), .ZN(G393));
  AOI21_X1  g0764(.A(new_n628), .B1(new_n901), .B2(new_n903), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n912), .B1(new_n906), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n913), .A2(new_n635), .A3(new_n966), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n906), .A2(new_n696), .A3(new_n965), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n893), .A2(new_n692), .A3(new_n894), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n694), .B1(new_n478), .B2(new_n215), .C1(new_n237), .C2(new_n679), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n762), .B1(new_n970), .B2(KEYINPUT108), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(KEYINPUT108), .B2(new_n970), .ZN(new_n972));
  AOI22_X1  g0772(.A1(G283), .A2(new_n732), .B1(new_n730), .B2(G322), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n973), .B(new_n286), .C1(new_n773), .C2(new_n718), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT111), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n710), .A2(new_n872), .B1(new_n701), .B2(new_n771), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT52), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n714), .A2(new_n770), .B1(new_n704), .B2(new_n436), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G116), .B2(new_n870), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n975), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n710), .A2(new_n265), .B1(new_n701), .B2(new_n723), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT109), .Z(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(KEYINPUT51), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(KEYINPUT51), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n714), .A2(new_n238), .B1(new_n704), .B2(new_n391), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n726), .A2(new_n393), .ZN(new_n986));
  NOR4_X1   g0786(.A1(new_n985), .A2(new_n766), .A3(new_n986), .A4(new_n286), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n712), .A2(new_n202), .B1(new_n722), .B2(new_n778), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT110), .Z(new_n989));
  NAND3_X1  g0789(.A1(new_n984), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n980), .B1(new_n983), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n972), .B1(new_n991), .B2(new_n693), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n968), .B1(new_n969), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n967), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(KEYINPUT112), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT112), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n967), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(G390));
  INV_X1    g0798(.A(new_n850), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n849), .B1(new_n843), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n657), .A2(new_n616), .A3(new_n753), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n754), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n808), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT113), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n850), .B1(new_n835), .B2(new_n830), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n808), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n1001), .B2(new_n754), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1005), .ZN(new_n1009));
  OAI21_X1  g0809(.A(KEYINPUT113), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1000), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n809), .A2(new_n620), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1012), .B(new_n1000), .C1(new_n1006), .C2(new_n1010), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n675), .A2(new_n856), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1017), .B(new_n590), .C1(new_n659), .C2(new_n414), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n672), .A2(G330), .A3(new_n673), .A4(new_n789), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n810), .A2(G330), .B1(new_n1019), .B2(new_n1007), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n758), .A2(new_n842), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1020), .A2(new_n754), .A3(new_n1001), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1018), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OR3_X1    g0824(.A1(new_n1016), .A2(KEYINPUT114), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(KEYINPUT114), .B1(new_n1016), .B2(new_n1024), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n635), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n1016), .B2(new_n1024), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1000), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1004), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1008), .A2(new_n1009), .A3(KEYINPUT113), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n1012), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1034), .A2(new_n697), .A3(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT115), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(KEYINPUT115), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n847), .A2(new_n848), .A3(new_n688), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n763), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n698), .B1(new_n260), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n712), .A2(new_n934), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT53), .ZN(new_n1043));
  XOR2_X1   g0843(.A(KEYINPUT54), .B(G143), .Z(new_n1044));
  AOI22_X1  g0844(.A1(new_n705), .A2(new_n1044), .B1(new_n719), .B2(G50), .ZN(new_n1045));
  INV_X1    g0845(.A(G128), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1043), .B(new_n1045), .C1(new_n1046), .C2(new_n710), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G132), .A2(new_n702), .B1(new_n715), .B2(G137), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n286), .B1(new_n730), .B2(G125), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n723), .C2(new_n726), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G283), .A2(new_n776), .B1(new_n705), .B2(G97), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n415), .B2(new_n701), .C1(new_n398), .C2(new_n714), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n291), .B1(new_n732), .B2(G87), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n730), .A2(G294), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n986), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n781), .A4(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1047), .A2(new_n1050), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1041), .B1(new_n1057), .B2(new_n693), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1037), .A2(new_n1038), .B1(new_n1039), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1029), .A2(new_n1059), .ZN(G378));
  NAND3_X1  g0860(.A1(new_n1034), .A2(new_n1024), .A3(new_n1035), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1018), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT119), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT119), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1061), .A2(new_n1065), .A3(new_n1062), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT55), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n301), .B2(new_n305), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n305), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n589), .A2(KEYINPUT55), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n270), .A2(new_n613), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1069), .B(new_n1071), .C1(new_n270), .C2(new_n613), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1075), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n837), .A2(G330), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n837), .B2(G330), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n852), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n837), .A2(G330), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1079), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n837), .A2(G330), .A3(new_n1079), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n853), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1082), .A2(new_n1087), .A3(KEYINPUT118), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT118), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1089), .B(new_n852), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT57), .B1(new_n1067), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT57), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1061), .A2(new_n1065), .A3(new_n1062), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1065), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n635), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1092), .A2(new_n1098), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1046), .A2(new_n701), .B1(new_n714), .B2(new_n785), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n732), .A2(new_n1044), .B1(new_n705), .B2(G137), .ZN(new_n1101));
  INV_X1    g0901(.A(G125), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n710), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1100), .B(new_n1103), .C1(G150), .C2(new_n870), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT59), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n719), .A2(G159), .ZN(new_n1108));
  AOI211_X1 g0908(.A(G33), .B(G41), .C1(new_n730), .C2(G124), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT116), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n702), .B2(G107), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n701), .A2(KEYINPUT116), .A3(new_n773), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1112), .A2(new_n881), .A3(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n390), .A2(new_n704), .B1(new_n718), .B2(new_n201), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G116), .B2(new_n776), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G77), .A2(new_n732), .B1(new_n730), .B2(G283), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n286), .A2(new_n279), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G97), .B2(new_n715), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT58), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1118), .B(new_n238), .C1(G33), .C2(G41), .ZN(new_n1124));
  AND4_X1   g0924(.A1(new_n1110), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n698), .B1(G50), .B2(new_n1040), .C1(new_n1125), .C2(new_n765), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n1084), .B2(new_n688), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n1091), .B2(new_n697), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1099), .A2(new_n1128), .ZN(G375));
  OAI21_X1  g0929(.A(new_n291), .B1(new_n718), .B2(new_n201), .ZN(new_n1130));
  INV_X1    g0930(.A(G137), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n710), .A2(new_n785), .B1(new_n701), .B2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1130), .B(new_n1132), .C1(G50), .C2(new_n870), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n712), .A2(new_n723), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n704), .A2(new_n265), .B1(new_n722), .B2(new_n1046), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(new_n715), .C2(new_n1044), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n398), .A2(new_n704), .B1(new_n710), .B2(new_n436), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n714), .A2(new_n415), .B1(new_n722), .B2(new_n770), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n478), .A2(new_n712), .B1(new_n701), .B2(new_n768), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1140), .A2(new_n879), .A3(new_n937), .A4(new_n291), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1133), .A2(new_n1136), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n698), .B1(G68), .B2(new_n1040), .C1(new_n1142), .C2(new_n765), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1007), .B2(new_n688), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n697), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1024), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n915), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1145), .A2(new_n1062), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(G381));
  INV_X1    g0950(.A(G375), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1029), .A2(new_n1059), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(G390), .A2(G387), .ZN(new_n1153));
  NOR4_X1   g0953(.A1(G381), .A2(G393), .A3(G384), .A4(G396), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(G407));
  NAND2_X1  g0955(.A1(new_n614), .A2(G213), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT120), .Z(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1151), .A2(new_n1152), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(G407), .A2(new_n1159), .A3(G213), .ZN(G409));
  OAI21_X1  g0960(.A(new_n1147), .B1(new_n1149), .B2(KEYINPUT60), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT122), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1027), .B1(new_n1149), .B2(KEYINPUT60), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n1146), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n791), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(G384), .A3(new_n1146), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(G2897), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n1156), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1170), .A2(G2897), .A3(new_n1158), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT124), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(G378), .B(new_n1128), .C1(new_n1092), .C2(new_n1098), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1091), .B(new_n915), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1127), .B1(new_n1180), .B2(new_n697), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n1152), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(KEYINPUT121), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT121), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1178), .A2(new_n1183), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1156), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1173), .A2(KEYINPUT124), .A3(new_n1174), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1177), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(G393), .B(new_n750), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(G390), .A2(G387), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n1153), .ZN(new_n1194));
  OR2_X1    g0994(.A1(G390), .A2(G387), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(G390), .A2(G387), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(new_n1191), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1158), .B1(new_n1178), .B2(new_n1183), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(KEYINPUT63), .A3(new_n1171), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT61), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1185), .A2(new_n1156), .A3(new_n1171), .A4(new_n1187), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1205));
  OAI211_X1 g1005(.A(new_n1190), .B(new_n1202), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1201), .B1(new_n1175), .B2(new_n1199), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1199), .A2(KEYINPUT62), .A3(new_n1171), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT62), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1203), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT125), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1208), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1203), .A2(KEYINPUT125), .A3(new_n1209), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1207), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1206), .B1(new_n1214), .B2(new_n1198), .ZN(G405));
  NAND2_X1  g1015(.A1(new_n1170), .A2(KEYINPUT126), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1198), .B(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1151), .A2(G378), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n1178), .C1(KEYINPUT126), .C2(new_n1170), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1217), .B(new_n1220), .Z(G402));
endmodule


