

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  NAND2_X1 U324 ( .A1(n563), .A2(n569), .ZN(n292) );
  INV_X1 U325 ( .A(KEYINPUT70), .ZN(n304) );
  XNOR2_X1 U326 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U327 ( .A(n307), .B(n306), .ZN(n308) );
  AND2_X1 U328 ( .A1(n558), .A2(n451), .ZN(n575) );
  INV_X1 U329 ( .A(G204GAT), .ZN(n453) );
  XOR2_X1 U330 ( .A(n556), .B(KEYINPUT28), .Z(n521) );
  XNOR2_X1 U331 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U332 ( .A(n456), .B(n455), .ZN(G1353GAT) );
  XOR2_X1 U333 ( .A(G64GAT), .B(G92GAT), .Z(n294) );
  XNOR2_X1 U334 ( .A(G176GAT), .B(G204GAT), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n294), .B(n293), .ZN(n383) );
  XOR2_X1 U336 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n296) );
  XNOR2_X1 U337 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U339 ( .A(G120GAT), .B(G71GAT), .Z(n415) );
  XOR2_X1 U340 ( .A(G99GAT), .B(G85GAT), .Z(n328) );
  XNOR2_X1 U341 ( .A(n415), .B(n328), .ZN(n298) );
  XOR2_X1 U342 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U344 ( .A(n300), .B(n299), .Z(n302) );
  NAND2_X1 U345 ( .A1(G230GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n302), .B(n301), .ZN(n307) );
  XNOR2_X1 U347 ( .A(G106GAT), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n303), .B(G148GAT), .ZN(n410) );
  XNOR2_X1 U349 ( .A(n410), .B(KEYINPUT71), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n383), .B(n308), .ZN(n310) );
  XNOR2_X1 U351 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n309) );
  XOR2_X1 U352 ( .A(n309), .B(KEYINPUT69), .Z(n345) );
  XNOR2_X1 U353 ( .A(n310), .B(n345), .ZN(n470) );
  XOR2_X1 U354 ( .A(G92GAT), .B(G106GAT), .Z(n312) );
  XNOR2_X1 U355 ( .A(G134GAT), .B(G218GAT), .ZN(n311) );
  XNOR2_X1 U356 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U357 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n314) );
  XNOR2_X1 U358 ( .A(KEYINPUT79), .B(KEYINPUT10), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U360 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U361 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n318) );
  NAND2_X1 U362 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U363 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U364 ( .A(KEYINPUT9), .B(n319), .ZN(n320) );
  XNOR2_X1 U365 ( .A(n321), .B(n320), .ZN(n326) );
  XOR2_X1 U366 ( .A(KEYINPUT7), .B(KEYINPUT67), .Z(n323) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G29GAT), .ZN(n322) );
  XNOR2_X1 U368 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U369 ( .A(KEYINPUT8), .B(n324), .Z(n354) );
  INV_X1 U370 ( .A(n354), .ZN(n325) );
  XNOR2_X1 U371 ( .A(n326), .B(n325), .ZN(n331) );
  XNOR2_X1 U372 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n327) );
  XNOR2_X1 U373 ( .A(n327), .B(G162GAT), .ZN(n404) );
  XNOR2_X1 U374 ( .A(n404), .B(n328), .ZN(n329) );
  XOR2_X1 U375 ( .A(G36GAT), .B(G190GAT), .Z(n382) );
  XOR2_X1 U376 ( .A(n329), .B(n382), .Z(n330) );
  XOR2_X1 U377 ( .A(n331), .B(n330), .Z(n570) );
  XOR2_X1 U378 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n333) );
  XNOR2_X1 U379 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n332) );
  XNOR2_X1 U380 ( .A(n333), .B(n332), .ZN(n340) );
  XOR2_X1 U381 ( .A(G155GAT), .B(G78GAT), .Z(n335) );
  XNOR2_X1 U382 ( .A(G127GAT), .B(G71GAT), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U384 ( .A(G8GAT), .B(G183GAT), .Z(n386) );
  XOR2_X1 U385 ( .A(n336), .B(n386), .Z(n338) );
  XNOR2_X1 U386 ( .A(G22GAT), .B(G211GAT), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U388 ( .A(n340), .B(n339), .ZN(n349) );
  XOR2_X1 U389 ( .A(KEYINPUT82), .B(KEYINPUT15), .Z(n342) );
  NAND2_X1 U390 ( .A1(G231GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U391 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U392 ( .A(n343), .B(KEYINPUT14), .Z(n347) );
  XNOR2_X1 U393 ( .A(G15GAT), .B(G1GAT), .ZN(n344) );
  XNOR2_X1 U394 ( .A(n344), .B(KEYINPUT68), .ZN(n361) );
  XOR2_X1 U395 ( .A(n361), .B(n345), .Z(n346) );
  XNOR2_X1 U396 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U397 ( .A(n349), .B(n348), .ZN(n483) );
  INV_X1 U398 ( .A(KEYINPUT41), .ZN(n350) );
  XNOR2_X1 U399 ( .A(n350), .B(n470), .ZN(n500) );
  INV_X1 U400 ( .A(n500), .ZN(n563) );
  XOR2_X1 U401 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n352) );
  XNOR2_X1 U402 ( .A(G113GAT), .B(G8GAT), .ZN(n351) );
  XNOR2_X1 U403 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n365) );
  XOR2_X1 U405 ( .A(G141GAT), .B(G22GAT), .Z(n400) );
  XOR2_X1 U406 ( .A(G197GAT), .B(G50GAT), .Z(n356) );
  XNOR2_X1 U407 ( .A(G169GAT), .B(G36GAT), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U409 ( .A(n400), .B(n357), .Z(n359) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U412 ( .A(n360), .B(KEYINPUT65), .Z(n363) );
  XNOR2_X1 U413 ( .A(n361), .B(KEYINPUT66), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U415 ( .A(n365), .B(n364), .ZN(n576) );
  NAND2_X1 U416 ( .A1(n563), .A2(n576), .ZN(n368) );
  XOR2_X1 U417 ( .A(KEYINPUT108), .B(KEYINPUT46), .Z(n366) );
  XNOR2_X1 U418 ( .A(KEYINPUT107), .B(n366), .ZN(n367) );
  XNOR2_X1 U419 ( .A(n368), .B(n367), .ZN(n369) );
  AND2_X1 U420 ( .A1(n483), .A2(n369), .ZN(n370) );
  XNOR2_X1 U421 ( .A(n370), .B(KEYINPUT109), .ZN(n371) );
  NOR2_X1 U422 ( .A1(n570), .A2(n371), .ZN(n372) );
  XNOR2_X1 U423 ( .A(n372), .B(KEYINPUT47), .ZN(n379) );
  XOR2_X1 U424 ( .A(n570), .B(KEYINPUT98), .Z(n373) );
  XNOR2_X1 U425 ( .A(n373), .B(KEYINPUT36), .ZN(n583) );
  NOR2_X1 U426 ( .A1(n483), .A2(n583), .ZN(n374) );
  XNOR2_X1 U427 ( .A(n374), .B(KEYINPUT45), .ZN(n375) );
  NAND2_X1 U428 ( .A1(n375), .A2(n470), .ZN(n376) );
  NOR2_X1 U429 ( .A1(n576), .A2(n376), .ZN(n377) );
  XOR2_X1 U430 ( .A(KEYINPUT110), .B(n377), .Z(n378) );
  NAND2_X1 U431 ( .A1(n379), .A2(n378), .ZN(n381) );
  XNOR2_X1 U432 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n380) );
  XNOR2_X1 U433 ( .A(n381), .B(n380), .ZN(n524) );
  XOR2_X1 U434 ( .A(n383), .B(n382), .Z(n385) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U436 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U437 ( .A(n387), .B(n386), .Z(n394) );
  XOR2_X1 U438 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n389) );
  XNOR2_X1 U439 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n388) );
  XNOR2_X1 U440 ( .A(n389), .B(n388), .ZN(n414) );
  XOR2_X1 U441 ( .A(KEYINPUT21), .B(G218GAT), .Z(n391) );
  XNOR2_X1 U442 ( .A(KEYINPUT88), .B(G211GAT), .ZN(n390) );
  XNOR2_X1 U443 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U444 ( .A(G197GAT), .B(n392), .Z(n411) );
  XNOR2_X1 U445 ( .A(n414), .B(n411), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n394), .B(n393), .ZN(n475) );
  XOR2_X1 U447 ( .A(KEYINPUT122), .B(n475), .Z(n395) );
  NOR2_X1 U448 ( .A1(n524), .A2(n395), .ZN(n396) );
  XNOR2_X1 U449 ( .A(n396), .B(KEYINPUT54), .ZN(n558) );
  XOR2_X1 U450 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n398) );
  XNOR2_X1 U451 ( .A(KEYINPUT22), .B(G204GAT), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U453 ( .A(n400), .B(n399), .Z(n402) );
  NAND2_X1 U454 ( .A1(G228GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U455 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U456 ( .A(n403), .B(KEYINPUT23), .Z(n406) );
  XNOR2_X1 U457 ( .A(n404), .B(KEYINPUT87), .ZN(n405) );
  XNOR2_X1 U458 ( .A(n406), .B(n405), .ZN(n409) );
  XOR2_X1 U459 ( .A(G155GAT), .B(KEYINPUT3), .Z(n408) );
  XNOR2_X1 U460 ( .A(KEYINPUT2), .B(KEYINPUT89), .ZN(n407) );
  XNOR2_X1 U461 ( .A(n408), .B(n407), .ZN(n441) );
  XOR2_X1 U462 ( .A(n409), .B(n441), .Z(n413) );
  XNOR2_X1 U463 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U464 ( .A(n413), .B(n412), .ZN(n556) );
  XOR2_X1 U465 ( .A(n415), .B(n414), .Z(n417) );
  XNOR2_X1 U466 ( .A(G99GAT), .B(G190GAT), .ZN(n416) );
  XNOR2_X1 U467 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U468 ( .A(KEYINPUT86), .B(G176GAT), .Z(n419) );
  NAND2_X1 U469 ( .A1(G227GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U470 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U471 ( .A(n421), .B(n420), .Z(n426) );
  XOR2_X1 U472 ( .A(KEYINPUT85), .B(G183GAT), .Z(n423) );
  XNOR2_X1 U473 ( .A(G43GAT), .B(G15GAT), .ZN(n422) );
  XNOR2_X1 U474 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U475 ( .A(n424), .B(KEYINPUT20), .ZN(n425) );
  XNOR2_X1 U476 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U477 ( .A(KEYINPUT0), .B(G134GAT), .Z(n428) );
  XNOR2_X1 U478 ( .A(KEYINPUT84), .B(G127GAT), .ZN(n427) );
  XNOR2_X1 U479 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U480 ( .A(G113GAT), .B(n429), .Z(n450) );
  XNOR2_X1 U481 ( .A(n430), .B(n450), .ZN(n569) );
  INV_X1 U482 ( .A(n569), .ZN(n560) );
  NAND2_X1 U483 ( .A1(n556), .A2(n560), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n431), .B(KEYINPUT26), .ZN(n538) );
  XOR2_X1 U485 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n433) );
  NAND2_X1 U486 ( .A1(G225GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U488 ( .A(KEYINPUT92), .B(n434), .ZN(n448) );
  XOR2_X1 U489 ( .A(KEYINPUT1), .B(KEYINPUT91), .Z(n436) );
  XNOR2_X1 U490 ( .A(G141GAT), .B(G120GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U492 ( .A(KEYINPUT93), .B(G57GAT), .Z(n438) );
  XNOR2_X1 U493 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U495 ( .A(n440), .B(n439), .Z(n446) );
  XOR2_X1 U496 ( .A(G85GAT), .B(G162GAT), .Z(n443) );
  XNOR2_X1 U497 ( .A(G29GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U499 ( .A(G148GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n511) );
  INV_X1 U503 ( .A(n511), .ZN(n555) );
  NOR2_X1 U504 ( .A1(n538), .A2(n555), .ZN(n451) );
  INV_X1 U505 ( .A(KEYINPUT124), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n575), .B(n452), .ZN(n584) );
  OR2_X1 U507 ( .A1(n470), .A2(n584), .ZN(n456) );
  XOR2_X1 U508 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n454) );
  INV_X1 U509 ( .A(n475), .ZN(n515) );
  NOR2_X1 U510 ( .A1(n560), .A2(n515), .ZN(n457) );
  NOR2_X1 U511 ( .A1(n556), .A2(n457), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n458), .B(KEYINPUT95), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT25), .ZN(n462) );
  XOR2_X1 U514 ( .A(n475), .B(KEYINPUT94), .Z(n460) );
  XNOR2_X1 U515 ( .A(KEYINPUT27), .B(n460), .ZN(n464) );
  NOR2_X1 U516 ( .A1(n538), .A2(n464), .ZN(n461) );
  NOR2_X1 U517 ( .A1(n462), .A2(n461), .ZN(n463) );
  NOR2_X1 U518 ( .A1(n555), .A2(n463), .ZN(n466) );
  NOR2_X1 U519 ( .A1(n511), .A2(n464), .ZN(n540) );
  NAND2_X1 U520 ( .A1(n540), .A2(n521), .ZN(n526) );
  NOR2_X1 U521 ( .A1(n526), .A2(n569), .ZN(n465) );
  NOR2_X1 U522 ( .A1(n466), .A2(n465), .ZN(n484) );
  XOR2_X1 U523 ( .A(KEYINPUT16), .B(KEYINPUT83), .Z(n468) );
  OR2_X1 U524 ( .A1(n570), .A2(n483), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n468), .B(n467), .ZN(n469) );
  NOR2_X1 U526 ( .A1(n484), .A2(n469), .ZN(n501) );
  NAND2_X1 U527 ( .A1(n470), .A2(n576), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n471), .B(KEYINPUT75), .ZN(n488) );
  NAND2_X1 U529 ( .A1(n501), .A2(n488), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT96), .B(n472), .Z(n481) );
  NAND2_X1 U531 ( .A1(n481), .A2(n555), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(KEYINPUT34), .ZN(n474) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n474), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n481), .A2(n475), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U537 ( .A1(n481), .A2(n569), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U539 ( .A(G15GAT), .B(n479), .Z(G1326GAT) );
  INV_X1 U540 ( .A(n521), .ZN(n480) );
  NAND2_X1 U541 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n482), .B(G22GAT), .ZN(G1327GAT) );
  INV_X1 U543 ( .A(n483), .ZN(n580) );
  NOR2_X1 U544 ( .A1(n484), .A2(n580), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n485), .B(KEYINPUT99), .ZN(n486) );
  NOR2_X1 U546 ( .A1(n583), .A2(n486), .ZN(n487) );
  XOR2_X1 U547 ( .A(KEYINPUT37), .B(n487), .Z(n510) );
  NAND2_X1 U548 ( .A1(n510), .A2(n488), .ZN(n489) );
  XNOR2_X1 U549 ( .A(KEYINPUT38), .B(n489), .ZN(n497) );
  NOR2_X1 U550 ( .A1(n497), .A2(n511), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n497), .A2(n515), .ZN(n492) );
  XOR2_X1 U554 ( .A(KEYINPUT100), .B(n492), .Z(n493) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(n493), .ZN(G1329GAT) );
  XNOR2_X1 U556 ( .A(KEYINPUT40), .B(KEYINPUT101), .ZN(n495) );
  NOR2_X1 U557 ( .A1(n560), .A2(n497), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  NOR2_X1 U560 ( .A1(n521), .A2(n497), .ZN(n498) );
  XOR2_X1 U561 ( .A(KEYINPUT102), .B(n498), .Z(n499) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  NOR2_X1 U563 ( .A1(n576), .A2(n500), .ZN(n509) );
  NAND2_X1 U564 ( .A1(n509), .A2(n501), .ZN(n506) );
  NOR2_X1 U565 ( .A1(n511), .A2(n506), .ZN(n502) );
  XOR2_X1 U566 ( .A(G57GAT), .B(n502), .Z(n503) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U568 ( .A1(n515), .A2(n506), .ZN(n504) );
  XOR2_X1 U569 ( .A(G64GAT), .B(n504), .Z(G1333GAT) );
  NOR2_X1 U570 ( .A1(n560), .A2(n506), .ZN(n505) );
  XOR2_X1 U571 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  NOR2_X1 U572 ( .A1(n521), .A2(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n510), .A2(n509), .ZN(n520) );
  NOR2_X1 U576 ( .A1(n511), .A2(n520), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NOR2_X1 U580 ( .A1(n515), .A2(n520), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G92GAT), .B(KEYINPUT105), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1337GAT) );
  NOR2_X1 U583 ( .A1(n560), .A2(n520), .ZN(n518) );
  XOR2_X1 U584 ( .A(KEYINPUT106), .B(n518), .Z(n519) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n519), .ZN(G1338GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U587 ( .A(KEYINPUT44), .B(n522), .Z(n523) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  OR2_X1 U589 ( .A1(n524), .A2(n560), .ZN(n525) );
  NOR2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n535) );
  NAND2_X1 U591 ( .A1(n576), .A2(n535), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n529) );
  NAND2_X1 U594 ( .A1(n535), .A2(n563), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(G1341GAT) );
  NAND2_X1 U596 ( .A1(n580), .A2(n535), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n530), .B(KEYINPUT50), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n533) );
  XNOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U602 ( .A(KEYINPUT112), .B(n534), .Z(n537) );
  NAND2_X1 U603 ( .A1(n535), .A2(n570), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n543) );
  NOR2_X1 U606 ( .A1(n524), .A2(n538), .ZN(n539) );
  NAND2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(KEYINPUT115), .B(n541), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n553), .A2(n576), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  NAND2_X1 U612 ( .A1(n553), .A2(n563), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n546) );
  XNOR2_X1 U614 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n545) );
  XNOR2_X1 U615 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .Z(n547) );
  XNOR2_X1 U617 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  XOR2_X1 U619 ( .A(G155GAT), .B(KEYINPUT121), .Z(n552) );
  NAND2_X1 U620 ( .A1(n553), .A2(n580), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n552), .B(n551), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n570), .A2(n553), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n554), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  AND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(KEYINPUT55), .ZN(n572) );
  NOR2_X1 U627 ( .A1(n572), .A2(n560), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n576), .A2(n567), .ZN(n562) );
  XOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT123), .Z(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(G1348GAT) );
  XNOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n565) );
  NOR2_X1 U632 ( .A1(n292), .A2(n572), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(n566), .ZN(G1349GAT) );
  NAND2_X1 U635 ( .A1(n580), .A2(n567), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  OR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT58), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n578) );
  XNOR2_X1 U642 ( .A(n575), .B(KEYINPUT124), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n576), .A2(n581), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n586) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(G218GAT), .B(n587), .Z(G1355GAT) );
endmodule

