

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  INV_X1 U325 ( .A(KEYINPUT84), .ZN(n425) );
  XNOR2_X1 U326 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U327 ( .A(n449), .B(KEYINPUT106), .ZN(n522) );
  XNOR2_X1 U328 ( .A(n433), .B(n432), .ZN(n524) );
  XOR2_X1 U329 ( .A(n397), .B(n396), .Z(n517) );
  XOR2_X1 U330 ( .A(KEYINPUT10), .B(n357), .Z(n293) );
  XOR2_X1 U331 ( .A(G162GAT), .B(n380), .Z(n294) );
  XNOR2_X1 U332 ( .A(n458), .B(KEYINPUT45), .ZN(n459) );
  XNOR2_X1 U333 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U334 ( .A(n388), .B(G134GAT), .ZN(n389) );
  XNOR2_X1 U335 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U336 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U337 ( .A(n358), .B(n293), .ZN(n359) );
  XNOR2_X1 U338 ( .A(n476), .B(KEYINPUT121), .ZN(n477) );
  XNOR2_X1 U339 ( .A(n428), .B(n427), .ZN(n431) );
  XNOR2_X1 U340 ( .A(n360), .B(n359), .ZN(n538) );
  INV_X1 U341 ( .A(G106GAT), .ZN(n450) );
  INV_X1 U342 ( .A(G43GAT), .ZN(n455) );
  XNOR2_X1 U343 ( .A(KEYINPUT122), .B(G169GAT), .ZN(n480) );
  XNOR2_X1 U344 ( .A(n450), .B(KEYINPUT44), .ZN(n451) );
  XNOR2_X1 U345 ( .A(n455), .B(KEYINPUT40), .ZN(n456) );
  XNOR2_X1 U346 ( .A(n481), .B(n480), .ZN(G1348GAT) );
  XNOR2_X1 U347 ( .A(n457), .B(n456), .ZN(G1330GAT) );
  XOR2_X1 U348 ( .A(G50GAT), .B(G162GAT), .Z(n345) );
  XOR2_X1 U349 ( .A(KEYINPUT88), .B(KEYINPUT21), .Z(n296) );
  XNOR2_X1 U350 ( .A(G197GAT), .B(G218GAT), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n404) );
  XNOR2_X1 U352 ( .A(n345), .B(n404), .ZN(n297) );
  XOR2_X1 U353 ( .A(G22GAT), .B(G155GAT), .Z(n361) );
  XNOR2_X1 U354 ( .A(n297), .B(n361), .ZN(n302) );
  XNOR2_X1 U355 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n298), .B(KEYINPUT2), .ZN(n380) );
  XOR2_X1 U357 ( .A(n380), .B(KEYINPUT87), .Z(n300) );
  NAND2_X1 U358 ( .A1(G228GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U359 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U360 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U361 ( .A(G148GAT), .B(G106GAT), .Z(n304) );
  XNOR2_X1 U362 ( .A(G204GAT), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U364 ( .A(KEYINPUT69), .B(n305), .Z(n315) );
  XOR2_X1 U365 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n307) );
  XNOR2_X1 U366 ( .A(G211GAT), .B(KEYINPUT23), .ZN(n306) );
  XNOR2_X1 U367 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n315), .B(n308), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n475) );
  XOR2_X1 U370 ( .A(n475), .B(KEYINPUT28), .Z(n514) );
  INV_X1 U371 ( .A(G85GAT), .ZN(n314) );
  XOR2_X1 U372 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n312) );
  XNOR2_X1 U373 ( .A(G99GAT), .B(G92GAT), .ZN(n311) );
  XNOR2_X1 U374 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n346) );
  XNOR2_X1 U376 ( .A(n346), .B(n315), .ZN(n326) );
  XOR2_X1 U377 ( .A(G176GAT), .B(G64GAT), .Z(n413) );
  XOR2_X1 U378 ( .A(KEYINPUT68), .B(KEYINPUT31), .Z(n317) );
  XNOR2_X1 U379 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n316) );
  XNOR2_X1 U380 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U381 ( .A(n413), .B(n318), .Z(n320) );
  NAND2_X1 U382 ( .A1(G230GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U384 ( .A(n321), .B(KEYINPUT72), .Z(n324) );
  XNOR2_X1 U385 ( .A(G71GAT), .B(G57GAT), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n322), .B(KEYINPUT13), .ZN(n365) );
  XNOR2_X1 U387 ( .A(n365), .B(KEYINPUT33), .ZN(n323) );
  XNOR2_X1 U388 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U389 ( .A(n326), .B(n325), .ZN(n578) );
  XNOR2_X1 U390 ( .A(KEYINPUT41), .B(n578), .ZN(n550) );
  XOR2_X1 U391 ( .A(KEYINPUT100), .B(n550), .Z(n558) );
  XOR2_X1 U392 ( .A(G197GAT), .B(G141GAT), .Z(n328) );
  XNOR2_X1 U393 ( .A(G169GAT), .B(G15GAT), .ZN(n327) );
  XNOR2_X1 U394 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U395 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n330) );
  XNOR2_X1 U396 ( .A(G22GAT), .B(G8GAT), .ZN(n329) );
  XNOR2_X1 U397 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U398 ( .A(n332), .B(n331), .ZN(n343) );
  XOR2_X1 U399 ( .A(KEYINPUT66), .B(G1GAT), .Z(n362) );
  XOR2_X1 U400 ( .A(G113GAT), .B(G36GAT), .Z(n334) );
  XNOR2_X1 U401 ( .A(G43GAT), .B(G50GAT), .ZN(n333) );
  XNOR2_X1 U402 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U403 ( .A(n362), .B(n335), .Z(n337) );
  NAND2_X1 U404 ( .A1(G229GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U405 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U406 ( .A(n338), .B(KEYINPUT29), .Z(n341) );
  XNOR2_X1 U407 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n339) );
  XNOR2_X1 U408 ( .A(n339), .B(KEYINPUT7), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n347), .B(KEYINPUT67), .ZN(n340) );
  XNOR2_X1 U410 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U411 ( .A(n343), .B(n342), .ZN(n464) );
  NAND2_X1 U412 ( .A1(n558), .A2(n464), .ZN(n344) );
  XNOR2_X1 U413 ( .A(n344), .B(KEYINPUT101), .ZN(n504) );
  XOR2_X1 U414 ( .A(n346), .B(n345), .Z(n349) );
  XOR2_X1 U415 ( .A(G43GAT), .B(G134GAT), .Z(n420) );
  XNOR2_X1 U416 ( .A(n347), .B(n420), .ZN(n348) );
  XNOR2_X1 U417 ( .A(n349), .B(n348), .ZN(n360) );
  XOR2_X1 U418 ( .A(KEYINPUT73), .B(KEYINPUT9), .Z(n351) );
  XNOR2_X1 U419 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n350) );
  XNOR2_X1 U420 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U421 ( .A(G36GAT), .B(KEYINPUT75), .Z(n405) );
  XOR2_X1 U422 ( .A(n352), .B(n405), .Z(n354) );
  XNOR2_X1 U423 ( .A(G190GAT), .B(G218GAT), .ZN(n353) );
  XNOR2_X1 U424 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U425 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n356) );
  NAND2_X1 U426 ( .A1(G232GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U427 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n538), .B(KEYINPUT36), .ZN(n587) );
  XOR2_X1 U429 ( .A(G8GAT), .B(G211GAT), .Z(n412) );
  XOR2_X1 U430 ( .A(n412), .B(n361), .Z(n364) );
  XOR2_X1 U431 ( .A(G15GAT), .B(G127GAT), .Z(n419) );
  XNOR2_X1 U432 ( .A(n362), .B(n419), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n364), .B(n363), .ZN(n369) );
  XOR2_X1 U434 ( .A(n365), .B(KEYINPUT76), .Z(n367) );
  NAND2_X1 U435 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U437 ( .A(n369), .B(n368), .Z(n377) );
  XOR2_X1 U438 ( .A(KEYINPUT14), .B(G64GAT), .Z(n371) );
  XNOR2_X1 U439 ( .A(G183GAT), .B(G78GAT), .ZN(n370) );
  XNOR2_X1 U440 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U441 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n373) );
  XNOR2_X1 U442 ( .A(KEYINPUT12), .B(KEYINPUT77), .ZN(n372) );
  XNOR2_X1 U443 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U445 ( .A(n377), .B(n376), .ZN(n482) );
  XOR2_X1 U446 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n379) );
  XNOR2_X1 U447 ( .A(KEYINPUT91), .B(KEYINPUT5), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n397) );
  NAND2_X1 U449 ( .A1(G225GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n294), .B(n381), .ZN(n390) );
  XOR2_X1 U451 ( .A(G85GAT), .B(G148GAT), .Z(n383) );
  XNOR2_X1 U452 ( .A(G29GAT), .B(G127GAT), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U454 ( .A(KEYINPUT90), .B(G57GAT), .Z(n385) );
  XNOR2_X1 U455 ( .A(G1GAT), .B(G155GAT), .ZN(n384) );
  XNOR2_X1 U456 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U457 ( .A(n387), .B(n386), .Z(n388) );
  XOR2_X1 U458 ( .A(n391), .B(KEYINPUT6), .Z(n395) );
  XOR2_X1 U459 ( .A(G120GAT), .B(KEYINPUT79), .Z(n393) );
  XNOR2_X1 U460 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n392) );
  XNOR2_X1 U461 ( .A(n393), .B(n392), .ZN(n429) );
  XNOR2_X1 U462 ( .A(n429), .B(KEYINPUT89), .ZN(n394) );
  XNOR2_X1 U463 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U464 ( .A(G183GAT), .B(KEYINPUT19), .Z(n399) );
  XNOR2_X1 U465 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n398) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U467 ( .A(KEYINPUT18), .B(KEYINPUT82), .Z(n401) );
  XNOR2_X1 U468 ( .A(G190GAT), .B(KEYINPUT83), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U470 ( .A(n403), .B(n402), .Z(n433) );
  XOR2_X1 U471 ( .A(n405), .B(n404), .Z(n407) );
  NAND2_X1 U472 ( .A1(G226GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U473 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U474 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n409) );
  XNOR2_X1 U475 ( .A(G204GAT), .B(G92GAT), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U477 ( .A(n411), .B(n410), .Z(n415) );
  XNOR2_X1 U478 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U479 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n433), .B(n416), .ZN(n520) );
  XNOR2_X1 U481 ( .A(KEYINPUT27), .B(n520), .ZN(n437) );
  NOR2_X1 U482 ( .A1(n517), .A2(n437), .ZN(n543) );
  NAND2_X1 U483 ( .A1(n543), .A2(n514), .ZN(n525) );
  XOR2_X1 U484 ( .A(KEYINPUT85), .B(KEYINPUT80), .Z(n418) );
  XNOR2_X1 U485 ( .A(G176GAT), .B(G71GAT), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n418), .B(n417), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U488 ( .A(KEYINPUT20), .B(G99GAT), .Z(n421) );
  XNOR2_X1 U489 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U490 ( .A(n424), .B(n423), .Z(n428) );
  NAND2_X1 U491 ( .A1(G227GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n429), .B(KEYINPUT81), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U494 ( .A(KEYINPUT86), .B(n524), .Z(n434) );
  NOR2_X1 U495 ( .A1(n525), .A2(n434), .ZN(n435) );
  XOR2_X1 U496 ( .A(KEYINPUT94), .B(n435), .Z(n445) );
  NAND2_X1 U497 ( .A1(n524), .A2(n475), .ZN(n436) );
  XOR2_X1 U498 ( .A(KEYINPUT26), .B(n436), .Z(n571) );
  INV_X1 U499 ( .A(n437), .ZN(n438) );
  NAND2_X1 U500 ( .A1(n571), .A2(n438), .ZN(n442) );
  NOR2_X1 U501 ( .A1(n524), .A2(n520), .ZN(n439) );
  NOR2_X1 U502 ( .A1(n475), .A2(n439), .ZN(n440) );
  XNOR2_X1 U503 ( .A(n440), .B(KEYINPUT25), .ZN(n441) );
  NAND2_X1 U504 ( .A1(n442), .A2(n441), .ZN(n443) );
  NAND2_X1 U505 ( .A1(n517), .A2(n443), .ZN(n444) );
  NAND2_X1 U506 ( .A1(n445), .A2(n444), .ZN(n485) );
  NAND2_X1 U507 ( .A1(n482), .A2(n485), .ZN(n446) );
  XOR2_X1 U508 ( .A(KEYINPUT99), .B(n446), .Z(n447) );
  NOR2_X1 U509 ( .A1(n587), .A2(n447), .ZN(n448) );
  XOR2_X1 U510 ( .A(KEYINPUT37), .B(n448), .Z(n453) );
  NAND2_X1 U511 ( .A1(n504), .A2(n453), .ZN(n449) );
  NOR2_X1 U512 ( .A1(n514), .A2(n522), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(G1339GAT) );
  NOR2_X1 U514 ( .A1(n464), .A2(n578), .ZN(n486) );
  NAND2_X1 U515 ( .A1(n453), .A2(n486), .ZN(n454) );
  XNOR2_X1 U516 ( .A(KEYINPUT38), .B(n454), .ZN(n501) );
  NOR2_X1 U517 ( .A1(n501), .A2(n524), .ZN(n457) );
  INV_X1 U518 ( .A(n464), .ZN(n572) );
  NOR2_X1 U519 ( .A1(n482), .A2(n587), .ZN(n460) );
  INV_X1 U520 ( .A(KEYINPUT110), .ZN(n458) );
  NOR2_X1 U521 ( .A1(n578), .A2(n461), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT111), .ZN(n463) );
  NOR2_X1 U523 ( .A1(n463), .A2(n572), .ZN(n471) );
  XOR2_X1 U524 ( .A(KEYINPUT47), .B(KEYINPUT109), .Z(n469) );
  XOR2_X1 U525 ( .A(KEYINPUT108), .B(n482), .Z(n563) );
  NOR2_X1 U526 ( .A1(n464), .A2(n550), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n465), .B(KEYINPUT46), .ZN(n466) );
  NOR2_X1 U528 ( .A1(n563), .A2(n466), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n467), .A2(n538), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U531 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n472), .B(KEYINPUT48), .ZN(n545) );
  NOR2_X1 U533 ( .A1(n520), .A2(n545), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n473), .B(KEYINPUT54), .ZN(n474) );
  NAND2_X1 U535 ( .A1(n474), .A2(n517), .ZN(n569) );
  NOR2_X1 U536 ( .A1(n475), .A2(n569), .ZN(n478) );
  INV_X1 U537 ( .A(KEYINPUT55), .ZN(n476) );
  NOR2_X1 U538 ( .A1(n524), .A2(n479), .ZN(n566) );
  NAND2_X1 U539 ( .A1(n572), .A2(n566), .ZN(n481) );
  INV_X1 U540 ( .A(n482), .ZN(n582) );
  NAND2_X1 U541 ( .A1(n538), .A2(n582), .ZN(n483) );
  XOR2_X1 U542 ( .A(KEYINPUT16), .B(n483), .Z(n484) );
  AND2_X1 U543 ( .A1(n485), .A2(n484), .ZN(n503) );
  NAND2_X1 U544 ( .A1(n486), .A2(n503), .ZN(n495) );
  NOR2_X1 U545 ( .A1(n517), .A2(n495), .ZN(n488) );
  XNOR2_X1 U546 ( .A(KEYINPUT34), .B(KEYINPUT95), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(n489), .ZN(G1324GAT) );
  NOR2_X1 U549 ( .A1(n520), .A2(n495), .ZN(n490) );
  XOR2_X1 U550 ( .A(G8GAT), .B(n490), .Z(G1325GAT) );
  NOR2_X1 U551 ( .A1(n495), .A2(n524), .ZN(n494) );
  XOR2_X1 U552 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n492) );
  XNOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NOR2_X1 U556 ( .A1(n514), .A2(n495), .ZN(n496) );
  XOR2_X1 U557 ( .A(KEYINPUT98), .B(n496), .Z(n497) );
  XNOR2_X1 U558 ( .A(G22GAT), .B(n497), .ZN(G1327GAT) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  NOR2_X1 U560 ( .A1(n501), .A2(n517), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U562 ( .A1(n501), .A2(n520), .ZN(n500) );
  XOR2_X1 U563 ( .A(G36GAT), .B(n500), .Z(G1329GAT) );
  NOR2_X1 U564 ( .A1(n514), .A2(n501), .ZN(n502) );
  XOR2_X1 U565 ( .A(G50GAT), .B(n502), .Z(G1331GAT) );
  NAND2_X1 U566 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U567 ( .A(KEYINPUT102), .B(n505), .ZN(n513) );
  NOR2_X1 U568 ( .A1(n517), .A2(n513), .ZN(n506) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n506), .Z(n507) );
  XNOR2_X1 U570 ( .A(KEYINPUT42), .B(n507), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n513), .A2(n520), .ZN(n509) );
  XNOR2_X1 U572 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G64GAT), .B(n510), .ZN(G1333GAT) );
  NOR2_X1 U575 ( .A1(n513), .A2(n524), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(G1334GAT) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  NOR2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NOR2_X1 U581 ( .A1(n522), .A2(n517), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(KEYINPUT107), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  NOR2_X1 U584 ( .A1(n522), .A2(n520), .ZN(n521) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n521), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n524), .ZN(n523) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n523), .Z(G1338GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n530) );
  INV_X1 U589 ( .A(n524), .ZN(n527) );
  NOR2_X1 U590 ( .A1(n525), .A2(n545), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U592 ( .A(KEYINPUT112), .B(n528), .Z(n539) );
  NAND2_X1 U593 ( .A1(n539), .A2(n572), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U597 ( .A1(n539), .A2(n558), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n537) );
  XOR2_X1 U600 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n535) );
  NAND2_X1 U601 ( .A1(n563), .A2(n539), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n541) );
  INV_X1 U605 ( .A(n538), .ZN(n565) );
  NAND2_X1 U606 ( .A1(n539), .A2(n565), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U608 ( .A(G134GAT), .B(n542), .Z(G1343GAT) );
  NAND2_X1 U609 ( .A1(n543), .A2(n571), .ZN(n544) );
  NOR2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n572), .A2(n554), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n548) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n552) );
  INV_X1 U616 ( .A(n554), .ZN(n549) );
  NOR2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(n552), .B(n551), .Z(G1345GAT) );
  NAND2_X1 U619 ( .A1(n582), .A2(n554), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n556) );
  NAND2_X1 U622 ( .A1(n554), .A2(n565), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n566), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT123), .Z(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n562) );
  XOR2_X1 U628 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n574) );
  INV_X1 U636 ( .A(n569), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n586) );
  INV_X1 U638 ( .A(n586), .ZN(n583) );
  NAND2_X1 U639 ( .A1(n583), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(n575), .B(KEYINPUT59), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n580) );
  NAND2_X1 U645 ( .A1(n583), .A2(n578), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  XOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT127), .Z(n585) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

