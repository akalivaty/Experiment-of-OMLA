//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(KEYINPUT22), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n205), .B1(new_n212), .B2(KEYINPUT29), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT74), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(G148gat), .ZN(new_n216));
  INV_X1    g015(.A(G148gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(KEYINPUT74), .A3(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(G148gat), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT75), .A4(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n216), .A2(new_n219), .A3(new_n218), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT75), .ZN(new_n222));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  OR3_X1    g022(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n221), .A2(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT73), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n217), .A2(G141gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n215), .A2(G148gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n217), .A2(G141gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n219), .A2(new_n230), .A3(KEYINPUT73), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n223), .A2(KEYINPUT2), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n223), .A2(KEYINPUT72), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n223), .A2(KEYINPUT72), .ZN(new_n235));
  INV_X1    g034(.A(G155gat), .ZN(new_n236));
  INV_X1    g035(.A(G162gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n220), .A2(new_n225), .B1(new_n233), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n213), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(KEYINPUT76), .A3(new_n205), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n233), .A2(new_n239), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n221), .A2(new_n222), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n223), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n220), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(new_n247), .A3(new_n205), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT76), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT29), .B1(new_n243), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n212), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n242), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G228gat), .ZN(new_n254));
  INV_X1    g053(.A(G233gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n256), .B(new_n242), .C1(new_n251), .C2(new_n252), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n204), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(G22gat), .B1(new_n260), .B2(KEYINPUT83), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n260), .A2(KEYINPUT83), .A3(G22gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n259), .ZN(new_n264));
  INV_X1    g063(.A(new_n204), .ZN(new_n265));
  OAI22_X1  g064(.A1(new_n262), .A2(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n263), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n264), .A2(new_n265), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(new_n268), .A3(new_n261), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G226gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(new_n255), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(KEYINPUT29), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT26), .ZN(new_n277));
  INV_X1    g076(.A(G169gat), .ZN(new_n278));
  INV_X1    g077(.A(G176gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n277), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n279), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n276), .A2(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  NOR3_X1   g085(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT67), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n275), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  OAI211_X1 g089(.A(KEYINPUT66), .B(new_n289), .C1(new_n290), .C2(KEYINPUT27), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT27), .ZN(new_n294));
  AOI21_X1  g093(.A(G190gat), .B1(new_n294), .B2(G183gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n290), .A2(KEYINPUT27), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n291), .A2(new_n295), .A3(new_n292), .A4(new_n296), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n288), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n286), .A2(KEYINPUT23), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  AND4_X1   g104(.A1(new_n302), .A2(new_n303), .A3(new_n281), .A4(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n275), .A2(KEYINPUT24), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(G183gat), .A3(G190gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n290), .A2(new_n289), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT65), .ZN(new_n312));
  OR3_X1    g111(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n307), .A2(new_n309), .B1(new_n290), .B2(new_n289), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n303), .A2(new_n281), .A3(new_n305), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT25), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT70), .B1(new_n301), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n303), .A2(new_n281), .A3(new_n305), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n310), .A2(new_n311), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n323), .A2(KEYINPUT25), .B1(new_n314), .B2(new_n306), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n282), .A2(new_n276), .A3(new_n283), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n285), .A2(new_n286), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT67), .B1(new_n286), .B2(new_n277), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n329), .A2(new_n298), .A3(new_n275), .A4(new_n299), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n324), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n274), .B1(new_n320), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n318), .A3(new_n315), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n333), .A2(new_n271), .A3(new_n255), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n252), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(G8gat), .B(G36gat), .Z(new_n336));
  XOR2_X1   g135(.A(G64gat), .B(G92gat), .Z(new_n337));
  XOR2_X1   g136(.A(new_n336), .B(new_n337), .Z(new_n338));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n272), .A3(new_n331), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n333), .A2(new_n273), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n212), .A3(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n335), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n338), .B(KEYINPUT71), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n335), .B2(new_n341), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT30), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n335), .A2(new_n338), .A3(new_n341), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT30), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(G127gat), .A2(G134gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT68), .ZN(new_n352));
  NAND2_X1  g151(.A1(G127gat), .A2(G134gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(G127gat), .A2(G134gat), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT68), .B1(new_n355), .B2(new_n350), .ZN(new_n356));
  INV_X1    g155(.A(G113gat), .ZN(new_n357));
  INV_X1    g156(.A(G120gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n360));
  NAND2_X1  g159(.A1(G113gat), .A2(G120gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n354), .A2(new_n356), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n355), .A2(new_n350), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT1), .B1(new_n357), .B2(new_n358), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n364), .A2(new_n352), .A3(new_n361), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n333), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT64), .ZN(new_n370));
  INV_X1    g169(.A(new_n367), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n324), .A2(new_n371), .A3(new_n330), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT32), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT33), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G15gat), .B(G43gat), .Z(new_n377));
  XNOR2_X1  g176(.A(G71gat), .B(G99gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n374), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n379), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n373), .B(KEYINPUT32), .C1(new_n375), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT34), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n372), .ZN(new_n385));
  INV_X1    g184(.A(new_n370), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI211_X1 g186(.A(KEYINPUT34), .B(new_n370), .C1(new_n368), .C2(new_n372), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n383), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n380), .A3(new_n382), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n349), .A2(KEYINPUT35), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n270), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT6), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n243), .A2(new_n250), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n371), .B1(new_n240), .B2(new_n205), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT77), .B(KEYINPUT5), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n244), .A2(new_n247), .A3(new_n367), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT4), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT81), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT80), .B1(new_n406), .B2(KEYINPUT4), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n409), .B2(new_n411), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n400), .B(new_n405), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n244), .A2(new_n247), .A3(new_n367), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n404), .B1(new_n417), .B2(new_n407), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n367), .B1(new_n244), .B2(new_n247), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n404), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n421), .A2(new_n402), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G57gat), .B(G85gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT79), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n428), .B(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n396), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n428), .B(new_n429), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT84), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT84), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n414), .B2(new_n423), .ZN(new_n438));
  OR3_X1    g237(.A1(new_n432), .A2(KEYINPUT87), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT6), .A3(new_n431), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT87), .B1(new_n432), .B2(new_n438), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n395), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n444));
  AOI211_X1 g243(.A(new_n396), .B(new_n433), .C1(new_n414), .C2(new_n423), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n398), .B1(new_n250), .B2(new_n243), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT80), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(new_n415), .B2(new_n416), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n406), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT81), .B1(new_n406), .B2(KEYINPUT4), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n453), .A2(new_n405), .B1(new_n419), .B2(new_n422), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT6), .B1(new_n454), .B2(new_n433), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n424), .A2(new_n431), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n445), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n444), .B1(new_n457), .B2(new_n349), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n454), .A2(new_n433), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n440), .B1(new_n432), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n349), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(KEYINPUT82), .A3(new_n461), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n391), .A2(new_n392), .B1(KEYINPUT69), .B2(new_n383), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n383), .A2(KEYINPUT69), .A3(new_n389), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n270), .A2(new_n458), .A3(new_n462), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT35), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n443), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n458), .A2(new_n462), .B1(new_n269), .B2(new_n266), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT36), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n383), .A2(KEYINPUT69), .ZN(new_n472));
  INV_X1    g271(.A(new_n392), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n389), .B1(new_n380), .B2(new_n382), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n471), .B1(new_n475), .B2(new_n464), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n393), .A2(KEYINPUT36), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n470), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n438), .B1(new_n345), .B2(new_n348), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n400), .B1(new_n412), .B2(new_n413), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT39), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n404), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n415), .A2(new_n420), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(new_n403), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n453), .B2(new_n403), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n485), .A3(new_n437), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n487), .A2(KEYINPUT40), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n488), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n482), .A2(new_n485), .A3(new_n437), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n479), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT86), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n479), .A2(new_n489), .A3(KEYINPUT86), .A4(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT37), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n335), .A2(new_n497), .A3(new_n341), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n212), .B1(new_n332), .B2(new_n334), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n339), .A2(new_n252), .A3(new_n340), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(KEYINPUT37), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n343), .A2(KEYINPUT38), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n503), .A2(new_n346), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n333), .A2(KEYINPUT70), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n325), .B1(new_n324), .B2(new_n330), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n273), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n334), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n212), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n339), .A2(new_n212), .A3(new_n340), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT37), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n338), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(KEYINPUT88), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT88), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n497), .B1(new_n335), .B2(new_n341), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(new_n338), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n516), .A3(new_n498), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT38), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n517), .B2(KEYINPUT38), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n504), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n496), .B(new_n270), .C1(new_n442), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n478), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n469), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT93), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G1gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n527), .A3(G1gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT16), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(G8gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n536));
  XOR2_X1   g335(.A(G43gat), .B(G50gat), .Z(new_n537));
  INV_X1    g336(.A(KEYINPUT15), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT91), .B(G29gat), .ZN(new_n540));
  OR3_X1    g339(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n540), .A2(G36gat), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n537), .A2(new_n538), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n535), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n546), .B(KEYINPUT17), .ZN(new_n550));
  INV_X1    g349(.A(new_n535), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT18), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(KEYINPUT18), .A3(new_n554), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n549), .B1(new_n535), .B2(new_n546), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n554), .B(KEYINPUT13), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G113gat), .B(G141gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(G169gat), .B(G197gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n567), .B(KEYINPUT12), .Z(new_n568));
  XOR2_X1   g367(.A(new_n562), .B(new_n568), .Z(new_n569));
  NOR2_X1   g368(.A1(new_n525), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  OR2_X1    g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT9), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G57gat), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT95), .B1(new_n575), .B2(G64gat), .ZN(new_n576));
  INV_X1    g375(.A(G64gat), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(G57gat), .B2(new_n577), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n575), .A2(KEYINPUT95), .A3(G64gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n574), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT96), .Z(new_n581));
  XNOR2_X1  g380(.A(G57gat), .B(G64gat), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n571), .B(new_n572), .C1(new_n582), .C2(new_n573), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G127gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n551), .B1(new_n584), .B2(new_n585), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(G155gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT99), .B(KEYINPUT7), .ZN(new_n601));
  INV_X1    g400(.A(G85gat), .ZN(new_n602));
  INV_X1    g401(.A(G92gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  AOI22_X1  g406(.A1(KEYINPUT8), .A2(new_n607), .B1(new_n602), .B2(new_n603), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G99gat), .B(G106gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n550), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n611), .ZN(new_n613));
  AND2_X1   g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n613), .A2(new_n546), .B1(KEYINPUT41), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT100), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n614), .A2(KEYINPUT41), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT97), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT98), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n617), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(G190gat), .B(G218gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n584), .A2(new_n611), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(KEYINPUT101), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT10), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n584), .A2(new_n611), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n629), .A2(KEYINPUT10), .ZN(new_n634));
  OR3_X1    g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n631), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n633), .B1(new_n636), .B2(new_n628), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n600), .A2(new_n627), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n570), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n460), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n529), .ZN(G1324gat));
  NOR2_X1   g447(.A1(new_n646), .A2(new_n461), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT42), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT102), .Z(new_n654));
  INV_X1    g453(.A(G8gat), .ZN(new_n655));
  OAI221_X1 g454(.A(new_n654), .B1(new_n652), .B2(new_n651), .C1(new_n655), .C2(new_n649), .ZN(G1325gat));
  INV_X1    g455(.A(new_n646), .ZN(new_n657));
  INV_X1    g456(.A(new_n393), .ZN(new_n658));
  AOI21_X1  g457(.A(G15gat), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT103), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT104), .B1(new_n476), .B2(new_n477), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT36), .B1(new_n463), .B2(new_n465), .ZN(new_n662));
  INV_X1    g461(.A(new_n477), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n666), .A2(G15gat), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n660), .B1(new_n657), .B2(new_n667), .ZN(G1326gat));
  NOR2_X1   g467(.A1(new_n646), .A2(new_n270), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n524), .B2(new_n627), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n442), .A2(new_n395), .B1(new_n467), .B2(KEYINPUT35), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n470), .A2(new_n666), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n522), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n676), .A2(new_n522), .A3(KEYINPUT106), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n627), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(KEYINPUT44), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n674), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n676), .A2(new_n522), .A3(KEYINPUT106), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT106), .B1(new_n676), .B2(new_n522), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n469), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(KEYINPUT107), .A3(new_n683), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n673), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n569), .A2(KEYINPUT105), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n569), .A2(KEYINPUT105), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n599), .A2(new_n644), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT108), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n673), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n688), .A2(KEYINPUT107), .A3(new_n683), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT107), .B1(new_n688), .B2(new_n683), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n701));
  INV_X1    g500(.A(new_n695), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n696), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n540), .B1(new_n705), .B2(new_n460), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n570), .A2(new_n627), .A3(new_n694), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n460), .A2(new_n540), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT45), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(new_n711), .ZN(G1328gat));
  INV_X1    g511(.A(G36gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n707), .A2(new_n713), .A3(new_n349), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT109), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT46), .ZN(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n705), .B2(new_n461), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1329gat));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719));
  INV_X1    g518(.A(G43gat), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n690), .A2(new_n695), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n721), .B2(new_n666), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n707), .A2(new_n720), .A3(new_n658), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT47), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n696), .A2(new_n703), .A3(new_n666), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(new_n726), .A3(G43gat), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n723), .A2(KEYINPUT47), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n726), .B1(new_n725), .B2(G43gat), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n719), .B(new_n724), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n725), .A2(G43gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT110), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(new_n727), .A3(new_n728), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n719), .B1(new_n735), .B2(new_n724), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n732), .A2(new_n736), .ZN(G1330gat));
  INV_X1    g536(.A(G50gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n270), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n707), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n690), .A2(new_n270), .A3(new_n695), .ZN(new_n741));
  OAI211_X1 g540(.A(KEYINPUT48), .B(new_n740), .C1(new_n741), .C2(new_n738), .ZN(new_n742));
  INV_X1    g541(.A(new_n740), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n704), .A2(new_n739), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(G50gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(G1331gat));
  INV_X1    g546(.A(new_n644), .ZN(new_n748));
  NOR4_X1   g547(.A1(new_n693), .A2(new_n600), .A3(new_n627), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n688), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n460), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(new_n575), .ZN(G1332gat));
  INV_X1    g551(.A(new_n750), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n461), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT113), .Z(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1333gat));
  NOR3_X1   g557(.A1(new_n750), .A2(G71gat), .A3(new_n393), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n753), .A2(new_n666), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n759), .B1(G71gat), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n753), .A2(new_n739), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g563(.A1(new_n693), .A2(new_n599), .A3(new_n748), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n700), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G85gat), .B1(new_n767), .B2(new_n460), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n693), .A2(new_n599), .A3(new_n682), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(new_n688), .A3(KEYINPUT51), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  OR2_X1    g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n769), .A2(new_n688), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n772), .B(new_n773), .C1(KEYINPUT51), .C2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n748), .B1(new_n775), .B2(KEYINPUT115), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(KEYINPUT115), .B2(new_n775), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n457), .A2(new_n602), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n768), .B1(new_n777), .B2(new_n778), .ZN(G1336gat));
  AOI21_X1  g578(.A(new_n603), .B1(new_n766), .B2(new_n349), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n774), .A2(KEYINPUT116), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT51), .Z(new_n782));
  NOR3_X1   g581(.A1(new_n748), .A2(G92gat), .A3(new_n461), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n775), .A2(new_n783), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n785), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n784), .A2(new_n785), .B1(new_n780), .B2(new_n787), .ZN(G1337gat));
  INV_X1    g587(.A(new_n666), .ZN(new_n789));
  OAI21_X1  g588(.A(G99gat), .B1(new_n767), .B2(new_n789), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n393), .A2(G99gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n777), .B2(new_n791), .ZN(G1338gat));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n766), .B2(new_n739), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n748), .A2(new_n270), .A3(G106gat), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n782), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n775), .A2(new_n795), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n797), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n796), .A2(new_n797), .B1(new_n794), .B2(new_n799), .ZN(G1339gat));
  NAND3_X1  g599(.A1(new_n645), .A2(new_n692), .A3(new_n691), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n633), .B1(new_n632), .B2(new_n634), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n635), .A2(KEYINPUT54), .A3(new_n802), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n803), .B(new_n641), .C1(KEYINPUT54), .C2(new_n635), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n642), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n691), .B2(new_n692), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n562), .A2(new_n568), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n553), .A2(new_n554), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n559), .A2(new_n560), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n567), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n644), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n814), .B(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n682), .B1(new_n809), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n627), .A2(new_n810), .A3(new_n813), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n818), .A2(new_n808), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(KEYINPUT118), .B(new_n801), .C1(new_n820), .C2(new_n599), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n599), .B1(new_n817), .B2(new_n819), .ZN(new_n823));
  INV_X1    g622(.A(new_n801), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n460), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(new_n270), .A3(new_n466), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n349), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n693), .A2(new_n357), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT119), .Z(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n826), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n460), .A2(new_n349), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n833), .A2(new_n270), .A3(new_n658), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(G113gat), .B1(new_n835), .B2(new_n569), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n832), .A2(new_n836), .ZN(G1340gat));
  OAI21_X1  g636(.A(G120gat), .B1(new_n835), .B2(new_n748), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT120), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n840), .B(G120gat), .C1(new_n835), .C2(new_n748), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n644), .A2(new_n358), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT121), .Z(new_n844));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n845), .ZN(G1341gat));
  NAND3_X1  g645(.A1(new_n829), .A2(new_n589), .A3(new_n599), .ZN(new_n847));
  OAI21_X1  g646(.A(G127gat), .B1(new_n835), .B2(new_n600), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1342gat));
  NOR2_X1   g648(.A1(new_n682), .A2(new_n349), .ZN(new_n850));
  INV_X1    g649(.A(G134gat), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OR3_X1    g651(.A1(new_n828), .A2(KEYINPUT56), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n835), .B2(new_n682), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT56), .B1(new_n828), .B2(new_n852), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(G1343gat));
  NOR2_X1   g655(.A1(new_n666), .A2(new_n270), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NOR4_X1   g657(.A1(new_n826), .A2(new_n460), .A3(new_n349), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n569), .A2(G141gat), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT58), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n270), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n814), .B1(new_n808), .B2(new_n569), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n682), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n599), .B1(new_n865), .B2(new_n819), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n863), .B1(new_n866), .B2(new_n824), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n821), .A2(new_n739), .A3(new_n825), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(new_n862), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n789), .A2(new_n834), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n870), .A2(new_n569), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n861), .B1(new_n872), .B2(new_n215), .ZN(new_n873));
  INV_X1    g672(.A(new_n870), .ZN(new_n874));
  INV_X1    g673(.A(new_n871), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n693), .A3(new_n875), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n876), .A2(G141gat), .B1(new_n859), .B2(new_n860), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n873), .B1(new_n877), .B2(new_n878), .ZN(G1344gat));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  AOI211_X1 g679(.A(new_n880), .B(G148gat), .C1(new_n859), .C2(new_n644), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n821), .A2(new_n825), .A3(new_n863), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n866), .B1(new_n569), .B2(new_n645), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n862), .B1(new_n883), .B2(new_n270), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886));
  AOI211_X1 g685(.A(new_n880), .B(new_n748), .C1(new_n871), .C2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n885), .B(new_n887), .C1(new_n886), .C2(new_n871), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n870), .A2(new_n748), .A3(new_n871), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(KEYINPUT59), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n881), .B1(new_n890), .B2(G148gat), .ZN(G1345gat));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n875), .ZN(new_n892));
  OAI21_X1  g691(.A(G155gat), .B1(new_n892), .B2(new_n600), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n859), .A2(new_n236), .A3(new_n599), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1346gat));
  OAI21_X1  g694(.A(G162gat), .B1(new_n892), .B2(new_n682), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n827), .A2(new_n237), .A3(new_n850), .A4(new_n857), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1347gat));
  NOR3_X1   g697(.A1(new_n457), .A2(new_n461), .A3(new_n393), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n821), .A2(new_n825), .A3(new_n270), .A4(new_n899), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(new_n278), .A3(new_n569), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n270), .A2(new_n349), .A3(new_n466), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n821), .A2(new_n825), .A3(new_n460), .A4(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT123), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n693), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n901), .B1(new_n905), .B2(new_n278), .ZN(G1348gat));
  NOR2_X1   g705(.A1(new_n748), .A2(G176gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n900), .A2(new_n748), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n908), .B(new_n909), .C1(new_n279), .C2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n903), .A2(new_n912), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n913), .A2(new_n914), .A3(new_n907), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n910), .A2(new_n279), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT124), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n911), .A2(new_n917), .ZN(G1349gat));
  NOR2_X1   g717(.A1(new_n290), .A2(KEYINPUT27), .ZN(new_n919));
  INV_X1    g718(.A(new_n296), .ZN(new_n920));
  OR4_X1    g719(.A1(new_n919), .A2(new_n903), .A3(new_n920), .A4(new_n600), .ZN(new_n921));
  OAI21_X1  g720(.A(G183gat), .B1(new_n900), .B2(new_n600), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n924));
  NAND2_X1  g723(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n921), .A2(new_n925), .A3(new_n922), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n900), .B2(new_n682), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT61), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n682), .A2(G190gat), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n904), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n904), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(G1351gat));
  NOR4_X1   g733(.A1(new_n826), .A2(new_n457), .A3(new_n461), .A4(new_n858), .ZN(new_n935));
  AOI21_X1  g734(.A(G197gat), .B1(new_n935), .B2(new_n693), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n457), .A2(new_n461), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n789), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n938), .B1(new_n882), .B2(new_n884), .ZN(new_n939));
  INV_X1    g738(.A(G197gat), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n569), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n936), .B1(new_n939), .B2(new_n941), .ZN(G1352gat));
  XOR2_X1   g741(.A(KEYINPUT127), .B(G204gat), .Z(new_n943));
  NAND2_X1  g742(.A1(new_n644), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n935), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n948));
  INV_X1    g747(.A(new_n939), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(new_n748), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n947), .B(new_n948), .C1(new_n950), .C2(new_n943), .ZN(G1353gat));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n207), .A3(new_n599), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n939), .A2(new_n599), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n953), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n953), .B2(G211gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(G1354gat));
  OAI21_X1  g755(.A(G218gat), .B1(new_n949), .B2(new_n682), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n935), .A2(new_n208), .A3(new_n627), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1355gat));
endmodule


