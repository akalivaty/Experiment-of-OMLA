

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U553 ( .A1(n681), .A2(n992), .ZN(n690) );
  INV_X1 U554 ( .A(n842), .ZN(n984) );
  INV_X2 U555 ( .A(n520), .ZN(n879) );
  BUF_X1 U556 ( .A(n545), .Z(n527) );
  NOR2_X1 U557 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  NAND2_X2 U558 ( .A1(n761), .A2(n680), .ZN(n727) );
  NOR2_X2 U559 ( .A1(n554), .A2(n553), .ZN(G160) );
  INV_X1 U560 ( .A(KEYINPUT64), .ZN(n754) );
  INV_X1 U561 ( .A(KEYINPUT33), .ZN(n756) );
  INV_X1 U562 ( .A(G2104), .ZN(n525) );
  NOR2_X1 U563 ( .A1(n531), .A2(n530), .ZN(G164) );
  XOR2_X1 U564 ( .A(KEYINPUT17), .B(n519), .Z(n547) );
  INV_X1 U565 ( .A(n547), .ZN(n520) );
  NAND2_X1 U566 ( .A1(n879), .A2(G138), .ZN(n521) );
  XNOR2_X1 U567 ( .A(n521), .B(KEYINPUT84), .ZN(n523) );
  AND2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n882) );
  NAND2_X1 U569 ( .A1(G114), .A2(n882), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n531) );
  NAND2_X1 U571 ( .A1(n525), .A2(G2105), .ZN(n524) );
  XNOR2_X2 U572 ( .A(n524), .B(KEYINPUT65), .ZN(n884) );
  NAND2_X1 U573 ( .A1(n884), .A2(G126), .ZN(n529) );
  NOR2_X1 U574 ( .A1(n525), .A2(G2105), .ZN(n526) );
  XNOR2_X1 U575 ( .A(n526), .B(KEYINPUT66), .ZN(n545) );
  NAND2_X1 U576 ( .A1(G102), .A2(n527), .ZN(n528) );
  NAND2_X1 U577 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n643) );
  NAND2_X1 U579 ( .A1(n643), .A2(G89), .ZN(n532) );
  XNOR2_X1 U580 ( .A(n532), .B(KEYINPUT4), .ZN(n534) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n618) );
  XOR2_X1 U582 ( .A(G651), .B(KEYINPUT68), .Z(n537) );
  NOR2_X2 U583 ( .A1(n618), .A2(n537), .ZN(n644) );
  NAND2_X1 U584 ( .A1(G76), .A2(n644), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U586 ( .A(KEYINPUT5), .B(n535), .ZN(n543) );
  NOR2_X2 U587 ( .A1(G651), .A2(n618), .ZN(n648) );
  NAND2_X1 U588 ( .A1(n648), .A2(G51), .ZN(n536) );
  XOR2_X1 U589 ( .A(KEYINPUT73), .B(n536), .Z(n540) );
  NOR2_X1 U590 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n538), .Z(n573) );
  BUF_X1 U592 ( .A(n573), .Z(n649) );
  NAND2_X1 U593 ( .A1(G63), .A2(n649), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U595 ( .A(KEYINPUT6), .B(n541), .Z(n542) );
  NAND2_X1 U596 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U597 ( .A(KEYINPUT7), .B(n544), .ZN(G168) );
  XOR2_X1 U598 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U599 ( .A1(n545), .A2(G101), .ZN(n546) );
  XOR2_X1 U600 ( .A(KEYINPUT23), .B(n546), .Z(n550) );
  NAND2_X1 U601 ( .A1(n547), .A2(G137), .ZN(n548) );
  XOR2_X1 U602 ( .A(KEYINPUT67), .B(n548), .Z(n549) );
  NAND2_X1 U603 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U604 ( .A1(G125), .A2(n884), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G113), .A2(n882), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n553) );
  AND2_X1 U607 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  NAND2_X1 U611 ( .A1(G7), .A2(G661), .ZN(n555) );
  XOR2_X1 U612 ( .A(n555), .B(KEYINPUT10), .Z(n927) );
  NAND2_X1 U613 ( .A1(n927), .A2(G567), .ZN(n556) );
  XOR2_X1 U614 ( .A(KEYINPUT11), .B(n556), .Z(G234) );
  NAND2_X1 U615 ( .A1(n573), .A2(G56), .ZN(n557) );
  XOR2_X1 U616 ( .A(KEYINPUT14), .B(n557), .Z(n563) );
  NAND2_X1 U617 ( .A1(n643), .A2(G81), .ZN(n558) );
  XNOR2_X1 U618 ( .A(n558), .B(KEYINPUT12), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G68), .A2(n644), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U621 ( .A(KEYINPUT13), .B(n561), .Z(n562) );
  NOR2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n648), .A2(G43), .ZN(n564) );
  NAND2_X1 U624 ( .A1(n565), .A2(n564), .ZN(n992) );
  INV_X1 U625 ( .A(G860), .ZN(n594) );
  OR2_X1 U626 ( .A1(n992), .A2(n594), .ZN(G153) );
  NAND2_X1 U627 ( .A1(n643), .A2(G90), .ZN(n567) );
  NAND2_X1 U628 ( .A1(G77), .A2(n644), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U630 ( .A(KEYINPUT9), .B(n568), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n649), .A2(G64), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n648), .A2(G52), .ZN(n569) );
  AND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n571), .ZN(G301) );
  NAND2_X1 U635 ( .A1(n643), .A2(G92), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G66), .A2(n573), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U638 ( .A1(n648), .A2(G54), .ZN(n577) );
  NAND2_X1 U639 ( .A1(G79), .A2(n644), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U642 ( .A(KEYINPUT15), .B(n580), .Z(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT72), .B(n581), .Z(n842) );
  NOR2_X1 U644 ( .A1(n842), .A2(G868), .ZN(n583) );
  INV_X1 U645 ( .A(G868), .ZN(n663) );
  NOR2_X1 U646 ( .A1(n663), .A2(G301), .ZN(n582) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(G284) );
  NAND2_X1 U648 ( .A1(G78), .A2(n644), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G65), .A2(n649), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G91), .A2(n643), .ZN(n586) );
  XNOR2_X1 U652 ( .A(KEYINPUT71), .B(n586), .ZN(n587) );
  NOR2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n648), .A2(G53), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(G299) );
  NOR2_X1 U656 ( .A1(G286), .A2(n663), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n591), .B(KEYINPUT74), .ZN(n593) );
  NOR2_X1 U658 ( .A1(G299), .A2(G868), .ZN(n592) );
  NOR2_X1 U659 ( .A1(n593), .A2(n592), .ZN(G297) );
  NAND2_X1 U660 ( .A1(n594), .A2(G559), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n595), .A2(n984), .ZN(n596) );
  XNOR2_X1 U662 ( .A(n596), .B(KEYINPUT75), .ZN(n597) );
  XOR2_X1 U663 ( .A(KEYINPUT16), .B(n597), .Z(G148) );
  NOR2_X1 U664 ( .A1(G868), .A2(n992), .ZN(n600) );
  NAND2_X1 U665 ( .A1(n984), .A2(G868), .ZN(n598) );
  NOR2_X1 U666 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U667 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U668 ( .A1(G123), .A2(n884), .ZN(n601) );
  XNOR2_X1 U669 ( .A(n601), .B(KEYINPUT18), .ZN(n602) );
  XNOR2_X1 U670 ( .A(n602), .B(KEYINPUT76), .ZN(n604) );
  NAND2_X1 U671 ( .A1(G111), .A2(n882), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U673 ( .A1(G135), .A2(n879), .ZN(n606) );
  NAND2_X1 U674 ( .A1(G99), .A2(n527), .ZN(n605) );
  NAND2_X1 U675 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n931) );
  XNOR2_X1 U677 ( .A(G2096), .B(n931), .ZN(n609) );
  INV_X1 U678 ( .A(G2100), .ZN(n914) );
  NAND2_X1 U679 ( .A1(n609), .A2(n914), .ZN(G156) );
  NAND2_X1 U680 ( .A1(G559), .A2(n984), .ZN(n661) );
  XNOR2_X1 U681 ( .A(n992), .B(n661), .ZN(n610) );
  NOR2_X1 U682 ( .A1(n610), .A2(G860), .ZN(n617) );
  NAND2_X1 U683 ( .A1(n643), .A2(G93), .ZN(n612) );
  NAND2_X1 U684 ( .A1(G67), .A2(n649), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U686 ( .A1(n648), .A2(G55), .ZN(n614) );
  NAND2_X1 U687 ( .A1(G80), .A2(n644), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n615) );
  OR2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n664) );
  XOR2_X1 U690 ( .A(n617), .B(n664), .Z(G145) );
  NAND2_X1 U691 ( .A1(G49), .A2(n648), .ZN(n620) );
  NAND2_X1 U692 ( .A1(G87), .A2(n618), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U694 ( .A1(n649), .A2(n621), .ZN(n624) );
  NAND2_X1 U695 ( .A1(G74), .A2(G651), .ZN(n622) );
  XOR2_X1 U696 ( .A(KEYINPUT77), .B(n622), .Z(n623) );
  NAND2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U698 ( .A(KEYINPUT78), .B(n625), .ZN(G288) );
  NAND2_X1 U699 ( .A1(G61), .A2(n649), .ZN(n626) );
  XOR2_X1 U700 ( .A(KEYINPUT79), .B(n626), .Z(n628) );
  NAND2_X1 U701 ( .A1(n643), .A2(G86), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U703 ( .A(KEYINPUT80), .B(n629), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n644), .A2(G73), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n630), .B(KEYINPUT2), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n631), .B(KEYINPUT81), .ZN(n632) );
  NOR2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n648), .A2(G48), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U710 ( .A1(n643), .A2(G88), .ZN(n637) );
  NAND2_X1 U711 ( .A1(G62), .A2(n649), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n648), .A2(G50), .ZN(n638) );
  XOR2_X1 U714 ( .A(KEYINPUT82), .B(n638), .Z(n639) );
  NOR2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U716 ( .A1(G75), .A2(n644), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(n641), .ZN(G303) );
  INV_X1 U718 ( .A(G303), .ZN(G166) );
  NAND2_X1 U719 ( .A1(n643), .A2(G85), .ZN(n646) );
  NAND2_X1 U720 ( .A1(G72), .A2(n644), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U722 ( .A(KEYINPUT69), .B(n647), .ZN(n654) );
  NAND2_X1 U723 ( .A1(n648), .A2(G47), .ZN(n651) );
  NAND2_X1 U724 ( .A1(G60), .A2(n649), .ZN(n650) );
  NAND2_X1 U725 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U726 ( .A(KEYINPUT70), .B(n652), .Z(n653) );
  NAND2_X1 U727 ( .A1(n654), .A2(n653), .ZN(G290) );
  XNOR2_X1 U728 ( .A(G288), .B(KEYINPUT19), .ZN(n655) );
  XOR2_X1 U729 ( .A(n655), .B(n664), .Z(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(G305), .ZN(n659) );
  XOR2_X1 U731 ( .A(G299), .B(G166), .Z(n657) );
  XNOR2_X1 U732 ( .A(n657), .B(G290), .ZN(n658) );
  XNOR2_X1 U733 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n660), .B(n992), .ZN(n844) );
  XNOR2_X1 U735 ( .A(n844), .B(n661), .ZN(n662) );
  NOR2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n666) );
  NOR2_X1 U737 ( .A1(G868), .A2(n664), .ZN(n665) );
  NOR2_X1 U738 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2084), .A2(G2078), .ZN(n667) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U745 ( .A1(G220), .A2(G219), .ZN(n671) );
  XNOR2_X1 U746 ( .A(KEYINPUT22), .B(n671), .ZN(n672) );
  NAND2_X1 U747 ( .A1(n672), .A2(G96), .ZN(n673) );
  NOR2_X1 U748 ( .A1(n673), .A2(G218), .ZN(n674) );
  XNOR2_X1 U749 ( .A(n674), .B(KEYINPUT83), .ZN(n893) );
  NAND2_X1 U750 ( .A1(n893), .A2(G2106), .ZN(n678) );
  NAND2_X1 U751 ( .A1(G69), .A2(G120), .ZN(n675) );
  NOR2_X1 U752 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U753 ( .A1(G108), .A2(n676), .ZN(n894) );
  NAND2_X1 U754 ( .A1(n894), .A2(G567), .ZN(n677) );
  NAND2_X1 U755 ( .A1(n678), .A2(n677), .ZN(n895) );
  NAND2_X1 U756 ( .A1(G661), .A2(G483), .ZN(n679) );
  NOR2_X1 U757 ( .A1(n895), .A2(n679), .ZN(n841) );
  NAND2_X1 U758 ( .A1(n841), .A2(G36), .ZN(G176) );
  INV_X1 U759 ( .A(G301), .ZN(G171) );
  NOR2_X1 U760 ( .A1(G164), .A2(G1384), .ZN(n761) );
  NAND2_X1 U761 ( .A1(G160), .A2(G40), .ZN(n760) );
  XOR2_X1 U762 ( .A(KEYINPUT88), .B(n760), .Z(n680) );
  AND2_X1 U763 ( .A1(n727), .A2(G1341), .ZN(n681) );
  AND2_X1 U764 ( .A1(n690), .A2(n984), .ZN(n684) );
  INV_X1 U765 ( .A(G1996), .ZN(n900) );
  NOR2_X1 U766 ( .A1(n727), .A2(n900), .ZN(n683) );
  INV_X1 U767 ( .A(KEYINPUT26), .ZN(n682) );
  XNOR2_X1 U768 ( .A(n683), .B(n682), .ZN(n691) );
  NAND2_X1 U769 ( .A1(n684), .A2(n691), .ZN(n688) );
  INV_X1 U770 ( .A(n727), .ZN(n715) );
  BUF_X1 U771 ( .A(n715), .Z(n729) );
  NOR2_X1 U772 ( .A1(n729), .A2(G1348), .ZN(n686) );
  NOR2_X1 U773 ( .A1(G2067), .A2(n727), .ZN(n685) );
  NOR2_X1 U774 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U775 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U776 ( .A(n689), .B(KEYINPUT94), .ZN(n694) );
  AND2_X1 U777 ( .A1(n691), .A2(n690), .ZN(n692) );
  OR2_X1 U778 ( .A1(n984), .A2(n692), .ZN(n693) );
  NAND2_X1 U779 ( .A1(n694), .A2(n693), .ZN(n700) );
  INV_X1 U780 ( .A(G299), .ZN(n702) );
  XOR2_X1 U781 ( .A(KEYINPUT91), .B(KEYINPUT27), .Z(n696) );
  NAND2_X1 U782 ( .A1(n715), .A2(G2072), .ZN(n695) );
  XNOR2_X1 U783 ( .A(n696), .B(n695), .ZN(n698) );
  XOR2_X1 U784 ( .A(G1956), .B(KEYINPUT92), .Z(n1004) );
  NOR2_X1 U785 ( .A1(n729), .A2(n1004), .ZN(n697) );
  NOR2_X1 U786 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U787 ( .A1(n702), .A2(n701), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n700), .A2(n699), .ZN(n706) );
  NOR2_X1 U789 ( .A1(n702), .A2(n701), .ZN(n704) );
  XNOR2_X1 U790 ( .A(KEYINPUT28), .B(KEYINPUT93), .ZN(n703) );
  XNOR2_X1 U791 ( .A(n704), .B(n703), .ZN(n705) );
  NAND2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U793 ( .A(n707), .B(KEYINPUT29), .ZN(n712) );
  XNOR2_X1 U794 ( .A(G2078), .B(KEYINPUT90), .ZN(n708) );
  XNOR2_X1 U795 ( .A(n708), .B(KEYINPUT25), .ZN(n959) );
  NOR2_X1 U796 ( .A1(n959), .A2(n727), .ZN(n710) );
  AND2_X1 U797 ( .A1(n727), .A2(G1961), .ZN(n709) );
  NOR2_X1 U798 ( .A1(n710), .A2(n709), .ZN(n714) );
  AND2_X1 U799 ( .A1(G171), .A2(n714), .ZN(n711) );
  NOR2_X2 U800 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U801 ( .A(KEYINPUT95), .B(n713), .ZN(n726) );
  NOR2_X1 U802 ( .A1(G171), .A2(n714), .ZN(n722) );
  NOR2_X1 U803 ( .A1(n715), .A2(G1966), .ZN(n716) );
  NOR2_X1 U804 ( .A1(G2084), .A2(n727), .ZN(n740) );
  NOR2_X1 U805 ( .A1(n716), .A2(n740), .ZN(n717) );
  NAND2_X1 U806 ( .A1(G8), .A2(n717), .ZN(n718) );
  XNOR2_X1 U807 ( .A(n718), .B(KEYINPUT30), .ZN(n719) );
  XNOR2_X1 U808 ( .A(KEYINPUT96), .B(n719), .ZN(n720) );
  NOR2_X1 U809 ( .A1(G168), .A2(n720), .ZN(n721) );
  NOR2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U811 ( .A(n723), .B(KEYINPUT97), .ZN(n724) );
  XNOR2_X1 U812 ( .A(n724), .B(KEYINPUT31), .ZN(n725) );
  NAND2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n742) );
  NAND2_X1 U814 ( .A1(n742), .A2(G286), .ZN(n736) );
  NOR2_X1 U815 ( .A1(G2090), .A2(n727), .ZN(n728) );
  XNOR2_X1 U816 ( .A(n728), .B(KEYINPUT98), .ZN(n732) );
  INV_X1 U817 ( .A(G8), .ZN(n730) );
  OR2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n801) );
  NOR2_X1 U819 ( .A1(n801), .A2(G1971), .ZN(n731) );
  NOR2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U821 ( .A(KEYINPUT99), .B(n733), .Z(n734) );
  NAND2_X1 U822 ( .A1(n734), .A2(G303), .ZN(n735) );
  NAND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U824 ( .A(n737), .B(KEYINPUT100), .ZN(n738) );
  NAND2_X1 U825 ( .A1(n738), .A2(G8), .ZN(n739) );
  XNOR2_X1 U826 ( .A(n739), .B(KEYINPUT32), .ZN(n795) );
  NAND2_X1 U827 ( .A1(G8), .A2(n740), .ZN(n741) );
  XOR2_X1 U828 ( .A(KEYINPUT89), .B(n741), .Z(n746) );
  NOR2_X1 U829 ( .A1(G1966), .A2(n801), .ZN(n744) );
  INV_X1 U830 ( .A(n742), .ZN(n743) );
  NOR2_X1 U831 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U832 ( .A1(n746), .A2(n745), .ZN(n794) );
  NAND2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n980) );
  INV_X1 U834 ( .A(n980), .ZN(n747) );
  OR2_X1 U835 ( .A1(n747), .A2(n801), .ZN(n751) );
  INV_X1 U836 ( .A(n751), .ZN(n748) );
  AND2_X1 U837 ( .A1(n794), .A2(n748), .ZN(n749) );
  NAND2_X1 U838 ( .A1(n795), .A2(n749), .ZN(n753) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n758) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n758), .A2(n750), .ZN(n981) );
  OR2_X1 U842 ( .A1(n751), .A2(n981), .ZN(n752) );
  NAND2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n755) );
  XNOR2_X1 U844 ( .A(n755), .B(n754), .ZN(n757) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n791) );
  NAND2_X1 U846 ( .A1(n758), .A2(KEYINPUT33), .ZN(n759) );
  NOR2_X1 U847 ( .A1(n759), .A2(n801), .ZN(n789) );
  XOR2_X1 U848 ( .A(G1981), .B(G305), .Z(n993) );
  NOR2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U850 ( .A(KEYINPUT85), .B(n762), .Z(n822) );
  NAND2_X1 U851 ( .A1(G141), .A2(n879), .ZN(n764) );
  NAND2_X1 U852 ( .A1(G117), .A2(n882), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n527), .A2(G105), .ZN(n765) );
  XNOR2_X1 U855 ( .A(n765), .B(KEYINPUT38), .ZN(n766) );
  XNOR2_X1 U856 ( .A(n766), .B(KEYINPUT87), .ZN(n767) );
  NOR2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n884), .A2(G129), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n866) );
  AND2_X1 U860 ( .A1(n866), .A2(G1996), .ZN(n938) );
  NAND2_X1 U861 ( .A1(G131), .A2(n879), .ZN(n772) );
  NAND2_X1 U862 ( .A1(G95), .A2(n527), .ZN(n771) );
  NAND2_X1 U863 ( .A1(n772), .A2(n771), .ZN(n776) );
  NAND2_X1 U864 ( .A1(G119), .A2(n884), .ZN(n774) );
  NAND2_X1 U865 ( .A1(G107), .A2(n882), .ZN(n773) );
  NAND2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n775) );
  OR2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n870) );
  AND2_X1 U868 ( .A1(n870), .A2(G1991), .ZN(n932) );
  OR2_X1 U869 ( .A1(n938), .A2(n932), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n822), .A2(n777), .ZN(n811) );
  NAND2_X1 U871 ( .A1(G140), .A2(n879), .ZN(n779) );
  NAND2_X1 U872 ( .A1(G104), .A2(n527), .ZN(n778) );
  NAND2_X1 U873 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U874 ( .A(KEYINPUT34), .B(n780), .ZN(n785) );
  NAND2_X1 U875 ( .A1(G128), .A2(n884), .ZN(n782) );
  NAND2_X1 U876 ( .A1(G116), .A2(n882), .ZN(n781) );
  NAND2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U878 ( .A(n783), .B(KEYINPUT35), .Z(n784) );
  NOR2_X1 U879 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U880 ( .A(KEYINPUT36), .B(n786), .Z(n787) );
  XOR2_X1 U881 ( .A(KEYINPUT86), .B(n787), .Z(n873) );
  XNOR2_X1 U882 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NOR2_X1 U883 ( .A1(n873), .A2(n820), .ZN(n948) );
  NAND2_X1 U884 ( .A1(n822), .A2(n948), .ZN(n819) );
  AND2_X1 U885 ( .A1(n811), .A2(n819), .ZN(n805) );
  NAND2_X1 U886 ( .A1(n993), .A2(n805), .ZN(n788) );
  NOR2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n807) );
  NAND2_X1 U889 ( .A1(G8), .A2(G166), .ZN(n792) );
  NOR2_X1 U890 ( .A1(G2090), .A2(n792), .ZN(n793) );
  XNOR2_X1 U891 ( .A(n793), .B(KEYINPUT101), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U894 ( .A1(n798), .A2(n801), .ZN(n803) );
  NOR2_X1 U895 ( .A1(G1981), .A2(G305), .ZN(n799) );
  XOR2_X1 U896 ( .A(n799), .B(KEYINPUT24), .Z(n800) );
  OR2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U901 ( .A(n808), .B(KEYINPUT102), .ZN(n810) );
  XNOR2_X1 U902 ( .A(G1986), .B(G290), .ZN(n990) );
  NAND2_X1 U903 ( .A1(n822), .A2(n990), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n826) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n866), .ZN(n929) );
  INV_X1 U906 ( .A(n811), .ZN(n814) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n870), .ZN(n934) );
  NOR2_X1 U909 ( .A1(n812), .A2(n934), .ZN(n813) );
  NOR2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U911 ( .A1(n929), .A2(n815), .ZN(n816) );
  XOR2_X1 U912 ( .A(n816), .B(KEYINPUT39), .Z(n817) );
  XNOR2_X1 U913 ( .A(KEYINPUT103), .B(n817), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n873), .A2(n820), .ZN(n946) );
  NAND2_X1 U916 ( .A1(n821), .A2(n946), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U918 ( .A(n824), .B(KEYINPUT104), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U920 ( .A(n827), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U921 ( .A(G1348), .B(G2454), .ZN(n828) );
  XNOR2_X1 U922 ( .A(n828), .B(G2430), .ZN(n829) );
  XNOR2_X1 U923 ( .A(n829), .B(G1341), .ZN(n835) );
  XOR2_X1 U924 ( .A(G2443), .B(G2427), .Z(n831) );
  XNOR2_X1 U925 ( .A(G2438), .B(G2446), .ZN(n830) );
  XNOR2_X1 U926 ( .A(n831), .B(n830), .ZN(n833) );
  XOR2_X1 U927 ( .A(G2451), .B(G2435), .Z(n832) );
  XNOR2_X1 U928 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U929 ( .A(n835), .B(n834), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n836), .A2(G14), .ZN(n923) );
  XNOR2_X1 U931 ( .A(KEYINPUT105), .B(n923), .ZN(G401) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n927), .ZN(G217) );
  NAND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n837) );
  XOR2_X1 U934 ( .A(KEYINPUT106), .B(n837), .Z(n838) );
  NAND2_X1 U935 ( .A1(n838), .A2(G661), .ZN(n839) );
  XOR2_X1 U936 ( .A(KEYINPUT107), .B(n839), .Z(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U938 ( .A1(n841), .A2(n840), .ZN(G188) );
  XOR2_X1 U939 ( .A(G301), .B(n842), .Z(n843) );
  XNOR2_X1 U940 ( .A(n843), .B(G286), .ZN(n845) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(n846) );
  NOR2_X1 U942 ( .A1(G37), .A2(n846), .ZN(G397) );
  NAND2_X1 U943 ( .A1(n882), .A2(G112), .ZN(n848) );
  NAND2_X1 U944 ( .A1(G100), .A2(n527), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U946 ( .A(KEYINPUT112), .B(n849), .ZN(n854) );
  NAND2_X1 U947 ( .A1(G124), .A2(n884), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U949 ( .A1(n879), .A2(G136), .ZN(n851) );
  NAND2_X1 U950 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U951 ( .A1(n854), .A2(n853), .ZN(G162) );
  NAND2_X1 U952 ( .A1(G118), .A2(n882), .ZN(n863) );
  NAND2_X1 U953 ( .A1(n884), .A2(G130), .ZN(n855) );
  XNOR2_X1 U954 ( .A(KEYINPUT113), .B(n855), .ZN(n861) );
  NAND2_X1 U955 ( .A1(G142), .A2(n879), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G106), .A2(n527), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(KEYINPUT114), .B(n858), .Z(n859) );
  XNOR2_X1 U959 ( .A(KEYINPUT45), .B(n859), .ZN(n860) );
  NOR2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n864), .B(n931), .ZN(n865) );
  XOR2_X1 U963 ( .A(n866), .B(n865), .Z(n878) );
  XOR2_X1 U964 ( .A(KEYINPUT119), .B(KEYINPUT46), .Z(n868) );
  XNOR2_X1 U965 ( .A(G162), .B(KEYINPUT118), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U967 ( .A(n869), .B(KEYINPUT48), .Z(n872) );
  XOR2_X1 U968 ( .A(n870), .B(KEYINPUT115), .Z(n871) );
  XNOR2_X1 U969 ( .A(n872), .B(n871), .ZN(n874) );
  XOR2_X1 U970 ( .A(n874), .B(n873), .Z(n876) );
  XNOR2_X1 U971 ( .A(G160), .B(G164), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U973 ( .A(n878), .B(n877), .ZN(n891) );
  NAND2_X1 U974 ( .A1(G139), .A2(n879), .ZN(n881) );
  NAND2_X1 U975 ( .A1(G103), .A2(n527), .ZN(n880) );
  NAND2_X1 U976 ( .A1(n881), .A2(n880), .ZN(n890) );
  NAND2_X1 U977 ( .A1(n882), .A2(G115), .ZN(n883) );
  XNOR2_X1 U978 ( .A(KEYINPUT117), .B(n883), .ZN(n887) );
  NAND2_X1 U979 ( .A1(n884), .A2(G127), .ZN(n885) );
  XOR2_X1 U980 ( .A(KEYINPUT116), .B(n885), .Z(n886) );
  NOR2_X1 U981 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U982 ( .A(n888), .B(KEYINPUT47), .ZN(n889) );
  NOR2_X1 U983 ( .A1(n890), .A2(n889), .ZN(n941) );
  XNOR2_X1 U984 ( .A(n891), .B(n941), .ZN(n892) );
  NOR2_X1 U985 ( .A1(G37), .A2(n892), .ZN(G395) );
  INV_X1 U987 ( .A(G120), .ZN(G236) );
  INV_X1 U988 ( .A(G96), .ZN(G221) );
  INV_X1 U989 ( .A(G69), .ZN(G235) );
  NOR2_X1 U990 ( .A1(n894), .A2(n893), .ZN(G325) );
  INV_X1 U991 ( .A(G325), .ZN(G261) );
  INV_X1 U992 ( .A(n895), .ZN(G319) );
  XOR2_X1 U993 ( .A(G1976), .B(G1971), .Z(n897) );
  XNOR2_X1 U994 ( .A(G1986), .B(G1961), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n908) );
  XOR2_X1 U996 ( .A(KEYINPUT109), .B(G2474), .Z(n899) );
  XNOR2_X1 U997 ( .A(G1991), .B(KEYINPUT111), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n904) );
  XNOR2_X1 U999 ( .A(G1981), .B(n900), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(G1966), .B(G1956), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1002 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1003 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1005 ( .A(n908), .B(n907), .Z(G229) );
  XOR2_X1 U1006 ( .A(G2096), .B(KEYINPUT43), .Z(n910) );
  XNOR2_X1 U1007 ( .A(G2090), .B(G2678), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(n911), .B(KEYINPUT42), .Z(n913) );
  XNOR2_X1 U1010 ( .A(G2072), .B(G2067), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n918) );
  XNOR2_X1 U1012 ( .A(KEYINPUT108), .B(n914), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(G2084), .B(G2078), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(n918), .B(n917), .ZN(G227) );
  NOR2_X1 U1016 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(KEYINPUT120), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(n920), .B(n919), .ZN(n925) );
  NOR2_X1 U1019 ( .A1(G397), .A2(G395), .ZN(n921) );
  XOR2_X1 U1020 ( .A(KEYINPUT121), .B(n921), .Z(n922) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(G319), .A2(n926), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  INV_X1 U1026 ( .A(n927), .ZN(G223) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1029 ( .A(KEYINPUT51), .B(n930), .Z(n940) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n936) );
  XOR2_X1 U1031 ( .A(G2084), .B(G160), .Z(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n952) );
  XOR2_X1 U1036 ( .A(G2072), .B(n941), .Z(n943) );
  XOR2_X1 U1037 ( .A(G164), .B(G2078), .Z(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(KEYINPUT50), .B(n944), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(n945), .B(KEYINPUT122), .ZN(n950) );
  INV_X1 U1041 ( .A(n946), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(KEYINPUT52), .B(n953), .ZN(n954) );
  INV_X1 U1046 ( .A(KEYINPUT55), .ZN(n973) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n973), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n955), .A2(G29), .ZN(n1032) );
  XOR2_X1 U1049 ( .A(G29), .B(KEYINPUT124), .Z(n976) );
  XOR2_X1 U1050 ( .A(G32), .B(G1996), .Z(n956) );
  NAND2_X1 U1051 ( .A1(n956), .A2(G28), .ZN(n965) );
  XNOR2_X1 U1052 ( .A(G2072), .B(G33), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G25), .B(G1991), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n963) );
  XOR2_X1 U1055 ( .A(n959), .B(G27), .Z(n961) );
  XNOR2_X1 U1056 ( .A(G2067), .B(G26), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1060 ( .A(KEYINPUT53), .B(n966), .Z(n970) );
  XNOR2_X1 U1061 ( .A(KEYINPUT54), .B(G34), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n967), .B(KEYINPUT123), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(G2084), .B(n968), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(G35), .B(G2090), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n974) );
  XOR2_X1 U1067 ( .A(n974), .B(n973), .Z(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(G11), .A2(n977), .ZN(n1030) );
  INV_X1 U1070 ( .A(G16), .ZN(n1026) );
  XOR2_X1 U1071 ( .A(n1026), .B(KEYINPUT56), .Z(n1002) );
  XOR2_X1 U1072 ( .A(G299), .B(G1956), .Z(n979) );
  NAND2_X1 U1073 ( .A1(G1971), .A2(G303), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n988) );
  XOR2_X1 U1077 ( .A(G171), .B(G1961), .Z(n986) );
  XOR2_X1 U1078 ( .A(n984), .B(G1348), .Z(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(KEYINPUT126), .B(n991), .ZN(n1000) );
  XNOR2_X1 U1083 ( .A(n992), .B(G1341), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G168), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(n995), .B(KEYINPUT57), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(KEYINPUT125), .B(n996), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1028) );
  XNOR2_X1 U1091 ( .A(KEYINPUT127), .B(G1961), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1003), .B(G5), .ZN(n1016) );
  XNOR2_X1 U1093 ( .A(n1004), .B(G20), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(G1341), .B(G19), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(G1981), .B(G6), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(KEYINPUT59), .B(G1348), .Z(n1009) );
  XNOR2_X1 U1099 ( .A(G4), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1101 ( .A(KEYINPUT60), .B(n1012), .Z(n1014) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G21), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1023) );
  XNOR2_X1 U1105 ( .A(G1986), .B(G24), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(G1971), .B(G22), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XOR2_X1 U1108 ( .A(G1976), .B(G23), .Z(n1019) );
  NAND2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1110 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1033), .ZN(G150) );
  INV_X1 U1118 ( .A(G150), .ZN(G311) );
endmodule

