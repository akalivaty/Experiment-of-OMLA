//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G120gat), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT1), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G127gat), .B(G134gat), .ZN(new_n206));
  XOR2_X1   g005(.A(KEYINPUT70), .B(G113gat), .Z(new_n207));
  OAI211_X1 g006(.A(new_n205), .B(new_n206), .C1(new_n207), .C2(new_n204), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n205), .B1(new_n203), .B2(new_n204), .ZN(new_n209));
  INV_X1    g008(.A(new_n206), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n215), .A2(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT23), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT23), .ZN(new_n221));
  AND2_X1   g020(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n213), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n214), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(new_n217), .B2(KEYINPUT23), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n226), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n223), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n215), .A2(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(KEYINPUT67), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(KEYINPUT24), .ZN(new_n238));
  NAND2_X1  g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n238), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n236), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(KEYINPUT24), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT24), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(G183gat), .A3(G190gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n246), .B(KEYINPUT64), .C1(G183gat), .C2(G190gat), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n225), .A2(new_n235), .A3(new_n242), .A4(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(KEYINPUT68), .B(G183gat), .Z(new_n251));
  OAI21_X1  g050(.A(new_n246), .B1(new_n251), .B2(G190gat), .ZN(new_n252));
  INV_X1    g051(.A(G169gat), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n249), .B1(new_n232), .B2(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n252), .A2(new_n230), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT28), .ZN(new_n258));
  NOR2_X1   g057(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(new_n251), .B2(KEYINPUT27), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n260), .B2(G190gat), .ZN(new_n261));
  XOR2_X1   g060(.A(KEYINPUT27), .B(G183gat), .Z(new_n262));
  OR3_X1    g061(.A1(new_n262), .A2(new_n258), .A3(G190gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n265));
  OR3_X1    g064(.A1(new_n265), .A2(new_n214), .A3(KEYINPUT69), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n226), .A2(KEYINPUT26), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT69), .B1(new_n265), .B2(new_n214), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(new_n239), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n212), .B1(new_n257), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n255), .B1(new_n248), .B2(new_n249), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n239), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n273), .B1(new_n261), .B2(new_n263), .ZN(new_n274));
  INV_X1    g073(.A(new_n212), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G227gat), .ZN(new_n277));
  INV_X1    g076(.A(G233gat), .ZN(new_n278));
  OAI22_X1  g077(.A1(new_n271), .A2(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(KEYINPUT74), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n277), .A2(new_n278), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n257), .A2(new_n270), .A3(new_n212), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n275), .B1(new_n272), .B2(new_n274), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n280), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n282), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT34), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n281), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT32), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n284), .A2(new_n283), .A3(new_n285), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT71), .A4(new_n283), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G15gat), .B(G43gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G71gat), .B(G99gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n301), .A2(KEYINPUT72), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(KEYINPUT72), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(KEYINPUT33), .A3(new_n303), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n291), .A2(KEYINPUT75), .B1(new_n297), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n281), .A2(new_n288), .A3(new_n306), .A4(new_n290), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n295), .A2(new_n296), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT33), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(KEYINPUT32), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n311), .A3(new_n301), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n305), .A2(new_n307), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n307), .B1(new_n305), .B2(new_n312), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n202), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n305), .A2(new_n312), .ZN(new_n316));
  INV_X1    g115(.A(new_n307), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n305), .A2(new_n307), .A3(new_n312), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(KEYINPUT36), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G197gat), .B(G204gat), .ZN(new_n321));
  INV_X1    g120(.A(G211gat), .ZN(new_n322));
  INV_X1    g121(.A(G218gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(KEYINPUT22), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G211gat), .B(G218gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G141gat), .B(G148gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n329), .B1(KEYINPUT2), .B2(new_n330), .ZN(new_n331));
  OR2_X1    g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n330), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n330), .B(new_n332), .C1(new_n329), .C2(KEYINPUT2), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT79), .B1(new_n336), .B2(KEYINPUT3), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT79), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n334), .A2(new_n338), .A3(new_n339), .A4(new_n335), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n328), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G228gat), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n343), .A2(new_n344), .A3(new_n278), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n327), .A2(KEYINPUT29), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n346), .A2(KEYINPUT85), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n339), .B1(new_n346), .B2(KEYINPUT85), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n336), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n328), .A2(new_n342), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT3), .B1(new_n352), .B2(KEYINPUT84), .ZN(new_n353));
  OR3_X1    g152(.A1(new_n327), .A2(KEYINPUT84), .A3(KEYINPUT29), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI22_X1  g154(.A1(new_n355), .A2(new_n343), .B1(new_n344), .B2(new_n278), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT86), .B(G22gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n350), .A2(new_n356), .A3(new_n358), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363));
  INV_X1    g162(.A(G50gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n367), .B(KEYINPUT83), .Z(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n362), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n361), .A2(new_n367), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n357), .A2(G22gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT5), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n351), .A2(KEYINPUT80), .A3(new_n275), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(new_n336), .B2(new_n212), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n376), .B(new_n378), .C1(new_n351), .C2(new_n275), .ZN(new_n379));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n375), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n275), .B1(KEYINPUT3), .B2(new_n336), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n341), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n376), .A2(new_n385), .A3(new_n378), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n351), .A2(KEYINPUT4), .A3(new_n275), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n384), .A2(new_n380), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  XOR2_X1   g188(.A(G1gat), .B(G29gat), .Z(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G57gat), .B(G85gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n381), .B1(new_n341), .B2(new_n383), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n378), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n385), .B1(new_n336), .B2(new_n212), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n395), .A2(new_n397), .A3(new_n375), .A4(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n389), .A2(new_n394), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT6), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n394), .B1(new_n389), .B2(new_n399), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI211_X1 g203(.A(new_n401), .B(new_n394), .C1(new_n389), .C2(new_n399), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(G226gat), .A2(G233gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n408), .B1(new_n272), .B2(new_n274), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT78), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n411), .B(new_n408), .C1(new_n272), .C2(new_n274), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n342), .B1(new_n272), .B2(new_n274), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n407), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(KEYINPUT77), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT77), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n414), .B2(new_n407), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n413), .B(new_n328), .C1(new_n416), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n409), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT76), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n327), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n407), .B1(new_n257), .B2(new_n270), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(new_n407), .B2(new_n414), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT76), .B1(new_n424), .B2(new_n328), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n419), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n421), .B1(new_n420), .B2(new_n327), .ZN(new_n432));
  AOI211_X1 g231(.A(KEYINPUT76), .B(new_n328), .C1(new_n415), .C2(new_n409), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(new_n419), .A3(new_n429), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n435), .A3(KEYINPUT30), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT30), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n434), .A2(new_n437), .A3(new_n419), .A4(new_n429), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n406), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n315), .B(new_n320), .C1(new_n374), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n406), .A2(new_n435), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT37), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n419), .A2(new_n442), .A3(new_n422), .A4(new_n425), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n434), .A2(KEYINPUT87), .A3(new_n442), .A4(new_n419), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n429), .B1(new_n426), .B2(KEYINPUT37), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n441), .B1(new_n449), .B2(KEYINPUT38), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n442), .B1(new_n420), .B2(new_n328), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n413), .B1(new_n418), .B2(new_n416), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(new_n328), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n429), .A2(KEYINPUT38), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT88), .B1(new_n447), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n447), .A2(new_n455), .A3(KEYINPUT88), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n450), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n397), .A2(new_n384), .A3(new_n398), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n381), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n461), .A2(KEYINPUT39), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n379), .A2(new_n381), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(KEYINPUT39), .A3(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n462), .A2(KEYINPUT40), .A3(new_n394), .A4(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n403), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT40), .ZN(new_n468));
  INV_X1    g267(.A(new_n464), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n394), .B1(new_n461), .B2(KEYINPUT39), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n436), .A2(new_n467), .A3(new_n438), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n374), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n440), .B1(new_n459), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT35), .ZN(new_n477));
  INV_X1    g276(.A(new_n439), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n374), .B1(new_n313), .B2(new_n314), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n362), .A2(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(new_n318), .B2(new_n319), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n476), .A2(new_n477), .ZN(new_n483));
  NAND2_X1  g282(.A1(KEYINPUT89), .A2(KEYINPUT35), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n482), .A2(new_n439), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n475), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G113gat), .B(G141gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(G197gat), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT11), .B(G169gat), .Z(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT12), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G43gat), .B(G50gat), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n494), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n496));
  INV_X1    g295(.A(G36gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G43gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(KEYINPUT91), .A3(G50gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT15), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n495), .B(new_n500), .C1(new_n502), .C2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n499), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT90), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(new_n498), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n496), .A2(KEYINPUT90), .A3(new_n497), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n510), .A2(new_n511), .B1(G29gat), .B2(G36gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n494), .A2(KEYINPUT15), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT16), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(G1gat), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n515), .A2(G1gat), .ZN(new_n519));
  OAI21_X1  g318(.A(G8gat), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G8gat), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n517), .B(new_n521), .C1(G1gat), .C2(new_n515), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n514), .B(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n525), .B(KEYINPUT13), .Z(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n520), .A2(new_n522), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n529));
  NAND2_X1  g328(.A1(G29gat), .A2(G36gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n530), .A3(new_n500), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n506), .B1(new_n501), .B2(new_n494), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n498), .A2(new_n509), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(new_n511), .A3(new_n499), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n513), .B1(new_n535), .B2(new_n530), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n529), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n507), .B(KEYINPUT17), .C1(new_n512), .C2(new_n513), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n528), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT93), .B1(new_n514), .B2(new_n523), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n528), .A2(new_n537), .A3(new_n538), .A4(KEYINPUT93), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n541), .A2(new_n542), .B1(G229gat), .B2(G233gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n527), .B1(new_n543), .B2(KEYINPUT18), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n542), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n545), .A2(KEYINPUT18), .A3(new_n525), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n493), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n525), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT18), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n543), .A2(KEYINPUT18), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n550), .A2(new_n492), .A3(new_n551), .A4(new_n527), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n547), .A2(new_n552), .A3(KEYINPUT94), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT94), .B1(new_n547), .B2(new_n552), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n487), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n557));
  INV_X1    g356(.A(G85gat), .ZN(new_n558));
  INV_X1    g357(.A(G92gat), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G99gat), .A2(G106gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n559), .ZN(new_n563));
  NAND4_X1  g362(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n560), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G99gat), .B(G106gat), .Z(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n537), .B(new_n538), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G190gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n568), .A2(new_n567), .ZN(new_n571));
  AND2_X1   g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n514), .A2(new_n571), .B1(KEYINPUT41), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n569), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n570), .B1(new_n569), .B2(new_n573), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n323), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n569), .A2(new_n573), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(G190gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(G218gat), .A3(new_n574), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT97), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n577), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G134gat), .B(G162gat), .Z(new_n585));
  INV_X1    g384(.A(new_n583), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n577), .A2(new_n580), .A3(new_n581), .A4(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n585), .B1(new_n584), .B2(new_n587), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(G57gat), .A2(G64gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT9), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G57gat), .A2(G64gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(KEYINPUT95), .A3(new_n596), .ZN(new_n598));
  AND2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n597), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(G57gat), .A2(G64gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(new_n591), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n599), .A2(new_n600), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n595), .B(new_n604), .C1(new_n605), .C2(KEYINPUT95), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G127gat), .B(G155gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT20), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n610), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G183gat), .B(G211gat), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n523), .B1(KEYINPUT21), .B2(new_n607), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n615), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n590), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n606), .B(new_n602), .C1(new_n568), .C2(new_n567), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n565), .A2(new_n566), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n565), .A2(new_n566), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n607), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n628), .A2(KEYINPUT99), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n623), .A2(new_n626), .A3(new_n630), .A4(new_n627), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n571), .A2(KEYINPUT10), .A3(new_n607), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n622), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n623), .A2(new_n626), .ZN(new_n635));
  INV_X1    g434(.A(new_n622), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n634), .A2(new_n637), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n621), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n556), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n406), .B(KEYINPUT100), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT101), .B(G1gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1324gat));
  INV_X1    g451(.A(new_n647), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n436), .A2(new_n438), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n521), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT16), .B(G8gat), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n647), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT42), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(KEYINPUT42), .B2(new_n658), .ZN(G1325gat));
  NAND2_X1  g459(.A1(new_n315), .A2(new_n320), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(G15gat), .B1(new_n647), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n318), .A2(new_n319), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(G15gat), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n663), .B1(new_n647), .B2(new_n666), .ZN(G1326gat));
  NOR2_X1   g466(.A1(new_n647), .A2(new_n374), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT43), .B(G22gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  INV_X1    g469(.A(new_n645), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n619), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n590), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n649), .A2(G29gat), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n556), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(KEYINPUT102), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(KEYINPUT45), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n590), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(new_n475), .B2(new_n486), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g481(.A(KEYINPUT44), .B(new_n679), .C1(new_n475), .C2(new_n486), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n547), .A2(new_n552), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n672), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G29gat), .B1(new_n688), .B2(new_n649), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n678), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT45), .B1(new_n676), .B2(new_n677), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n690), .A2(new_n691), .ZN(G1328gat));
  NAND2_X1  g491(.A1(new_n556), .A2(new_n673), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n693), .A2(G36gat), .A3(new_n654), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT46), .ZN(new_n695));
  OAI21_X1  g494(.A(G36gat), .B1(new_n688), .B2(new_n654), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(G1329gat));
  NAND3_X1  g496(.A1(new_n684), .A2(new_n661), .A3(new_n687), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G43gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n665), .A2(G43gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n556), .A2(new_n673), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT103), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n556), .A2(new_n704), .A3(new_n673), .A4(new_n701), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n700), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n699), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n699), .B2(new_n706), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(G1330gat));
  OAI21_X1  g509(.A(new_n364), .B1(new_n693), .B2(new_n374), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n481), .A2(G50gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n688), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g513(.A(new_n458), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n456), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n473), .B1(new_n716), .B2(new_n450), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n480), .B(new_n485), .C1(new_n717), .C2(new_n440), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n621), .A2(new_n685), .A3(new_n671), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n648), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT105), .B(G57gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1332gat));
  AOI21_X1  g522(.A(new_n654), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT106), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n726), .B(new_n727), .Z(G1333gat));
  INV_X1    g527(.A(new_n720), .ZN(new_n729));
  OAI21_X1  g528(.A(G71gat), .B1(new_n729), .B2(new_n662), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n665), .A2(G71gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n720), .A2(new_n481), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g535(.A1(new_n620), .A2(new_n685), .A3(new_n671), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n682), .A2(new_n648), .A3(new_n683), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G85gat), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n620), .A2(new_n685), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n679), .B(new_n740), .C1(new_n475), .C2(new_n486), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n718), .A2(KEYINPUT51), .A3(new_n679), .A4(new_n740), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n743), .A2(new_n744), .A3(KEYINPUT108), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n741), .A2(new_n746), .A3(new_n742), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n648), .A2(new_n558), .A3(new_n645), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n739), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1336gat));
  NOR3_X1   g551(.A1(new_n654), .A2(G92gat), .A3(new_n671), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT110), .B1(new_n748), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n682), .A2(new_n655), .A3(new_n683), .A4(new_n737), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G92gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n748), .A2(KEYINPUT110), .A3(new_n754), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n744), .ZN(new_n761));
  AOI22_X1  g560(.A1(G92gat), .A2(new_n757), .B1(new_n761), .B2(new_n753), .ZN(new_n762));
  OAI22_X1  g561(.A1(new_n759), .A2(new_n760), .B1(new_n756), .B2(new_n762), .ZN(G1337gat));
  NAND3_X1  g562(.A1(new_n684), .A2(new_n661), .A3(new_n737), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G99gat), .ZN(new_n765));
  OR3_X1    g564(.A1(new_n665), .A2(G99gat), .A3(new_n671), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n748), .B2(new_n766), .ZN(G1338gat));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n682), .A2(new_n481), .A3(new_n683), .A4(new_n737), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT53), .B1(new_n769), .B2(G106gat), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n374), .A2(G106gat), .A3(new_n671), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n745), .A2(new_n747), .A3(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(G106gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n761), .A2(new_n771), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n768), .B1(new_n773), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n770), .A2(new_n772), .ZN(new_n779));
  AOI22_X1  g578(.A1(G106gat), .A2(new_n769), .B1(new_n761), .B2(new_n771), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n779), .B(KEYINPUT111), .C1(new_n774), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n781), .ZN(G1339gat));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n628), .A2(KEYINPUT99), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n784), .A2(new_n636), .A3(new_n632), .A4(new_n631), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n634), .A2(KEYINPUT54), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n787), .B(new_n622), .C1(new_n629), .C2(new_n633), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n642), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n783), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT113), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n634), .A2(KEYINPUT54), .A3(new_n785), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n792), .A2(KEYINPUT55), .A3(new_n642), .A4(new_n788), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n789), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(new_n792), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(new_n644), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT114), .B1(new_n791), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n790), .B(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n798), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n799), .A2(new_n685), .A3(new_n804), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n545), .A2(new_n525), .B1(new_n524), .B2(new_n526), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n491), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n552), .A2(new_n645), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n679), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n552), .A2(new_n807), .ZN(new_n810));
  AND4_X1   g609(.A1(new_n679), .A2(new_n799), .A3(new_n810), .A4(new_n804), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n619), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n646), .A2(new_n686), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n481), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n649), .A2(new_n655), .A3(new_n665), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(G113gat), .B1(new_n817), .B2(new_n555), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n649), .B1(new_n812), .B2(new_n813), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n820), .A2(new_n655), .A3(new_n479), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n685), .A3(new_n207), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n822), .ZN(G1340gat));
  AOI21_X1  g622(.A(G120gat), .B1(new_n821), .B2(new_n645), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n671), .A2(new_n204), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n816), .B2(new_n825), .ZN(G1341gat));
  AND2_X1   g625(.A1(new_n821), .A2(new_n620), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(G127gat), .B1(new_n827), .B2(new_n828), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n620), .A2(G127gat), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n829), .A2(new_n830), .B1(new_n816), .B2(new_n831), .ZN(G1342gat));
  NAND2_X1  g631(.A1(new_n679), .A2(new_n654), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT116), .ZN(new_n834));
  NOR4_X1   g633(.A1(new_n820), .A2(G134gat), .A3(new_n479), .A4(new_n834), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT56), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n816), .A2(new_n679), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n837), .A2(KEYINPUT117), .A3(G134gat), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT117), .B1(new_n837), .B2(G134gat), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(G1343gat));
  NOR2_X1   g639(.A1(new_n649), .A2(new_n655), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n662), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n812), .A2(new_n813), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT57), .B1(new_n844), .B2(new_n481), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n808), .B(KEYINPUT118), .ZN(new_n847));
  XNOR2_X1  g646(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n786), .B2(new_n789), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n795), .A2(new_n797), .A3(new_n644), .A4(new_n849), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n850), .A2(KEYINPUT120), .B1(new_n553), .B2(new_n554), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(KEYINPUT120), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n590), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n619), .B1(new_n854), .B2(new_n811), .ZN(new_n855));
  AOI211_X1 g654(.A(new_n846), .B(new_n374), .C1(new_n855), .C2(new_n813), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n843), .B1(new_n845), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G141gat), .B1(new_n857), .B2(new_n555), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n661), .A2(new_n374), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n819), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n655), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n555), .A2(G141gat), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT58), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n858), .A2(new_n859), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n859), .B1(new_n858), .B2(new_n864), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n685), .B(new_n843), .C1(new_n845), .C2(new_n856), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n868), .A2(G141gat), .B1(new_n862), .B2(new_n863), .ZN(new_n869));
  OAI22_X1  g668(.A1(new_n865), .A2(new_n866), .B1(new_n867), .B2(new_n869), .ZN(G1344gat));
  INV_X1    g669(.A(G148gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n862), .A2(new_n871), .A3(new_n645), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n842), .A2(KEYINPUT123), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n842), .A2(KEYINPUT123), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n645), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n646), .A2(new_n555), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n810), .B1(new_n588), .B2(new_n589), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n801), .A2(new_n802), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n880), .B1(new_n853), .B2(new_n590), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n877), .B1(new_n881), .B2(new_n620), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT124), .B(new_n877), .C1(new_n881), .C2(new_n620), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n481), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n846), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n374), .A2(new_n846), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n844), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n876), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n871), .B1(new_n890), .B2(KEYINPUT125), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892));
  INV_X1    g691(.A(new_n889), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n846), .B2(new_n886), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n892), .B1(new_n894), .B2(new_n876), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n873), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n645), .B(new_n843), .C1(new_n845), .C2(new_n856), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n871), .A2(KEYINPUT59), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n897), .A2(KEYINPUT122), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT122), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n872), .B1(new_n896), .B2(new_n901), .ZN(G1345gat));
  OAI21_X1  g701(.A(G155gat), .B1(new_n857), .B2(new_n619), .ZN(new_n903));
  INV_X1    g702(.A(G155gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n862), .A2(new_n904), .A3(new_n620), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1346gat));
  OAI21_X1  g705(.A(G162gat), .B1(new_n857), .B2(new_n590), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n834), .A2(G162gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n861), .B2(new_n908), .ZN(G1347gat));
  NAND2_X1  g708(.A1(new_n649), .A2(new_n655), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n665), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n814), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(G169gat), .B1(new_n913), .B2(new_n555), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n648), .B1(new_n812), .B2(new_n813), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n479), .A2(new_n654), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n685), .A2(new_n231), .A3(new_n233), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(G1348gat));
  OAI21_X1  g718(.A(G176gat), .B1(new_n913), .B2(new_n671), .ZN(new_n920));
  INV_X1    g719(.A(new_n917), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n220), .A3(new_n645), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1349gat));
  NAND2_X1  g722(.A1(new_n912), .A2(new_n620), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(new_n251), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n917), .A2(new_n262), .A3(new_n619), .ZN(new_n926));
  OR3_X1    g725(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT60), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT60), .B1(new_n925), .B2(new_n926), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1350gat));
  NAND3_X1  g728(.A1(new_n921), .A2(new_n570), .A3(new_n679), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n912), .A2(new_n679), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n932));
  AND4_X1   g731(.A1(KEYINPUT126), .A2(new_n931), .A3(new_n932), .A4(G190gat), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n570), .B1(new_n934), .B2(KEYINPUT61), .ZN(new_n935));
  AOI22_X1  g734(.A1(new_n931), .A2(new_n935), .B1(KEYINPUT126), .B2(new_n932), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n930), .B1(new_n933), .B2(new_n936), .ZN(G1351gat));
  AND3_X1   g736(.A1(new_n915), .A2(new_n655), .A3(new_n860), .ZN(new_n938));
  INV_X1    g737(.A(G197gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n939), .A3(new_n685), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT127), .Z(new_n941));
  NOR2_X1   g740(.A1(new_n910), .A2(new_n661), .ZN(new_n942));
  INV_X1    g741(.A(new_n887), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n893), .ZN(new_n944));
  OAI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n555), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n941), .A2(new_n945), .ZN(G1352gat));
  INV_X1    g745(.A(G204gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n938), .A2(new_n947), .A3(new_n645), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT62), .Z(new_n949));
  OAI21_X1  g748(.A(G204gat), .B1(new_n944), .B2(new_n671), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1353gat));
  NAND3_X1  g750(.A1(new_n938), .A2(new_n322), .A3(new_n620), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n620), .B(new_n942), .C1(new_n943), .C2(new_n893), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n953), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n953), .B2(G211gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(G1354gat));
  OAI21_X1  g755(.A(G218gat), .B1(new_n944), .B2(new_n590), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n938), .A2(new_n323), .A3(new_n679), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1355gat));
endmodule


