//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933;
  NOR2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202));
  AND2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  AOI211_X1 g007(.A(new_n202), .B(new_n203), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n203), .B2(new_n202), .ZN(new_n212));
  INV_X1    g011(.A(G141gat), .ZN(new_n213));
  INV_X1    g012(.A(G148gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(KEYINPUT76), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(new_n217), .A3(new_n204), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT77), .ZN(new_n219));
  XOR2_X1   g018(.A(G155gat), .B(G162gat), .Z(new_n220));
  AND3_X1   g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n219), .B1(new_n218), .B2(new_n220), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n210), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n218), .A2(new_n220), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT77), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(new_n229), .A3(new_n210), .ZN(new_n230));
  INV_X1    g029(.A(G113gat), .ZN(new_n231));
  INV_X1    g030(.A(G120gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g033(.A1(G113gat), .A2(G120gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n237));
  INV_X1    g036(.A(G134gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G127gat), .ZN(new_n239));
  INV_X1    g038(.A(G127gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G134gat), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n237), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT67), .B1(new_n238), .B2(G127gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n236), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n234), .B1(G113gat), .B2(G120gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n235), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(new_n239), .A3(new_n241), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n248), .A3(KEYINPUT78), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT78), .B1(new_n244), .B2(new_n248), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n224), .A2(new_n230), .A3(new_n252), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n244), .A2(new_n248), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n254), .B(new_n210), .C1(new_n221), .C2(new_n222), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT4), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n228), .A2(new_n257), .A3(new_n210), .A4(new_n254), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT5), .ZN(new_n260));
  NAND2_X1  g059(.A1(G225gat), .A2(G233gat), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n253), .A2(new_n259), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n209), .B1(new_n226), .B2(new_n227), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT78), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n249), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT80), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT80), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n252), .A2(new_n223), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n255), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n261), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n260), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT79), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n256), .A2(new_n258), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n255), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n276), .A2(new_n253), .A3(new_n277), .A4(new_n261), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n273), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n274), .B1(new_n273), .B2(new_n278), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n262), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G1gat), .B(G29gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT0), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G57gat), .ZN(new_n284));
  INV_X1    g083(.A(G85gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n286), .B(new_n262), .C1(new_n279), .C2(new_n280), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G8gat), .B(G36gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(G92gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT73), .B(G64gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  NAND2_X1  g094(.A1(G226gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298));
  NOR2_X1   g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(KEYINPUT23), .ZN(new_n300));
  NAND2_X1  g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(KEYINPUT24), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G183gat), .B(G190gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT65), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n300), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n309), .A2(G169gat), .A3(G176gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT64), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G169gat), .ZN(new_n314));
  INV_X1    g113(.A(G176gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT23), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT64), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(new_n311), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n298), .B1(new_n308), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT66), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT26), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n299), .A2(KEYINPUT66), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n311), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G183gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT27), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT27), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G183gat), .ZN(new_n329));
  INV_X1    g128(.A(G190gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT28), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT27), .B(G183gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(new_n330), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n325), .A2(new_n332), .A3(new_n301), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n311), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n298), .B1(new_n299), .B2(KEYINPUT23), .ZN(new_n338));
  OAI22_X1  g137(.A1(new_n337), .A2(new_n338), .B1(new_n307), .B2(new_n298), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n326), .A2(G190gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n330), .A2(G183gat), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n305), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(new_n302), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n297), .B1(new_n320), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G197gat), .B(G204gat), .Z(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT71), .B(G211gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G218gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT70), .B(KEYINPUT22), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G211gat), .B(G218gat), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n352), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n336), .A2(new_n344), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n307), .B1(new_n342), .B2(new_n302), .ZN(new_n357));
  INV_X1    g156(.A(new_n300), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n319), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT25), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT29), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n346), .B(new_n355), .C1(new_n361), .C2(new_n297), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT72), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(new_n320), .B2(new_n345), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n296), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n355), .B1(new_n366), .B2(new_n346), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n369));
  INV_X1    g168(.A(new_n355), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n356), .A2(new_n360), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n297), .B1(new_n371), .B2(new_n364), .ZN(new_n372));
  INV_X1    g171(.A(new_n346), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n369), .B(new_n370), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n295), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n362), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT37), .B1(new_n377), .B2(new_n367), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT38), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n295), .B(KEYINPUT74), .Z(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(KEYINPUT72), .A3(new_n362), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT37), .B1(new_n383), .B2(new_n374), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n376), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n384), .ZN(new_n386));
  INV_X1    g185(.A(new_n295), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n383), .A2(KEYINPUT37), .A3(new_n374), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n385), .B1(new_n389), .B2(KEYINPUT38), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n281), .A2(KEYINPUT6), .A3(new_n287), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n291), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n393));
  NOR2_X1   g192(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n394));
  NAND2_X1  g193(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n253), .A2(new_n259), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT39), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n272), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n286), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n268), .A2(new_n270), .A3(new_n255), .A4(new_n261), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT39), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n261), .B1(new_n253), .B2(new_n259), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n396), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n267), .B1(KEYINPUT3), .B2(new_n223), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n406), .A2(new_n230), .B1(new_n256), .B2(new_n258), .ZN(new_n407));
  OAI211_X1 g206(.A(KEYINPUT39), .B(new_n401), .C1(new_n407), .C2(new_n261), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n408), .A2(new_n286), .A3(new_n395), .A4(new_n399), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n394), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n288), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g210(.A(KEYINPUT30), .B(new_n295), .C1(new_n368), .C2(new_n375), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n383), .A2(new_n374), .A3(new_n380), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n387), .B1(new_n383), .B2(new_n374), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT75), .B1(new_n415), .B2(KEYINPUT30), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT75), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT30), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n376), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n393), .B1(new_n411), .B2(new_n420), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n412), .A2(new_n413), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n417), .B1(new_n376), .B2(new_n418), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n415), .A2(KEYINPUT75), .A3(KEYINPUT30), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n425), .A2(KEYINPUT86), .A3(new_n288), .A4(new_n410), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n355), .B1(new_n230), .B2(new_n364), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n427), .A2(KEYINPUT84), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n353), .A2(new_n429), .A3(new_n354), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n364), .B1(new_n354), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n229), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n432), .A2(new_n223), .B1(G228gat), .B2(G233gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n427), .A2(KEYINPUT84), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n355), .A2(new_n364), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n263), .B1(new_n436), .B2(new_n229), .ZN(new_n437));
  OAI211_X1 g236(.A(G228gat), .B(G233gat), .C1(new_n437), .C2(new_n427), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT31), .B(G50gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n440), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n435), .A2(new_n442), .A3(new_n438), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G78gat), .B(G106gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(G22gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n441), .A2(new_n446), .A3(new_n443), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n392), .A2(new_n421), .A3(new_n426), .A4(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(KEYINPUT87), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT68), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n371), .B(new_n254), .ZN(new_n454));
  NAND2_X1  g253(.A1(G227gat), .A2(G233gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n453), .B1(new_n456), .B2(KEYINPUT34), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(KEYINPUT34), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT34), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n454), .A2(KEYINPUT68), .A3(new_n459), .A4(new_n455), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(G15gat), .B(G43gat), .Z(new_n462));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n454), .A2(new_n455), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n464), .B1(new_n465), .B2(KEYINPUT33), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT32), .B1(new_n454), .B2(new_n455), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n466), .A2(new_n468), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n461), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n466), .A2(new_n468), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n457), .A2(new_n460), .A3(new_n458), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n469), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT69), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT36), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n477), .B(new_n478), .C1(new_n476), .C2(new_n472), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n472), .A2(new_n475), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT36), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n290), .A2(new_n289), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n273), .A2(new_n278), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT81), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n273), .A2(new_n274), .A3(new_n278), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n286), .B1(new_n487), .B2(new_n262), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n391), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n420), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT82), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n291), .A2(new_n391), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(KEYINPUT82), .A3(new_n420), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n448), .A2(new_n449), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n482), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n450), .A2(new_n480), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n493), .A2(new_n499), .A3(new_n495), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n477), .B1(new_n476), .B2(new_n472), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT35), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n502), .A2(new_n503), .A3(new_n450), .ZN(new_n504));
  INV_X1    g303(.A(new_n491), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n452), .A2(new_n498), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT91), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT92), .ZN(new_n510));
  INV_X1    g309(.A(G8gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT16), .ZN(new_n513));
  AOI21_X1  g312(.A(G1gat), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n512), .B(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT88), .ZN(new_n517));
  OR3_X1    g316(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n519), .A2(new_n520), .B1(G29gat), .B2(G36gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n520), .B2(new_n519), .ZN(new_n522));
  XNOR2_X1  g321(.A(G43gat), .B(G50gat), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n524), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n518), .B(KEYINPUT90), .Z(new_n527));
  INV_X1    g326(.A(new_n516), .ZN(new_n528));
  OAI221_X1 g327(.A(new_n526), .B1(KEYINPUT15), .B2(new_n523), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n515), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n525), .A2(new_n529), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n515), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n531), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT18), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n515), .B(new_n530), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n537), .B(KEYINPUT13), .Z(new_n541));
  AOI22_X1  g340(.A1(new_n538), .A2(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n531), .A2(new_n536), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(KEYINPUT18), .A3(new_n537), .ZN(new_n544));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT11), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(new_n314), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G197gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT12), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n542), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n549), .B1(new_n542), .B2(new_n544), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(G85gat), .A3(G92gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT95), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT7), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  XOR2_X1   g357(.A(G99gat), .B(G106gat), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT96), .ZN(new_n560));
  NAND2_X1  g359(.A1(G99gat), .A2(G106gat), .ZN(new_n561));
  INV_X1    g360(.A(G92gat), .ZN(new_n562));
  AOI22_X1  g361(.A1(KEYINPUT8), .A2(new_n561), .B1(new_n285), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n557), .A2(new_n558), .A3(new_n560), .A4(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n559), .A2(KEYINPUT96), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n532), .A2(new_n535), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT97), .ZN(new_n571));
  AND2_X1   g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n568), .A2(new_n533), .B1(KEYINPUT41), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G134gat), .B(G162gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n574), .B(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n578));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n574), .B(new_n575), .ZN(new_n582));
  INV_X1    g381(.A(new_n580), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT21), .ZN(new_n587));
  XOR2_X1   g386(.A(G57gat), .B(G64gat), .Z(new_n588));
  AND2_X1   g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n588), .B1(KEYINPUT9), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n591));
  NOR2_X1   g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n589), .A2(new_n592), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  OAI21_X1  g394(.A(new_n515), .B1(new_n587), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G183gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n598));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n597), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n595), .A2(new_n587), .ZN(new_n602));
  XOR2_X1   g401(.A(G127gat), .B(G155gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G211gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n601), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n595), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n568), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT10), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n566), .A2(new_n595), .A3(new_n567), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT98), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n608), .A2(new_n613), .A3(new_n609), .A4(new_n610), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n568), .A2(KEYINPUT10), .A3(new_n607), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT99), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT99), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n612), .A2(new_n618), .A3(new_n614), .A4(new_n615), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n617), .A2(new_n619), .B1(G230gat), .B2(G233gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n621), .B1(new_n608), .B2(new_n610), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G176gat), .ZN(new_n624));
  INV_X1    g423(.A(G204gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n620), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n616), .A2(new_n621), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n627), .B1(new_n630), .B2(new_n622), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n586), .A2(new_n606), .A3(new_n633), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n507), .A2(new_n552), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n494), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g437(.A(KEYINPUT16), .B(G8gat), .Z(new_n639));
  NAND4_X1  g438(.A1(new_n635), .A2(KEYINPUT42), .A3(new_n425), .A4(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT42), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n635), .A2(new_n425), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n639), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(G8gat), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n647), .A2(KEYINPUT101), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(KEYINPUT101), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n640), .B(new_n646), .C1(new_n648), .C2(new_n649), .ZN(G1325gat));
  INV_X1    g449(.A(G15gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n651), .A3(new_n502), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n635), .A2(new_n482), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n652), .B1(new_n653), .B2(new_n651), .ZN(G1326gat));
  NAND2_X1  g453(.A1(new_n635), .A2(new_n497), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT43), .B(G22gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1327gat));
  NOR2_X1   g456(.A1(new_n507), .A2(new_n586), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n632), .A2(new_n552), .A3(new_n606), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n660), .A2(G29gat), .A3(new_n494), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT45), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n507), .B2(new_n586), .ZN(new_n664));
  INV_X1    g463(.A(new_n495), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT82), .B1(new_n494), .B2(new_n420), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n497), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n482), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n421), .A2(new_n450), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n669), .A2(KEYINPUT87), .A3(new_n392), .A4(new_n426), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT87), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n451), .A2(new_n671), .ZN(new_n672));
  AND4_X1   g471(.A1(new_n667), .A2(new_n668), .A3(new_n670), .A4(new_n672), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n500), .A2(KEYINPUT35), .B1(new_n505), .B2(new_n504), .ZN(new_n674));
  OAI211_X1 g473(.A(KEYINPUT44), .B(new_n585), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n664), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n659), .ZN(new_n677));
  OAI21_X1  g476(.A(G29gat), .B1(new_n677), .B2(new_n494), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT102), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n662), .A2(new_n681), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(G1328gat));
  OR3_X1    g482(.A1(new_n660), .A2(G36gat), .A3(new_n420), .ZN(new_n684));
  AND2_X1   g483(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n685));
  NOR2_X1   g484(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G36gat), .B1(new_n677), .B2(new_n420), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n687), .B(new_n688), .C1(new_n685), .C2(new_n684), .ZN(G1329gat));
  OAI21_X1  g488(.A(G43gat), .B1(new_n677), .B2(new_n668), .ZN(new_n690));
  INV_X1    g489(.A(new_n502), .ZN(new_n691));
  OR3_X1    g490(.A1(new_n660), .A2(G43gat), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n695));
  AOI211_X1 g494(.A(G50gat), .B(new_n450), .C1(new_n660), .C2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n658), .A2(KEYINPUT104), .A3(new_n659), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n676), .A2(new_n497), .A3(new_n659), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n696), .A2(new_n697), .B1(new_n698), .B2(G50gat), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT48), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NOR2_X1   g502(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n699), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n702), .A2(new_n705), .ZN(G1331gat));
  NAND2_X1  g505(.A1(new_n452), .A2(new_n498), .ZN(new_n707));
  INV_X1    g506(.A(new_n674), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n606), .ZN(new_n710));
  INV_X1    g509(.A(new_n552), .ZN(new_n711));
  NOR4_X1   g510(.A1(new_n585), .A2(new_n710), .A3(new_n711), .A4(new_n633), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n636), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g515(.A1(new_n713), .A2(new_n420), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT49), .B(G64gat), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT106), .ZN(G1333gat));
  OR3_X1    g521(.A1(new_n713), .A2(G71gat), .A3(new_n691), .ZN(new_n723));
  OAI21_X1  g522(.A(G71gat), .B1(new_n713), .B2(new_n668), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g525(.A1(new_n714), .A2(new_n497), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g527(.A1(new_n606), .A2(new_n711), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n709), .A2(new_n585), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n658), .A2(KEYINPUT51), .A3(new_n729), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT51), .B1(new_n658), .B2(new_n729), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT108), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n632), .A2(new_n285), .A3(new_n636), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT109), .Z(new_n741));
  AND2_X1   g540(.A1(new_n729), .A2(new_n632), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n664), .A2(new_n675), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n664), .A2(new_n675), .A3(KEYINPUT107), .A4(new_n742), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n636), .A3(new_n746), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n739), .A2(new_n741), .B1(G85gat), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT110), .ZN(G1336gat));
  NAND4_X1  g548(.A1(new_n664), .A2(new_n675), .A3(new_n425), .A4(new_n742), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT52), .B1(new_n750), .B2(G92gat), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n633), .A2(G92gat), .A3(new_n420), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n738), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n732), .B2(new_n733), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n745), .A2(new_n425), .A3(new_n746), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(G92gat), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n754), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT111), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n761), .B(new_n754), .C1(new_n757), .C2(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(G1337gat));
  NAND3_X1  g562(.A1(new_n745), .A2(new_n482), .A3(new_n746), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT112), .B(G99gat), .Z(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR3_X1    g565(.A1(new_n633), .A2(new_n691), .A3(new_n765), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n738), .B2(new_n767), .ZN(G1338gat));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  OAI21_X1  g568(.A(G106gat), .B1(new_n743), .B2(new_n450), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n633), .A2(G106gat), .A3(new_n450), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n769), .B(new_n770), .C1(new_n738), .C2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n745), .A2(new_n497), .A3(new_n746), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(G106gat), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n771), .B(KEYINPUT113), .Z(new_n776));
  INV_X1    g575(.A(new_n733), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(new_n736), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n778), .A2(KEYINPUT114), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(KEYINPUT114), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n775), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n773), .B1(new_n781), .B2(new_n769), .ZN(G1339gat));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n626), .B1(new_n630), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT54), .B1(new_n616), .B2(new_n621), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n620), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n552), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n784), .B(KEYINPUT55), .C1(new_n620), .C2(new_n785), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n629), .B(new_n788), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  OAI22_X1  g592(.A1(new_n543), .A2(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n550), .B1(new_n548), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n632), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n585), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n629), .B1(new_n791), .B2(new_n792), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n786), .A2(new_n787), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n585), .A2(new_n795), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n710), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n634), .A2(new_n711), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n494), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n804), .A2(new_n420), .A3(new_n499), .ZN(new_n805));
  AOI21_X1  g604(.A(G113gat), .B1(new_n805), .B2(new_n711), .ZN(new_n806));
  AND4_X1   g605(.A1(new_n420), .A2(new_n804), .A3(new_n450), .A4(new_n502), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n552), .A2(new_n231), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(G1340gat));
  AOI21_X1  g608(.A(G120gat), .B1(new_n805), .B2(new_n632), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n633), .A2(new_n232), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n807), .B2(new_n811), .ZN(G1341gat));
  NAND3_X1  g611(.A1(new_n805), .A2(new_n240), .A3(new_n606), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n807), .A2(new_n606), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n240), .ZN(G1342gat));
  NAND3_X1  g614(.A1(new_n805), .A2(new_n238), .A3(new_n585), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n816), .A2(KEYINPUT56), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(KEYINPUT56), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n807), .A2(new_n585), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n817), .B(new_n818), .C1(new_n238), .C2(new_n819), .ZN(G1343gat));
  NOR3_X1   g619(.A1(new_n482), .A2(new_n494), .A3(new_n425), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n450), .B1(new_n802), .B2(new_n803), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n797), .A2(KEYINPUT116), .B1(new_n798), .B2(new_n800), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n827));
  AOI211_X1 g626(.A(new_n827), .B(new_n585), .C1(new_n793), .C2(new_n796), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n710), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n450), .B1(new_n829), .B2(new_n803), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n711), .B(new_n825), .C1(new_n830), .C2(new_n824), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(G141gat), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n482), .A2(new_n450), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n804), .A2(new_n420), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n213), .A3(new_n711), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT58), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n832), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(G1344gat));
  NAND3_X1  g639(.A1(new_n834), .A2(new_n214), .A3(new_n632), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842));
  NAND2_X1  g641(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n823), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  AOI211_X1 g646(.A(new_n450), .B(new_n847), .C1(new_n802), .C2(new_n803), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n632), .B(new_n821), .C1(new_n845), .C2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n214), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n823), .B1(new_n846), .B2(new_n844), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n823), .B2(new_n844), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n853), .A2(KEYINPUT118), .A3(new_n632), .A4(new_n821), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n842), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n825), .B1(new_n830), .B2(new_n824), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n633), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n842), .A2(G148gat), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n841), .B1(new_n855), .B2(new_n859), .ZN(G1345gat));
  OAI21_X1  g659(.A(G155gat), .B1(new_n856), .B2(new_n710), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n834), .A2(new_n205), .A3(new_n606), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1346gat));
  OAI21_X1  g662(.A(G162gat), .B1(new_n856), .B2(new_n586), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n834), .A2(new_n206), .A3(new_n585), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1347gat));
  NAND2_X1  g665(.A1(new_n802), .A2(new_n803), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n691), .A2(new_n420), .A3(new_n497), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n494), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(G169gat), .B1(new_n872), .B2(new_n552), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n867), .A2(new_n494), .A3(new_n425), .A4(new_n499), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n874), .A2(new_n875), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n552), .A2(G169gat), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n879), .A2(KEYINPUT120), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT120), .B1(new_n879), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n873), .B1(new_n881), .B2(new_n882), .ZN(G1348gat));
  NOR3_X1   g682(.A1(new_n872), .A2(new_n315), .A3(new_n633), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n877), .A2(new_n878), .A3(new_n633), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT122), .B1(new_n885), .B2(G176gat), .ZN(new_n886));
  INV_X1    g685(.A(new_n878), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n632), .A3(new_n876), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(new_n315), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n884), .B1(new_n886), .B2(new_n890), .ZN(G1349gat));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n869), .B(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n326), .B1(new_n893), .B2(new_n606), .ZN(new_n894));
  INV_X1    g693(.A(new_n874), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n333), .A3(new_n606), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT123), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT60), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G183gat), .B1(new_n872), .B2(new_n710), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n900));
  INV_X1    g699(.A(new_n897), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n898), .A2(new_n902), .ZN(G1350gat));
  NAND3_X1  g702(.A1(new_n879), .A2(new_n330), .A3(new_n585), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n870), .A2(new_n585), .A3(new_n871), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n905), .A2(new_n906), .A3(G190gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n905), .B2(G190gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(G1351gat));
  NAND2_X1  g708(.A1(new_n833), .A2(new_n425), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT124), .Z(new_n911));
  AND3_X1   g710(.A1(new_n867), .A2(new_n494), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(G197gat), .B1(new_n912), .B2(new_n711), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n668), .A2(new_n494), .A3(new_n425), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT125), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n915), .A2(G197gat), .A3(new_n711), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n913), .B1(new_n853), .B2(new_n916), .ZN(G1352gat));
  NAND3_X1  g716(.A1(new_n912), .A2(new_n625), .A3(new_n632), .ZN(new_n918));
  XOR2_X1   g717(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n853), .A2(new_n632), .A3(new_n915), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n625), .B2(new_n921), .ZN(G1353gat));
  INV_X1    g721(.A(G211gat), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n914), .A2(new_n710), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n853), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n710), .A2(new_n348), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n927), .B(new_n929), .C1(new_n925), .C2(new_n930), .ZN(G1354gat));
  AOI21_X1  g730(.A(G218gat), .B1(new_n912), .B2(new_n585), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n915), .A2(G218gat), .A3(new_n585), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n853), .B2(new_n933), .ZN(G1355gat));
endmodule


