

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U549 ( .A(n694), .B(n693), .ZN(n744) );
  INV_X1 U550 ( .A(KEYINPUT31), .ZN(n693) );
  NOR2_X1 U551 ( .A1(G651), .A2(G543), .ZN(n635) );
  NOR2_X2 U552 ( .A1(G2104), .A2(n517), .ZN(n596) );
  XNOR2_X2 U553 ( .A(n514), .B(n513), .ZN(n598) );
  INV_X1 U554 ( .A(KEYINPUT101), .ZN(n684) );
  XNOR2_X1 U555 ( .A(n684), .B(KEYINPUT30), .ZN(n685) );
  XNOR2_X1 U556 ( .A(n686), .B(n685), .ZN(n687) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n725) );
  XNOR2_X1 U558 ( .A(n726), .B(n725), .ZN(n729) );
  NOR2_X1 U559 ( .A1(G1966), .A2(n775), .ZN(n731) );
  XNOR2_X1 U560 ( .A(n682), .B(KEYINPUT64), .ZN(n706) );
  BUF_X1 U561 ( .A(n706), .Z(n735) );
  AND2_X1 U562 ( .A1(n517), .A2(G2104), .ZN(n518) );
  XNOR2_X1 U563 ( .A(n518), .B(KEYINPUT68), .ZN(n591) );
  NOR2_X1 U564 ( .A1(G651), .A2(n622), .ZN(n634) );
  XOR2_X1 U565 ( .A(KEYINPUT1), .B(n532), .Z(n642) );
  INV_X1 U566 ( .A(KEYINPUT66), .ZN(n525) );
  XNOR2_X1 U567 ( .A(KEYINPUT17), .B(KEYINPUT69), .ZN(n514) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n513) );
  NAND2_X1 U569 ( .A1(G137), .A2(n598), .ZN(n516) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n589) );
  NAND2_X1 U571 ( .A1(G113), .A2(n589), .ZN(n515) );
  NAND2_X1 U572 ( .A1(n516), .A2(n515), .ZN(n521) );
  INV_X1 U573 ( .A(G2105), .ZN(n517) );
  NAND2_X1 U574 ( .A1(n591), .A2(G101), .ZN(n519) );
  XNOR2_X1 U575 ( .A(n519), .B(KEYINPUT23), .ZN(n520) );
  NOR2_X1 U576 ( .A1(n521), .A2(n520), .ZN(n524) );
  NAND2_X1 U577 ( .A1(G125), .A2(n596), .ZN(n522) );
  XOR2_X1 U578 ( .A(KEYINPUT67), .B(n522), .Z(n523) );
  NAND2_X1 U579 ( .A1(n524), .A2(n523), .ZN(n526) );
  XNOR2_X2 U580 ( .A(n526), .B(n525), .ZN(G160) );
  AND2_X1 U581 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U582 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U583 ( .A(KEYINPUT71), .B(KEYINPUT9), .ZN(n530) );
  NAND2_X1 U584 ( .A1(G90), .A2(n635), .ZN(n528) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n622) );
  INV_X1 U586 ( .A(G651), .ZN(n531) );
  NOR2_X1 U587 ( .A1(n622), .A2(n531), .ZN(n638) );
  NAND2_X1 U588 ( .A1(G77), .A2(n638), .ZN(n527) );
  NAND2_X1 U589 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U590 ( .A(n530), .B(n529), .ZN(n536) );
  NAND2_X1 U591 ( .A1(G52), .A2(n634), .ZN(n534) );
  NOR2_X1 U592 ( .A1(G543), .A2(n531), .ZN(n532) );
  NAND2_X1 U593 ( .A1(G64), .A2(n642), .ZN(n533) );
  NAND2_X1 U594 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U595 ( .A1(n536), .A2(n535), .ZN(G171) );
  NAND2_X1 U596 ( .A1(G51), .A2(n634), .ZN(n538) );
  NAND2_X1 U597 ( .A1(G63), .A2(n642), .ZN(n537) );
  NAND2_X1 U598 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U599 ( .A(KEYINPUT6), .B(n539), .Z(n547) );
  NAND2_X1 U600 ( .A1(n638), .A2(G76), .ZN(n540) );
  XNOR2_X1 U601 ( .A(KEYINPUT75), .B(n540), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n635), .A2(G89), .ZN(n541) );
  XOR2_X1 U603 ( .A(n541), .B(KEYINPUT4), .Z(n542) );
  NOR2_X1 U604 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U605 ( .A(KEYINPUT76), .B(n544), .Z(n545) );
  XNOR2_X1 U606 ( .A(KEYINPUT5), .B(n545), .ZN(n546) );
  NAND2_X1 U607 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U608 ( .A(KEYINPUT7), .B(n548), .ZN(G168) );
  XOR2_X1 U609 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U610 ( .A1(G7), .A2(G661), .ZN(n549) );
  XNOR2_X1 U611 ( .A(n549), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U612 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n551) );
  INV_X1 U613 ( .A(G223), .ZN(n840) );
  NAND2_X1 U614 ( .A1(G567), .A2(n840), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(G234) );
  NAND2_X1 U616 ( .A1(n635), .A2(G81), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(KEYINPUT12), .ZN(n554) );
  NAND2_X1 U618 ( .A1(G68), .A2(n638), .ZN(n553) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(KEYINPUT13), .ZN(n557) );
  NAND2_X1 U621 ( .A1(G43), .A2(n634), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U623 ( .A1(n642), .A2(G56), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT14), .B(n558), .Z(n559) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n1014) );
  NAND2_X1 U626 ( .A1(n1014), .A2(G860), .ZN(G153) );
  INV_X1 U627 ( .A(G171), .ZN(G301) );
  NAND2_X1 U628 ( .A1(G54), .A2(n634), .ZN(n562) );
  NAND2_X1 U629 ( .A1(G79), .A2(n638), .ZN(n561) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G66), .A2(n642), .ZN(n564) );
  NAND2_X1 U632 ( .A1(G92), .A2(n635), .ZN(n563) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U634 ( .A(n565), .B(KEYINPUT73), .Z(n566) );
  NOR2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U636 ( .A(KEYINPUT15), .B(n568), .Z(n569) );
  XOR2_X1 U637 ( .A(KEYINPUT74), .B(n569), .Z(n995) );
  NOR2_X1 U638 ( .A1(n995), .A2(G868), .ZN(n571) );
  INV_X1 U639 ( .A(G868), .ZN(n653) );
  NOR2_X1 U640 ( .A1(n653), .A2(G301), .ZN(n570) );
  NOR2_X1 U641 ( .A1(n571), .A2(n570), .ZN(G284) );
  NAND2_X1 U642 ( .A1(G53), .A2(n634), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G65), .A2(n642), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U645 ( .A1(G91), .A2(n635), .ZN(n575) );
  NAND2_X1 U646 ( .A1(G78), .A2(n638), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n1001) );
  INV_X1 U649 ( .A(n1001), .ZN(G299) );
  XNOR2_X1 U650 ( .A(KEYINPUT77), .B(G868), .ZN(n578) );
  NOR2_X1 U651 ( .A1(G286), .A2(n578), .ZN(n580) );
  NOR2_X1 U652 ( .A1(G868), .A2(G299), .ZN(n579) );
  NOR2_X1 U653 ( .A1(n580), .A2(n579), .ZN(G297) );
  INV_X1 U654 ( .A(G860), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n581), .A2(G559), .ZN(n582) );
  INV_X1 U656 ( .A(n995), .ZN(n912) );
  NAND2_X1 U657 ( .A1(n582), .A2(n912), .ZN(n583) );
  XNOR2_X1 U658 ( .A(n583), .B(KEYINPUT78), .ZN(n584) );
  XNOR2_X1 U659 ( .A(KEYINPUT16), .B(n584), .ZN(G148) );
  NAND2_X1 U660 ( .A1(n1014), .A2(n653), .ZN(n587) );
  NOR2_X1 U661 ( .A1(G559), .A2(n653), .ZN(n585) );
  NAND2_X1 U662 ( .A1(n585), .A2(n912), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U664 ( .A(KEYINPUT79), .B(n588), .ZN(G282) );
  NAND2_X1 U665 ( .A1(G111), .A2(n589), .ZN(n590) );
  XNOR2_X1 U666 ( .A(n590), .B(KEYINPUT80), .ZN(n595) );
  INV_X1 U667 ( .A(n591), .ZN(n592) );
  INV_X1 U668 ( .A(n592), .ZN(n898) );
  NAND2_X1 U669 ( .A1(n898), .A2(G99), .ZN(n593) );
  XOR2_X1 U670 ( .A(KEYINPUT81), .B(n593), .Z(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G123), .A2(n596), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n597), .B(KEYINPUT18), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n598), .A2(G135), .ZN(n599) );
  NAND2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n978) );
  XOR2_X1 U677 ( .A(n978), .B(G2096), .Z(n603) );
  XNOR2_X1 U678 ( .A(KEYINPUT82), .B(n603), .ZN(n604) );
  NOR2_X1 U679 ( .A1(G2100), .A2(n604), .ZN(n605) );
  XNOR2_X1 U680 ( .A(KEYINPUT83), .B(n605), .ZN(G156) );
  NAND2_X1 U681 ( .A1(G55), .A2(n634), .ZN(n607) );
  NAND2_X1 U682 ( .A1(G67), .A2(n642), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U684 ( .A(KEYINPUT84), .B(n608), .ZN(n612) );
  NAND2_X1 U685 ( .A1(G93), .A2(n635), .ZN(n610) );
  NAND2_X1 U686 ( .A1(G80), .A2(n638), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n611) );
  OR2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n654) );
  NAND2_X1 U689 ( .A1(G559), .A2(n912), .ZN(n651) );
  XOR2_X1 U690 ( .A(n1014), .B(n651), .Z(n613) );
  NOR2_X1 U691 ( .A1(G860), .A2(n613), .ZN(n614) );
  XOR2_X1 U692 ( .A(n654), .B(n614), .Z(G145) );
  NAND2_X1 U693 ( .A1(G85), .A2(n635), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G72), .A2(n638), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n634), .A2(G47), .ZN(n617) );
  XOR2_X1 U697 ( .A(KEYINPUT70), .B(n617), .Z(n618) );
  NOR2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n642), .A2(G60), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(G290) );
  NAND2_X1 U701 ( .A1(G49), .A2(n634), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G87), .A2(n622), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U704 ( .A1(n642), .A2(n625), .ZN(n627) );
  NAND2_X1 U705 ( .A1(G651), .A2(G74), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(G288) );
  NAND2_X1 U707 ( .A1(G88), .A2(n635), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G75), .A2(n638), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G50), .A2(n634), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G62), .A2(n642), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U713 ( .A1(n633), .A2(n632), .ZN(G166) );
  NAND2_X1 U714 ( .A1(G48), .A2(n634), .ZN(n637) );
  NAND2_X1 U715 ( .A1(G86), .A2(n635), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n638), .A2(G73), .ZN(n639) );
  XOR2_X1 U718 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n642), .A2(G61), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(G305) );
  XNOR2_X1 U722 ( .A(G288), .B(KEYINPUT19), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n1001), .B(G166), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n646), .B(n645), .ZN(n647) );
  XOR2_X1 U725 ( .A(n647), .B(G305), .Z(n648) );
  XNOR2_X1 U726 ( .A(G290), .B(n648), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n1014), .B(n654), .ZN(n649) );
  XNOR2_X1 U728 ( .A(n650), .B(n649), .ZN(n909) );
  XOR2_X1 U729 ( .A(n909), .B(n651), .Z(n652) );
  NAND2_X1 U730 ( .A1(G868), .A2(n652), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n656), .A2(n655), .ZN(G295) );
  NAND2_X1 U733 ( .A1(G2078), .A2(G2084), .ZN(n657) );
  XNOR2_X1 U734 ( .A(n657), .B(KEYINPUT85), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n658), .B(KEYINPUT20), .ZN(n659) );
  NAND2_X1 U736 ( .A1(n659), .A2(G2090), .ZN(n660) );
  XNOR2_X1 U737 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U738 ( .A1(n661), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U740 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n663) );
  NAND2_X1 U741 ( .A1(G132), .A2(G82), .ZN(n662) );
  XNOR2_X1 U742 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n664), .A2(G96), .ZN(n665) );
  NOR2_X1 U744 ( .A1(n665), .A2(G218), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(KEYINPUT87), .ZN(n844) );
  NAND2_X1 U746 ( .A1(n844), .A2(G2106), .ZN(n670) );
  NAND2_X1 U747 ( .A1(G69), .A2(G120), .ZN(n667) );
  NOR2_X1 U748 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U749 ( .A1(G108), .A2(n668), .ZN(n845) );
  NAND2_X1 U750 ( .A1(n845), .A2(G567), .ZN(n669) );
  NAND2_X1 U751 ( .A1(n670), .A2(n669), .ZN(n846) );
  NAND2_X1 U752 ( .A1(G483), .A2(G661), .ZN(n671) );
  NOR2_X1 U753 ( .A1(n846), .A2(n671), .ZN(n843) );
  NAND2_X1 U754 ( .A1(n843), .A2(G36), .ZN(G176) );
  NAND2_X1 U755 ( .A1(n598), .A2(G138), .ZN(n673) );
  NAND2_X1 U756 ( .A1(G102), .A2(n898), .ZN(n672) );
  NAND2_X1 U757 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U758 ( .A(KEYINPUT88), .B(n674), .ZN(n678) );
  NAND2_X1 U759 ( .A1(G126), .A2(n596), .ZN(n676) );
  NAND2_X1 U760 ( .A1(G114), .A2(n589), .ZN(n675) );
  NAND2_X1 U761 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U762 ( .A1(n678), .A2(n677), .ZN(G164) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  NOR2_X1 U764 ( .A1(G2090), .A2(G303), .ZN(n679) );
  NAND2_X1 U765 ( .A1(G8), .A2(n679), .ZN(n680) );
  XNOR2_X1 U766 ( .A(n680), .B(KEYINPUT104), .ZN(n751) );
  NAND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n793) );
  XOR2_X1 U768 ( .A(KEYINPUT94), .B(n793), .Z(n681) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n794) );
  NAND2_X1 U770 ( .A1(n681), .A2(n794), .ZN(n682) );
  NAND2_X1 U771 ( .A1(n735), .A2(G8), .ZN(n775) );
  NOR2_X1 U772 ( .A1(n735), .A2(G2084), .ZN(n730) );
  NOR2_X1 U773 ( .A1(n731), .A2(n730), .ZN(n683) );
  NAND2_X1 U774 ( .A1(G8), .A2(n683), .ZN(n686) );
  NOR2_X1 U775 ( .A1(G168), .A2(n687), .ZN(n692) );
  INV_X1 U776 ( .A(n706), .ZN(n713) );
  XNOR2_X1 U777 ( .A(G1961), .B(KEYINPUT96), .ZN(n931) );
  NOR2_X1 U778 ( .A1(n713), .A2(n931), .ZN(n688) );
  XNOR2_X1 U779 ( .A(n688), .B(KEYINPUT97), .ZN(n690) );
  XNOR2_X1 U780 ( .A(G2078), .B(KEYINPUT25), .ZN(n947) );
  NAND2_X1 U781 ( .A1(n947), .A2(n713), .ZN(n689) );
  NAND2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n727) );
  NOR2_X1 U783 ( .A1(G171), .A2(n727), .ZN(n691) );
  NOR2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n694) );
  NAND2_X1 U785 ( .A1(G2072), .A2(n713), .ZN(n695) );
  XNOR2_X1 U786 ( .A(n695), .B(KEYINPUT27), .ZN(n697) );
  XOR2_X1 U787 ( .A(G1956), .B(KEYINPUT98), .Z(n926) );
  NOR2_X1 U788 ( .A1(n713), .A2(n926), .ZN(n696) );
  NOR2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n700) );
  NOR2_X1 U790 ( .A1(n700), .A2(n1001), .ZN(n699) );
  XNOR2_X1 U791 ( .A(KEYINPUT28), .B(KEYINPUT99), .ZN(n698) );
  XNOR2_X1 U792 ( .A(n699), .B(n698), .ZN(n724) );
  NAND2_X1 U793 ( .A1(n700), .A2(n1001), .ZN(n722) );
  NAND2_X1 U794 ( .A1(G1996), .A2(n713), .ZN(n703) );
  INV_X1 U795 ( .A(n703), .ZN(n702) );
  INV_X1 U796 ( .A(KEYINPUT26), .ZN(n701) );
  NAND2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U798 ( .A1(KEYINPUT26), .A2(n703), .ZN(n704) );
  NAND2_X1 U799 ( .A1(n705), .A2(n704), .ZN(n710) );
  NAND2_X1 U800 ( .A1(n706), .A2(G1341), .ZN(n707) );
  XNOR2_X1 U801 ( .A(KEYINPUT100), .B(n707), .ZN(n708) );
  AND2_X1 U802 ( .A1(n708), .A2(n1014), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n712) );
  INV_X1 U804 ( .A(KEYINPUT65), .ZN(n711) );
  XNOR2_X1 U805 ( .A(n712), .B(n711), .ZN(n717) );
  AND2_X1 U806 ( .A1(n735), .A2(G1348), .ZN(n715) );
  AND2_X1 U807 ( .A1(n713), .A2(G2067), .ZN(n714) );
  NOR2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n912), .A2(n718), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n717), .A2(n716), .ZN(n720) );
  OR2_X1 U811 ( .A1(n718), .A2(n912), .ZN(n719) );
  NAND2_X1 U812 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n726) );
  NAND2_X1 U815 ( .A1(n727), .A2(G171), .ZN(n728) );
  NAND2_X1 U816 ( .A1(n729), .A2(n728), .ZN(n742) );
  AND2_X1 U817 ( .A1(n744), .A2(n742), .ZN(n734) );
  AND2_X1 U818 ( .A1(G8), .A2(n730), .ZN(n732) );
  OR2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n733) );
  OR2_X1 U820 ( .A1(n734), .A2(n733), .ZN(n755) );
  INV_X1 U821 ( .A(G8), .ZN(n741) );
  NOR2_X1 U822 ( .A1(n735), .A2(G2090), .ZN(n737) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n775), .ZN(n736) );
  NOR2_X1 U824 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U825 ( .A(n738), .B(KEYINPUT102), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n739), .A2(G303), .ZN(n740) );
  OR2_X1 U827 ( .A1(n741), .A2(n740), .ZN(n745) );
  AND2_X1 U828 ( .A1(n742), .A2(n745), .ZN(n743) );
  NAND2_X1 U829 ( .A1(n744), .A2(n743), .ZN(n748) );
  INV_X1 U830 ( .A(n745), .ZN(n746) );
  OR2_X1 U831 ( .A1(n746), .A2(G286), .ZN(n747) );
  NAND2_X1 U832 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U833 ( .A(n749), .B(KEYINPUT32), .ZN(n757) );
  NAND2_X1 U834 ( .A1(n755), .A2(n757), .ZN(n750) );
  NAND2_X1 U835 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U836 ( .A1(n752), .A2(n775), .ZN(n771) );
  XOR2_X1 U837 ( .A(G1981), .B(G305), .Z(n1009) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n1000) );
  INV_X1 U839 ( .A(n1000), .ZN(n753) );
  OR2_X1 U840 ( .A1(n775), .A2(n753), .ZN(n759) );
  INV_X1 U841 ( .A(n759), .ZN(n754) );
  AND2_X1 U842 ( .A1(n755), .A2(n754), .ZN(n756) );
  AND2_X1 U843 ( .A1(n757), .A2(n756), .ZN(n763) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n764) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U846 ( .A1(n764), .A2(n758), .ZN(n1006) );
  OR2_X1 U847 ( .A1(n759), .A2(n1006), .ZN(n761) );
  INV_X1 U848 ( .A(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n767) );
  NAND2_X1 U851 ( .A1(n764), .A2(KEYINPUT33), .ZN(n765) );
  NOR2_X1 U852 ( .A1(n765), .A2(n775), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n1009), .A2(n768), .ZN(n769) );
  XOR2_X1 U855 ( .A(KEYINPUT103), .B(n769), .Z(n770) );
  NAND2_X1 U856 ( .A1(n771), .A2(n770), .ZN(n821) );
  NOR2_X1 U857 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XNOR2_X1 U858 ( .A(n772), .B(KEYINPUT24), .ZN(n773) );
  XNOR2_X1 U859 ( .A(KEYINPUT95), .B(n773), .ZN(n774) );
  NOR2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n819) );
  NAND2_X1 U861 ( .A1(G129), .A2(n596), .ZN(n777) );
  NAND2_X1 U862 ( .A1(G117), .A2(n589), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U864 ( .A(KEYINPUT92), .B(n778), .ZN(n782) );
  NAND2_X1 U865 ( .A1(n898), .A2(G105), .ZN(n779) );
  XNOR2_X1 U866 ( .A(n779), .B(KEYINPUT93), .ZN(n780) );
  XNOR2_X1 U867 ( .A(n780), .B(KEYINPUT38), .ZN(n781) );
  NOR2_X1 U868 ( .A1(n782), .A2(n781), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n598), .A2(G141), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n887) );
  NOR2_X1 U871 ( .A1(G1996), .A2(n887), .ZN(n974) );
  AND2_X1 U872 ( .A1(n887), .A2(G1996), .ZN(n792) );
  NAND2_X1 U873 ( .A1(n596), .A2(G119), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G95), .A2(n898), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G131), .A2(n598), .ZN(n788) );
  NAND2_X1 U877 ( .A1(G107), .A2(n589), .ZN(n787) );
  NAND2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n886) );
  INV_X1 U880 ( .A(G1991), .ZN(n796) );
  NOR2_X1 U881 ( .A1(n886), .A2(n796), .ZN(n791) );
  NOR2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n983) );
  NOR2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n822) );
  INV_X1 U884 ( .A(n822), .ZN(n795) );
  NOR2_X1 U885 ( .A1(n983), .A2(n795), .ZN(n824) );
  NOR2_X1 U886 ( .A1(G1986), .A2(G290), .ZN(n797) );
  AND2_X1 U887 ( .A1(n796), .A2(n886), .ZN(n979) );
  NOR2_X1 U888 ( .A1(n797), .A2(n979), .ZN(n798) );
  NOR2_X1 U889 ( .A1(n824), .A2(n798), .ZN(n799) );
  NOR2_X1 U890 ( .A1(n974), .A2(n799), .ZN(n800) );
  XNOR2_X1 U891 ( .A(n800), .B(KEYINPUT39), .ZN(n813) );
  XNOR2_X1 U892 ( .A(G2067), .B(KEYINPUT37), .ZN(n814) );
  XNOR2_X1 U893 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n805) );
  NAND2_X1 U894 ( .A1(G128), .A2(n596), .ZN(n802) );
  NAND2_X1 U895 ( .A1(G116), .A2(n589), .ZN(n801) );
  NAND2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U897 ( .A(n803), .B(KEYINPUT35), .ZN(n804) );
  XNOR2_X1 U898 ( .A(n805), .B(n804), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n598), .A2(G140), .ZN(n807) );
  NAND2_X1 U900 ( .A1(G104), .A2(n898), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U902 ( .A(KEYINPUT34), .B(n808), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U904 ( .A(KEYINPUT36), .B(n811), .ZN(n885) );
  NOR2_X1 U905 ( .A1(n814), .A2(n885), .ZN(n812) );
  XNOR2_X1 U906 ( .A(n812), .B(KEYINPUT91), .ZN(n971) );
  NAND2_X1 U907 ( .A1(n813), .A2(n971), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n885), .A2(n814), .ZN(n982) );
  NAND2_X1 U909 ( .A1(n815), .A2(n982), .ZN(n816) );
  XOR2_X1 U910 ( .A(KEYINPUT105), .B(n816), .Z(n817) );
  NAND2_X1 U911 ( .A1(n817), .A2(n822), .ZN(n827) );
  INV_X1 U912 ( .A(n827), .ZN(n818) );
  OR2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n829) );
  XOR2_X1 U915 ( .A(G1986), .B(G290), .Z(n1002) );
  NAND2_X1 U916 ( .A1(n1002), .A2(n971), .ZN(n823) );
  AND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n825) );
  OR2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n826) );
  AND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U920 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U921 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U922 ( .A(G1341), .B(G2454), .ZN(n831) );
  XNOR2_X1 U923 ( .A(n831), .B(G2430), .ZN(n832) );
  XNOR2_X1 U924 ( .A(n832), .B(G1348), .ZN(n838) );
  XOR2_X1 U925 ( .A(G2443), .B(G2427), .Z(n834) );
  XNOR2_X1 U926 ( .A(G2438), .B(G2446), .ZN(n833) );
  XNOR2_X1 U927 ( .A(n834), .B(n833), .ZN(n836) );
  XOR2_X1 U928 ( .A(G2451), .B(G2435), .Z(n835) );
  XNOR2_X1 U929 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U930 ( .A(n838), .B(n837), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n839), .A2(G14), .ZN(n915) );
  XOR2_X1 U932 ( .A(KEYINPUT106), .B(n915), .Z(G401) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n840), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U935 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U937 ( .A1(n843), .A2(n842), .ZN(G188) );
  NOR2_X1 U938 ( .A1(n845), .A2(n844), .ZN(G325) );
  XNOR2_X1 U939 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  INV_X1 U940 ( .A(n846), .ZN(G319) );
  XOR2_X1 U941 ( .A(G2100), .B(G2096), .Z(n848) );
  XNOR2_X1 U942 ( .A(G2090), .B(KEYINPUT43), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U944 ( .A(n849), .B(KEYINPUT108), .Z(n851) );
  XNOR2_X1 U945 ( .A(G2072), .B(G2678), .ZN(n850) );
  XNOR2_X1 U946 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U947 ( .A(KEYINPUT42), .B(G2084), .Z(n853) );
  XNOR2_X1 U948 ( .A(G2078), .B(G2067), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U950 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(G1986), .Z(n857) );
  XNOR2_X1 U952 ( .A(G1966), .B(G1971), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U954 ( .A(n858), .B(G1991), .Z(n860) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1976), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U957 ( .A(G2474), .B(G1981), .Z(n862) );
  XNOR2_X1 U958 ( .A(G1961), .B(G1956), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U961 ( .A1(n898), .A2(G100), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n865), .B(KEYINPUT110), .ZN(n868) );
  NAND2_X1 U963 ( .A1(G112), .A2(n589), .ZN(n866) );
  XOR2_X1 U964 ( .A(KEYINPUT109), .B(n866), .Z(n867) );
  NAND2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U966 ( .A1(G124), .A2(n596), .ZN(n869) );
  XNOR2_X1 U967 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n598), .A2(G136), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U970 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U971 ( .A1(n598), .A2(G139), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G103), .A2(n898), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n882) );
  NAND2_X1 U974 ( .A1(n589), .A2(G115), .ZN(n876) );
  XNOR2_X1 U975 ( .A(n876), .B(KEYINPUT114), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G127), .A2(n596), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U978 ( .A(KEYINPUT115), .B(n879), .ZN(n880) );
  XNOR2_X1 U979 ( .A(KEYINPUT47), .B(n880), .ZN(n881) );
  NOR2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n967) );
  XNOR2_X1 U981 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n883), .B(KEYINPUT116), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n889) );
  XOR2_X1 U984 ( .A(n887), .B(n886), .Z(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U986 ( .A(n890), .B(n978), .Z(n892) );
  XNOR2_X1 U987 ( .A(G164), .B(G162), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n905) );
  NAND2_X1 U989 ( .A1(G118), .A2(n589), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n893), .B(KEYINPUT112), .ZN(n896) );
  NAND2_X1 U991 ( .A1(G130), .A2(n596), .ZN(n894) );
  XOR2_X1 U992 ( .A(KEYINPUT111), .B(n894), .Z(n895) );
  NAND2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n903) );
  NAND2_X1 U994 ( .A1(n598), .A2(G142), .ZN(n897) );
  XOR2_X1 U995 ( .A(KEYINPUT113), .B(n897), .Z(n900) );
  NAND2_X1 U996 ( .A1(G106), .A2(n898), .ZN(n899) );
  NAND2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U998 ( .A(n901), .B(KEYINPUT45), .Z(n902) );
  NOR2_X1 U999 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n905), .B(n904), .Z(n906) );
  XNOR2_X1 U1001 ( .A(n967), .B(n906), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n907), .B(G160), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n908), .ZN(G395) );
  XOR2_X1 U1004 ( .A(KEYINPUT117), .B(n909), .Z(n911) );
  XNOR2_X1 U1005 ( .A(G171), .B(G286), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n913) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n914), .ZN(G397) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n915), .ZN(n918) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(G225) );
  XOR2_X1 U1015 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  XNOR2_X1 U1017 ( .A(G1348), .B(KEYINPUT59), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(n921), .B(G4), .ZN(n925) );
  XNOR2_X1 U1019 ( .A(G1341), .B(G19), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(G6), .B(G1981), .ZN(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n929) );
  XOR2_X1 U1023 ( .A(G20), .B(n926), .Z(n927) );
  XNOR2_X1 U1024 ( .A(KEYINPUT126), .B(n927), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(KEYINPUT60), .B(n930), .ZN(n935) );
  XNOR2_X1 U1027 ( .A(n931), .B(G5), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(G21), .B(G1966), .ZN(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n942) );
  XNOR2_X1 U1031 ( .A(G1971), .B(G22), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(G23), .B(G1976), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n939) );
  XOR2_X1 U1034 ( .A(G1986), .B(G24), .Z(n938) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(KEYINPUT58), .B(n940), .ZN(n941) );
  NOR2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(n943), .B(KEYINPUT61), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(G16), .B(KEYINPUT125), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(G11), .A2(n946), .ZN(n994) );
  XNOR2_X1 U1042 ( .A(G1991), .B(G25), .ZN(n956) );
  XNOR2_X1 U1043 ( .A(G27), .B(n947), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n949) );
  XNOR2_X1 U1045 ( .A(G1996), .B(G32), .ZN(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(G33), .B(G2072), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(KEYINPUT121), .B(n954), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(G28), .A2(n957), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(n958), .B(KEYINPUT53), .ZN(n961) );
  XOR2_X1 U1054 ( .A(G2084), .B(KEYINPUT54), .Z(n959) );
  XNOR2_X1 U1055 ( .A(G34), .B(n959), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G35), .B(G2090), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(G29), .A2(n964), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(n965), .B(KEYINPUT55), .ZN(n992) );
  XNOR2_X1 U1061 ( .A(G164), .B(G2078), .ZN(n966) );
  XNOR2_X1 U1062 ( .A(n966), .B(KEYINPUT119), .ZN(n969) );
  XOR2_X1 U1063 ( .A(G2072), .B(n967), .Z(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n970), .B(KEYINPUT50), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n977) );
  XOR2_X1 U1067 ( .A(G2090), .B(G162), .Z(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(n975), .B(KEYINPUT51), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n987) );
  XNOR2_X1 U1071 ( .A(G2084), .B(G160), .ZN(n981) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n985) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(KEYINPUT52), .B(n988), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(KEYINPUT120), .B(n989), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(G29), .A2(n990), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n1023) );
  XNOR2_X1 U1082 ( .A(KEYINPUT56), .B(G16), .ZN(n1020) );
  XNOR2_X1 U1083 ( .A(G301), .B(G1961), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(n995), .B(G1348), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(KEYINPUT122), .B(n998), .ZN(n1018) );
  NAND2_X1 U1087 ( .A1(G1971), .A2(G303), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1005) );
  XNOR2_X1 U1089 ( .A(n1001), .B(G1956), .ZN(n1003) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NAND2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(n1008), .B(KEYINPUT123), .ZN(n1013) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G168), .ZN(n1010) );
  NAND2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(n1011), .B(KEYINPUT57), .ZN(n1012) );
  NAND2_X1 U1097 ( .A1(n1013), .A2(n1012), .ZN(n1016) );
  XOR2_X1 U1098 ( .A(n1014), .B(G1341), .Z(n1015) );
  NOR2_X1 U1099 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1100 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1101 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1102 ( .A(n1021), .B(KEYINPUT124), .ZN(n1022) );
  NAND2_X1 U1103 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  XNOR2_X1 U1105 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1106 ( .A(G132), .ZN(G219) );
  INV_X1 U1107 ( .A(G120), .ZN(G236) );
  INV_X1 U1108 ( .A(G96), .ZN(G221) );
  INV_X1 U1109 ( .A(G82), .ZN(G220) );
  INV_X1 U1110 ( .A(G69), .ZN(G235) );
  INV_X1 U1111 ( .A(G108), .ZN(G238) );
endmodule

