//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n210), .A2(new_n211), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(new_n211), .B2(new_n210), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n219), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G87), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(G97), .B(G107), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n250), .A2(G223), .B1(G77), .B2(new_n248), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT66), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n252), .A2(new_n253), .A3(G222), .A4(new_n249), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n249), .ZN(new_n255));
  INV_X1    g0055(.A(G222), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT66), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n251), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  OAI211_X1 g0061(.A(G1), .B(G13), .C1(new_n244), .C2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n263), .B(KEYINPUT65), .C1(G41), .C2(G45), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n262), .A2(G274), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n267), .A2(KEYINPUT65), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n259), .A2(new_n267), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n269), .B1(G226), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n260), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G190), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n263), .A2(G20), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n212), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT67), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n279), .A3(new_n212), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n275), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G50), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n202), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n213), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(G20), .B2(new_n203), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n278), .A2(new_n280), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n282), .B(new_n285), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT9), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n273), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT69), .ZN(new_n297));
  INV_X1    g0097(.A(G200), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n272), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT10), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n273), .A2(new_n295), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n302), .B(new_n303), .C1(new_n304), .C2(new_n299), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n272), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(new_n294), .C1(G169), .C2(new_n272), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n301), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n252), .A2(G232), .A3(G1698), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n252), .A2(G226), .A3(new_n249), .ZN(new_n312));
  INV_X1    g0112(.A(G97), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n311), .B(new_n312), .C1(new_n244), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n259), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT13), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n265), .A2(new_n268), .B1(new_n270), .B2(G238), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n316), .B1(new_n315), .B2(new_n317), .ZN(new_n319));
  OAI21_X1  g0119(.A(G200), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n315), .A2(new_n317), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT13), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(G190), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n293), .ZN(new_n325));
  INV_X1    g0125(.A(G68), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G20), .ZN(new_n327));
  INV_X1    g0127(.A(G77), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n327), .B1(new_n287), .B2(new_n328), .C1(new_n290), .C2(new_n202), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT11), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n275), .A2(new_n277), .A3(new_n326), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT70), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n284), .A2(new_n326), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT12), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n325), .A2(KEYINPUT11), .A3(new_n329), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n332), .A2(new_n334), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n320), .A2(new_n324), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n318), .A2(new_n319), .ZN(new_n342));
  INV_X1    g0142(.A(G169), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(KEYINPUT71), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT14), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT14), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n344), .C1(new_n318), .C2(new_n319), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n342), .A2(G179), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n341), .B1(new_n350), .B2(new_n338), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n269), .B1(G244), .B2(new_n270), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n250), .A2(G238), .B1(G107), .B2(new_n248), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n252), .A2(G232), .A3(new_n249), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n259), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n306), .ZN(new_n358));
  INV_X1    g0158(.A(new_n277), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(G77), .A3(new_n274), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(G77), .B2(new_n283), .ZN(new_n361));
  INV_X1    g0161(.A(new_n286), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT68), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n365), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n363), .B1(new_n368), .B2(new_n287), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n361), .B1(new_n369), .B2(new_n277), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n352), .A2(new_n356), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(new_n343), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n358), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n357), .A2(G190), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n374), .B(new_n370), .C1(new_n298), .C2(new_n357), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n310), .A2(new_n351), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n252), .A2(G226), .A3(G1698), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n252), .A2(G223), .A3(new_n249), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G87), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n259), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n265), .A2(new_n268), .B1(new_n270), .B2(G232), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G169), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n381), .A2(new_n382), .A3(G179), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT7), .B1(new_n248), .B2(new_n213), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  AOI211_X1 g0188(.A(new_n388), .B(G20), .C1(new_n245), .C2(new_n247), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G58), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n326), .ZN(new_n392));
  OAI21_X1  g0192(.A(G20), .B1(new_n392), .B2(new_n201), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n289), .A2(G159), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n388), .B1(new_n252), .B2(G20), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n246), .A2(G33), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n401));
  OAI211_X1 g0201(.A(KEYINPUT7), .B(new_n213), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n326), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n398), .B1(new_n403), .B2(new_n395), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n397), .A2(new_n404), .A3(new_n277), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n286), .A2(new_n283), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n281), .B2(new_n286), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT72), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT72), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n409), .B(new_n406), .C1(new_n281), .C2(new_n286), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n405), .A2(KEYINPUT73), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT73), .B1(new_n405), .B2(new_n411), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n386), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n383), .A2(G200), .ZN(new_n415));
  XOR2_X1   g0215(.A(KEYINPUT74), .B(G190), .Z(new_n416));
  NAND3_X1  g0216(.A1(new_n381), .A2(new_n382), .A3(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n405), .A2(new_n415), .A3(new_n411), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT17), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n298), .B1(new_n381), .B2(new_n382), .ZN(new_n420));
  INV_X1    g0220(.A(new_n383), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n416), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(new_n405), .A4(new_n411), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n414), .A2(KEYINPUT18), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n426), .B(new_n386), .C1(new_n412), .C2(new_n413), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n376), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n245), .A2(new_n247), .A3(G244), .A4(new_n249), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT4), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n249), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G283), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n252), .A2(G250), .A3(G1698), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n432), .A2(new_n433), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n259), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT75), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(KEYINPUT75), .A3(new_n259), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n263), .B(G45), .C1(new_n261), .C2(KEYINPUT5), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT5), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G41), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n262), .B(G257), .C1(new_n442), .C2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n266), .A2(G1), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(G41), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .A4(G274), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT76), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n445), .A2(KEYINPUT76), .A3(new_n449), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n441), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G200), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n437), .A2(new_n452), .A3(new_n453), .ZN(new_n457));
  INV_X1    g0257(.A(G190), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G107), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G97), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT6), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n462), .B2(new_n238), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n464), .A2(new_n213), .B1(new_n328), .B2(new_n290), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n460), .B1(new_n399), .B2(new_n402), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n277), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n283), .A2(G97), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n263), .A2(G33), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n293), .A2(new_n283), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n468), .B1(new_n470), .B2(G97), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n459), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n456), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G116), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n244), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n245), .A2(new_n247), .A3(G238), .A4(new_n249), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT78), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n252), .A2(new_n480), .A3(G244), .A4(G1698), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n252), .A2(KEYINPUT78), .A3(G238), .A4(new_n249), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n245), .A2(new_n247), .A3(G244), .A4(G1698), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT79), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n479), .A2(new_n481), .A3(new_n482), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n259), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n262), .B(G250), .C1(G1), .C2(new_n266), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n446), .A2(G274), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n252), .A2(new_n213), .A3(G68), .ZN(new_n492));
  OR2_X1    g0292(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n213), .A2(G33), .A3(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NOR3_X1   g0298(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n493), .A2(G33), .A3(G97), .A4(new_n494), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n213), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n277), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n368), .A2(new_n284), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n368), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n470), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n491), .A2(new_n343), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n489), .B1(new_n485), .B2(new_n259), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n306), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n293), .A2(G87), .A3(new_n283), .A4(new_n469), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n502), .A2(new_n503), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n491), .B2(G200), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n508), .A2(G190), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n507), .A2(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n436), .A2(KEYINPUT75), .A3(new_n259), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT75), .B1(new_n436), .B2(new_n259), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n454), .B(new_n306), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT77), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT77), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n441), .A2(new_n519), .A3(new_n306), .A4(new_n454), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n457), .A2(new_n343), .B1(new_n467), .B2(new_n471), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n474), .A2(new_n514), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n252), .A2(G250), .A3(new_n249), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n252), .A2(G257), .A3(G1698), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G294), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n259), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n442), .A2(new_n444), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(new_n259), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G264), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n531), .A3(new_n449), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G200), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n527), .A2(new_n259), .B1(new_n530), .B2(G264), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(G190), .A3(new_n449), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT25), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n283), .B2(G107), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n284), .A2(KEYINPUT25), .A3(new_n460), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n470), .A2(G107), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT23), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n213), .B2(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n460), .A2(KEYINPUT23), .A3(G20), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n476), .A2(new_n213), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n245), .A2(new_n247), .A3(new_n213), .A4(G87), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT22), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT22), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n252), .A2(new_n549), .A3(new_n213), .A4(G87), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n546), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT24), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n277), .B1(new_n551), .B2(KEYINPUT24), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n540), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n536), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n534), .A2(G179), .A3(new_n449), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n343), .B1(new_n534), .B2(new_n449), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT81), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n532), .A2(G169), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n534), .A2(G179), .A3(new_n449), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT81), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n559), .A2(new_n563), .A3(new_n555), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT82), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n559), .A2(KEYINPUT82), .A3(new_n563), .A4(new_n555), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n556), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n245), .A2(new_n247), .A3(G257), .A4(new_n249), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n245), .A2(new_n247), .A3(G264), .A4(G1698), .ZN(new_n570));
  INV_X1    g0370(.A(G303), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n252), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n259), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n262), .B(G270), .C1(new_n442), .C2(new_n444), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n574), .A2(new_n449), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n343), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n283), .A2(G116), .A3(new_n469), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(new_n359), .B1(new_n475), .B2(new_n284), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n276), .A2(new_n212), .B1(G20), .B2(new_n475), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n434), .B(new_n213), .C1(G33), .C2(new_n313), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n579), .A2(KEYINPUT20), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT20), .B1(new_n579), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n576), .A2(KEYINPUT21), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n583), .A2(G179), .A3(new_n573), .A4(new_n575), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT21), .B1(new_n576), .B2(new_n583), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n573), .A2(new_n575), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n416), .ZN(new_n591));
  INV_X1    g0391(.A(new_n583), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n591), .B(new_n592), .C1(new_n298), .C2(new_n590), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n429), .A2(new_n523), .A3(new_n568), .A4(new_n594), .ZN(G372));
  NAND2_X1  g0395(.A1(new_n405), .A2(new_n411), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n386), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n426), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n405), .A2(new_n411), .B1(new_n384), .B2(new_n385), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT18), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n350), .A2(new_n338), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n358), .A2(new_n372), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n419), .A2(new_n424), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n340), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n601), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(new_n305), .A3(new_n301), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n609), .A2(new_n308), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n560), .A2(new_n561), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n555), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n556), .B1(new_n588), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n613), .A2(new_n522), .A3(new_n474), .A4(new_n514), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n506), .A2(new_n503), .A3(new_n502), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n509), .B(new_n615), .C1(G169), .C2(new_n508), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT26), .B1(new_n617), .B2(new_n514), .ZN(new_n618));
  INV_X1    g0418(.A(new_n511), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n513), .B(new_n619), .C1(new_n298), .C2(new_n508), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n522), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n614), .B(new_n616), .C1(new_n618), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n429), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n610), .A2(new_n625), .ZN(G369));
  AND2_X1   g0426(.A1(new_n213), .A2(G13), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n263), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n628), .A2(KEYINPUT27), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(KEYINPUT27), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(G213), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G343), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n633), .A2(new_n592), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n586), .B2(new_n587), .ZN(new_n635));
  INV_X1    g0435(.A(new_n594), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(new_n634), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT83), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT84), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n555), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n568), .B1(new_n642), .B2(new_n633), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n551), .A2(KEYINPUT24), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(new_n277), .A3(new_n552), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n611), .A2(KEYINPUT81), .B1(new_n645), .B2(new_n540), .ZN(new_n646));
  INV_X1    g0446(.A(new_n633), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n563), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n641), .A2(G330), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n588), .A2(new_n647), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n568), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n612), .A2(new_n647), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n650), .A2(new_n655), .ZN(G399));
  INV_X1    g0456(.A(new_n209), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(G41), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n499), .A2(new_n475), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(G1), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n216), .B2(new_n659), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT28), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT82), .B1(new_n646), .B2(new_n563), .ZN(new_n665));
  INV_X1    g0465(.A(new_n567), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n588), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n621), .A2(new_n556), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n474), .A2(new_n522), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT88), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT88), .B1(new_n474), .B2(new_n522), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n667), .B(new_n668), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n616), .B(KEYINPUT87), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n617), .A2(KEYINPUT26), .A3(new_n514), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n622), .B1(new_n522), .B2(new_n621), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT89), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(KEYINPUT29), .A4(new_n633), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT29), .ZN(new_n681));
  AOI211_X1 g0481(.A(new_n681), .B(new_n647), .C1(new_n673), .C2(new_n677), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n624), .A2(new_n633), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT89), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n680), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n568), .A2(new_n523), .A3(new_n594), .A4(new_n633), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n573), .A2(new_n575), .A3(G179), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n454), .A2(new_n687), .A3(new_n437), .A4(new_n534), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT85), .B1(new_n688), .B2(new_n491), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n532), .A2(new_n306), .A3(new_n589), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n508), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n689), .A2(KEYINPUT30), .B1(new_n455), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT30), .ZN(new_n693));
  OAI211_X1 g0493(.A(KEYINPUT85), .B(new_n693), .C1(new_n688), .C2(new_n491), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n633), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT86), .B1(new_n695), .B2(KEYINPUT31), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(KEYINPUT31), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n686), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n695), .A2(KEYINPUT86), .A3(KEYINPUT31), .ZN(new_n699));
  OAI21_X1  g0499(.A(G330), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT90), .B1(new_n685), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n685), .A2(KEYINPUT90), .A3(new_n700), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n664), .B1(new_n704), .B2(G1), .ZN(G364));
  NAND2_X1  g0505(.A1(new_n641), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n263), .B1(new_n627), .B2(G45), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n658), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n641), .A2(G330), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(G13), .A2(G33), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G20), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n639), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n212), .B1(G20), .B2(new_n343), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n657), .A2(new_n252), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(G45), .B2(new_n216), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(G45), .B2(new_n242), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n657), .A2(new_n248), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  XOR2_X1   g0524(.A(G355), .B(KEYINPUT91), .Z(new_n725));
  OAI22_X1  g0525(.A1(new_n724), .A2(new_n725), .B1(G116), .B2(new_n209), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n719), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n710), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n213), .A2(new_n306), .A3(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n458), .ZN(new_n730));
  INV_X1    g0530(.A(G311), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n248), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n416), .A2(new_n729), .ZN(new_n733));
  INV_X1    g0533(.A(G322), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n213), .A2(G179), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(G190), .A3(G200), .ZN(new_n736));
  OAI22_X1  g0536(.A1(new_n733), .A2(new_n734), .B1(new_n571), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G179), .A2(G200), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n213), .B1(new_n738), .B2(G190), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n732), .B(new_n737), .C1(G294), .C2(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n213), .A2(new_n306), .A3(new_n298), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT93), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(KEYINPUT93), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n743), .A2(new_n416), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G326), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n743), .A2(new_n458), .A3(new_n744), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT33), .B(G317), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n735), .A2(new_n458), .A3(G200), .ZN(new_n750));
  INV_X1    g0550(.A(G283), .ZN(new_n751));
  INV_X1    g0551(.A(G329), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n738), .A2(G20), .A3(new_n458), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT96), .Z(new_n755));
  NAND4_X1  g0555(.A1(new_n741), .A2(new_n746), .A3(new_n749), .A4(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G87), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n736), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n733), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n758), .B1(new_n759), .B2(G58), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(new_n313), .B2(new_n739), .ZN(new_n761));
  INV_X1    g0561(.A(new_n750), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n248), .B(new_n761), .C1(G107), .C2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n753), .ZN(new_n764));
  XOR2_X1   g0564(.A(KEYINPUT94), .B(G159), .Z(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT95), .Z(new_n767));
  INV_X1    g0567(.A(new_n745), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n763), .B1(KEYINPUT32), .B2(new_n767), .C1(new_n202), .C2(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n767), .A2(KEYINPUT32), .B1(G68), .B2(new_n747), .ZN(new_n770));
  INV_X1    g0570(.A(new_n730), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT92), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(KEYINPUT92), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n770), .B1(new_n328), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n756), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n728), .B1(new_n776), .B2(new_n718), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n711), .A2(new_n713), .B1(new_n717), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(G396));
  INV_X1    g0579(.A(new_n710), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n370), .A2(new_n633), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n604), .B1(new_n375), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n373), .A2(new_n647), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT97), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n683), .ZN(new_n786));
  INV_X1    g0586(.A(new_n616), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n675), .B2(new_n676), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n647), .B1(new_n788), .B2(new_n614), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n786), .A2(KEYINPUT98), .B1(new_n789), .B2(new_n784), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(KEYINPUT98), .B2(new_n786), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n780), .B1(new_n791), .B2(new_n700), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT99), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n792), .A2(new_n793), .B1(new_n700), .B2(new_n791), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n793), .B2(new_n792), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n718), .A2(new_n714), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n780), .B1(new_n328), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G132), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n252), .B1(new_n753), .B2(new_n798), .C1(new_n736), .C2(new_n202), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n750), .A2(new_n326), .B1(new_n739), .B2(new_n391), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n745), .A2(G137), .B1(new_n759), .B2(G143), .ZN(new_n801));
  INV_X1    g0601(.A(new_n747), .ZN(new_n802));
  INV_X1    g0602(.A(new_n765), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n801), .B1(new_n288), .B2(new_n802), .C1(new_n774), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT34), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n799), .B(new_n800), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n757), .A2(new_n750), .B1(new_n736), .B2(new_n460), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n248), .B1(new_n753), .B2(new_n731), .C1(new_n313), .C2(new_n739), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n808), .B(new_n809), .C1(G294), .C2(new_n759), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n768), .A2(new_n571), .B1(new_n802), .B2(new_n751), .ZN(new_n811));
  INV_X1    g0611(.A(new_n774), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(G116), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n806), .A2(new_n807), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n718), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n797), .B1(new_n814), .B2(new_n815), .C1(new_n784), .C2(new_n715), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n795), .A2(new_n816), .ZN(G384));
  INV_X1    g0617(.A(new_n464), .ZN(new_n818));
  OAI211_X1 g0618(.A(G116), .B(new_n214), .C1(new_n818), .C2(KEYINPUT35), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(KEYINPUT35), .B2(new_n818), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT36), .ZN(new_n821));
  OR3_X1    g0621(.A1(new_n216), .A2(new_n328), .A3(new_n392), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n202), .A2(G68), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n263), .B(G13), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n689), .A2(KEYINPUT30), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n691), .A2(new_n455), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n826), .A2(new_n694), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n647), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT31), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n695), .A2(KEYINPUT31), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n686), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n374), .A2(new_n370), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n357), .A2(new_n298), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n781), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n373), .ZN(new_n837));
  INV_X1    g0637(.A(new_n783), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n603), .A2(new_n647), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n339), .A2(new_n633), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n351), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n839), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n833), .A2(new_n844), .A3(KEYINPUT40), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n632), .B1(new_n412), .B2(new_n413), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT102), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n606), .A2(new_n848), .B1(new_n598), .B2(new_n600), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n419), .A2(new_n424), .A3(KEYINPUT102), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n418), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT73), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n596), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n405), .A2(KEYINPUT73), .A3(new_n411), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n853), .B1(new_n857), .B2(new_n386), .ZN(new_n858));
  AND4_X1   g0658(.A1(new_n405), .A2(new_n415), .A3(new_n411), .A4(new_n417), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n859), .A2(new_n599), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n847), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n847), .A2(new_n858), .B1(new_n861), .B2(KEYINPUT37), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n846), .B1(new_n851), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT103), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n397), .A2(new_n404), .A3(new_n325), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n411), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n632), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n386), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n855), .B2(new_n856), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n606), .B1(new_n870), .B2(new_n426), .ZN(new_n871));
  INV_X1    g0671(.A(new_n427), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n414), .A2(new_n847), .A3(new_n852), .A4(new_n418), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n866), .A2(new_n386), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n867), .A3(new_n418), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n873), .A2(KEYINPUT38), .A3(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n863), .A2(new_n864), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n864), .B1(new_n863), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n845), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n867), .B1(new_n425), .B2(new_n427), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n858), .A2(new_n847), .B1(KEYINPUT37), .B2(new_n876), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n846), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n885), .A2(KEYINPUT100), .A3(new_n879), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT100), .B1(new_n885), .B2(new_n879), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n833), .A2(new_n844), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n882), .B(G330), .C1(new_n889), .C2(KEYINPUT40), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n833), .A2(G330), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n429), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT104), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT100), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n883), .A2(new_n884), .A3(new_n846), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n873), .B2(new_n878), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n841), .B(new_n341), .C1(new_n350), .C2(new_n338), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n602), .A2(new_n633), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n784), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n695), .B(new_n830), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n905), .B2(new_n686), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n885), .A2(new_n879), .A3(KEYINPUT100), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n901), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n606), .A2(new_n848), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n601), .A3(new_n850), .ZN(new_n910));
  INV_X1    g0710(.A(new_n847), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n874), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT103), .B1(new_n915), .B2(new_n899), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n863), .A2(new_n864), .A3(new_n879), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n897), .A2(new_n908), .B1(new_n918), .B2(new_n845), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n429), .A3(new_n833), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n895), .A2(new_n896), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n429), .B(new_n680), .C1(new_n682), .C2(new_n684), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n610), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n896), .B1(new_n895), .B2(new_n920), .ZN(new_n926));
  OR3_X1    g0726(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n902), .A2(new_n903), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n624), .A2(new_n633), .A3(new_n784), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n928), .B1(new_n929), .B2(new_n838), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(new_n901), .A3(new_n907), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n885), .B2(new_n879), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n915), .A2(new_n899), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n933), .B1(new_n934), .B2(new_n932), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT101), .B1(new_n602), .B2(new_n647), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n602), .A2(KEYINPUT101), .A3(new_n647), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n931), .B1(new_n601), .B2(new_n632), .C1(new_n935), .C2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n925), .B1(new_n922), .B2(new_n926), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n927), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n263), .B2(new_n627), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n941), .B1(new_n927), .B2(new_n942), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n825), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT105), .ZN(G367));
  XNOR2_X1  g0747(.A(new_n669), .B(new_n670), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n472), .A2(new_n647), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n522), .B2(new_n633), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(new_n655), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT44), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n655), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT45), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n650), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n953), .A2(new_n650), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n652), .B1(new_n649), .B2(new_n651), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n706), .B(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n704), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n658), .B(KEYINPUT41), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n708), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n653), .A2(new_n948), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n948), .A2(new_n566), .A3(new_n567), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n647), .B1(new_n971), .B2(new_n522), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n514), .B1(new_n619), .B2(new_n633), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n787), .A2(new_n511), .A3(new_n647), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n970), .A2(new_n973), .B1(KEYINPUT43), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n977), .B(new_n978), .Z(new_n979));
  NAND2_X1  g0779(.A1(new_n958), .A2(new_n951), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n967), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n720), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n984), .A2(new_n235), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n719), .B1(new_n209), .B2(new_n368), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n710), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT107), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n812), .A2(G283), .B1(G311), .B2(new_n745), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n750), .A2(new_n313), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n248), .B1(new_n991), .B2(new_n753), .C1(new_n733), .C2(new_n571), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n990), .B(new_n992), .C1(G107), .C2(new_n740), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT108), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(KEYINPUT46), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n736), .A2(new_n475), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n736), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n997), .B(G116), .C1(new_n994), .C2(KEYINPUT46), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n747), .A2(G294), .B1(new_n998), .B2(new_n995), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n989), .A2(new_n993), .A3(new_n996), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(G137), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n736), .A2(new_n391), .B1(new_n1001), .B2(new_n753), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT109), .Z(new_n1003));
  AOI22_X1  g0803(.A1(new_n747), .A2(new_n765), .B1(new_n745), .B2(G143), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n739), .A2(new_n326), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n252), .B1(new_n750), .B2(new_n328), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G150), .C2(new_n759), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1004), .B(new_n1007), .C1(new_n202), .C2(new_n774), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1000), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT47), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n815), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n988), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n974), .A2(new_n975), .A3(new_n716), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n983), .A2(new_n1015), .ZN(G387));
  INV_X1    g0816(.A(new_n963), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n704), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n963), .A2(new_n702), .A3(new_n703), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n658), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n643), .A2(new_n648), .A3(new_n716), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n984), .B1(new_n232), .B2(G45), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n660), .B2(new_n723), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n286), .A2(G50), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT110), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n661), .B(new_n266), .C1(new_n326), .C2(new_n328), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1023), .A2(new_n1029), .B1(G107), .B2(new_n209), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n780), .B1(new_n1030), .B2(new_n719), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n736), .A2(new_n328), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n252), .B1(new_n753), .B2(new_n288), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n990), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n368), .A2(new_n739), .B1(new_n202), .B2(new_n733), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT111), .ZN(new_n1036));
  INV_X1    g0836(.A(G159), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .C1(new_n1037), .C2(new_n768), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n747), .A2(new_n362), .B1(G68), .B2(new_n771), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT112), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(new_n1036), .C2(new_n1035), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n747), .A2(G311), .B1(new_n745), .B2(G322), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n571), .B2(new_n774), .C1(new_n991), .C2(new_n733), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT48), .ZN(new_n1044));
  INV_X1    g0844(.A(G294), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1044), .B1(new_n751), .B2(new_n739), .C1(new_n1045), .C2(new_n736), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT49), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n252), .B1(new_n764), .B2(G326), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n475), .B2(new_n750), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1041), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1031), .B1(new_n1052), .B2(new_n815), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT113), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1017), .A2(new_n709), .B1(new_n1021), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1020), .A2(new_n1055), .ZN(G393));
  AOI21_X1  g0856(.A(new_n963), .B1(new_n702), .B2(new_n703), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n959), .A2(new_n960), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n659), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n959), .A2(KEYINPUT114), .A3(new_n960), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(KEYINPUT114), .B2(new_n959), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1059), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n951), .A2(G20), .A3(new_n715), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n984), .A2(new_n239), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n719), .B1(new_n209), .B2(new_n313), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n248), .B1(new_n764), .B2(G143), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n326), .B2(new_n736), .C1(new_n757), .C2(new_n750), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT116), .Z(new_n1068));
  OAI22_X1  g0868(.A1(new_n768), .A2(new_n288), .B1(new_n733), .B2(new_n1037), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n747), .A2(G50), .B1(G77), .B2(new_n740), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n286), .B2(new_n774), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n745), .A2(G317), .B1(new_n759), .B2(G311), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT52), .Z(new_n1077));
  OAI221_X1 g0877(.A(new_n248), .B1(new_n753), .B2(new_n734), .C1(new_n750), .C2(new_n460), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n997), .A2(G283), .B1(new_n740), .B2(G116), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n1045), .B2(new_n730), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(G303), .C2(new_n747), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1072), .A2(new_n1075), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n710), .B1(new_n1064), .B2(new_n1065), .C1(new_n1082), .C2(new_n815), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1063), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1061), .B2(new_n709), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1062), .A2(new_n1085), .ZN(G390));
  OAI21_X1  g0886(.A(KEYINPUT39), .B1(new_n899), .B2(new_n900), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n863), .A2(new_n932), .A3(new_n879), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n939), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1087), .B(new_n1088), .C1(new_n930), .C2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(G330), .B(new_n844), .C1(new_n698), .C2(new_n699), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT117), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n937), .B2(new_n938), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT101), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n603), .A2(new_n1094), .A3(new_n633), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(KEYINPUT117), .A3(new_n936), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n880), .B2(new_n881), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n647), .B1(new_n673), .B2(new_n677), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n837), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n928), .B1(new_n1100), .B2(new_n838), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1090), .B(new_n1091), .C1(new_n1098), .C2(new_n1101), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n647), .B(new_n782), .C1(new_n673), .C2(new_n677), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1103), .A2(new_n783), .B1(new_n902), .B2(new_n903), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n916), .B2(new_n917), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n783), .B1(new_n789), .B2(new_n784), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n939), .B1(new_n1107), .B2(new_n928), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1104), .A2(new_n1106), .B1(new_n935), .B2(new_n1108), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n833), .A2(new_n844), .A3(G330), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1102), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n935), .A2(new_n714), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n796), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n710), .B1(new_n362), .B2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n252), .B(new_n758), .C1(G294), .C2(new_n764), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n762), .A2(G68), .B1(new_n740), .B2(G77), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(new_n475), .C2(new_n733), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n812), .A2(G97), .B1(G107), .B2(new_n747), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n751), .B2(new_n768), .ZN(new_n1121));
  XOR2_X1   g0921(.A(KEYINPUT54), .B(G143), .Z(new_n1122));
  AOI22_X1  g0922(.A1(new_n812), .A2(new_n1122), .B1(G137), .B2(new_n747), .ZN(new_n1123));
  INV_X1    g0923(.A(G128), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n768), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n759), .A2(G132), .B1(G50), .B2(new_n762), .ZN(new_n1126));
  INV_X1    g0926(.A(G125), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n252), .B1(new_n753), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G159), .B2(new_n740), .ZN(new_n1129));
  OR3_X1    g0929(.A1(new_n736), .A2(KEYINPUT53), .A3(new_n288), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT53), .B1(new_n736), .B2(new_n288), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1126), .A2(new_n1129), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1119), .A2(new_n1121), .B1(new_n1125), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1116), .B1(new_n1133), .B2(new_n718), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1113), .A2(new_n709), .B1(new_n1114), .B2(new_n1134), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n923), .A2(new_n610), .A3(new_n893), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n928), .B1(new_n891), .B2(new_n785), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n783), .B1(new_n1099), .B2(new_n837), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n1138), .A3(new_n1091), .ZN(new_n1139));
  OAI211_X1 g0939(.A(G330), .B(new_n784), .C1(new_n698), .C2(new_n699), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1110), .B1(new_n1140), .B2(new_n928), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1141), .B2(new_n1107), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1136), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n659), .B1(new_n1113), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1112), .A2(new_n1143), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT118), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1106), .A2(new_n1104), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1090), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1110), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1150), .A2(new_n1102), .A3(new_n1136), .A4(new_n1142), .ZN(new_n1151));
  AND4_X1   g0951(.A1(KEYINPUT118), .A2(new_n1151), .A3(new_n658), .A4(new_n1146), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1135), .B1(new_n1147), .B2(new_n1152), .ZN(G378));
  OAI21_X1  g0953(.A(new_n1136), .B1(new_n1112), .B2(new_n1143), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n309), .A2(new_n294), .A3(new_n632), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n294), .A2(new_n632), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n301), .A2(new_n305), .A3(new_n308), .A4(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1158), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n919), .B2(G330), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n908), .A2(new_n897), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT121), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1158), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(KEYINPUT121), .A3(new_n1159), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  AND4_X1   g0972(.A1(G330), .A2(new_n1165), .A3(new_n1172), .A4(new_n882), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n941), .B1(new_n1164), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n890), .A2(new_n1162), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1165), .A2(new_n1172), .A3(G330), .A4(new_n882), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(new_n940), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1154), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n659), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1175), .A2(new_n940), .A3(new_n1176), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n940), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1183), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n1154), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1154), .A2(new_n1174), .A3(KEYINPUT57), .A4(new_n1177), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT122), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1180), .A2(new_n1184), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1183), .A2(new_n709), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n710), .B1(G50), .B2(new_n1115), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n252), .A2(G41), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G50), .B(new_n1191), .C1(new_n244), .C2(new_n261), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1191), .B1(new_n751), .B2(new_n753), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1005), .B(new_n1193), .C1(new_n505), .C2(new_n771), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n747), .A2(G97), .B1(new_n745), .B2(G116), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n750), .A2(new_n391), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1032), .B(new_n1196), .C1(new_n759), .C2(G107), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT58), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1192), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G33), .B(G41), .C1(new_n764), .C2(G124), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n759), .A2(G128), .B1(new_n997), .B2(new_n1122), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT119), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n730), .A2(new_n1001), .B1(new_n288), .B2(new_n739), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n747), .B2(G132), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(new_n1127), .C2(new_n768), .ZN(new_n1206));
  XOR2_X1   g1006(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1207));
  OAI221_X1 g1007(.A(new_n1201), .B1(new_n803), .B2(new_n750), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1200), .B1(new_n1199), .B2(new_n1198), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1190), .B1(new_n1210), .B2(new_n718), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n1172), .B2(new_n715), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1189), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1188), .A2(new_n1213), .ZN(G375));
  OR2_X1    g1014(.A1(new_n1136), .A2(new_n1142), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n965), .B(KEYINPUT123), .Z(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n1143), .A3(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n747), .A2(new_n1122), .B1(G137), .B2(new_n759), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n798), .B2(new_n768), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT126), .Z(new_n1220));
  OAI21_X1  g1020(.A(new_n252), .B1(new_n753), .B2(new_n1124), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n997), .A2(G159), .B1(new_n740), .B2(G50), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n288), .B2(new_n730), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1220), .A2(new_n1196), .A3(new_n1221), .A4(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT125), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n248), .B1(new_n750), .B2(new_n328), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n745), .A2(G294), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n460), .A2(new_n774), .B1(new_n802), .B2(new_n475), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n368), .A2(new_n739), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n997), .A2(G97), .B1(new_n764), .B2(G303), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n751), .B2(new_n733), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n718), .B1(new_n1224), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n710), .B1(G68), .B2(new_n1115), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT124), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n928), .B2(new_n714), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1142), .B2(new_n709), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1217), .A2(new_n1239), .ZN(G381));
  OR2_X1    g1040(.A1(G375), .A2(KEYINPUT127), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1242), .A2(new_n1135), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G375), .A2(KEYINPUT127), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1241), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(G393), .A2(G396), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OR3_X1    g1048(.A1(new_n1245), .A2(G387), .A3(new_n1248), .ZN(G407));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G343), .C2(new_n1245), .ZN(G409));
  INV_X1    g1050(.A(G213), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1251), .A2(G343), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(G2897), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT60), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1215), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1215), .A2(new_n1255), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1256), .A2(new_n658), .A3(new_n1143), .A4(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1258), .A2(G384), .A3(new_n1239), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G384), .B1(new_n1258), .B2(new_n1239), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1254), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1239), .ZN(new_n1262));
  INV_X1    g1062(.A(G384), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1258), .A2(G384), .A3(new_n1239), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1265), .A3(new_n1253), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1261), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1188), .A2(G378), .A3(new_n1213), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1189), .A2(new_n1212), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1216), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1178), .A2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1243), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1269), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1252), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT61), .B1(new_n1268), .B2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(G390), .A2(new_n983), .A3(new_n1015), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n981), .B1(new_n966), .B2(new_n708), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1015), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1062), .B(new_n1085), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(G393), .B(new_n778), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1278), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT63), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1286), .B1(new_n1276), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1252), .B1(new_n1269), .B2(new_n1273), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1277), .A2(new_n1285), .A3(new_n1289), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1290), .A2(new_n1293), .A3(new_n1287), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1290), .B2(new_n1267), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1293), .B1(new_n1290), .B2(new_n1287), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1294), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1292), .B1(new_n1298), .B2(new_n1285), .ZN(G405));
  AND2_X1   g1099(.A1(G375), .A2(new_n1243), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1269), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1287), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1300), .A2(new_n1287), .A3(new_n1301), .ZN(new_n1304));
  OAI22_X1  g1104(.A1(new_n1303), .A2(new_n1304), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1304), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(new_n1285), .A3(new_n1302), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(G402));
endmodule


