//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n211), .A2(new_n212), .B1(new_n202), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G68), .B2(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n215), .B1(new_n203), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n210), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT0), .Z(new_n231));
  NOR2_X1   g0031(.A1(G58), .A2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n234), .A2(new_n208), .A3(new_n235), .ZN(new_n236));
  NOR3_X1   g0036(.A1(new_n228), .A2(new_n231), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n225), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n216), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G270), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G97), .B(G107), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(KEYINPUT70), .ZN(new_n253));
  OR2_X1    g0053(.A1(new_n253), .A2(KEYINPUT9), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(KEYINPUT9), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT67), .A2(G58), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT8), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(new_n208), .A3(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G150), .ZN(new_n260));
  OAI21_X1  g0060(.A(G20), .B1(new_n233), .B2(G50), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n235), .ZN(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n262), .A2(new_n264), .B1(new_n219), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n264), .B1(new_n207), .B2(G20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G50), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(new_n269), .B2(new_n272), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n254), .B(new_n255), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n275), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n277), .A2(new_n253), .A3(KEYINPUT9), .A4(new_n273), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n207), .B(G274), .C1(G41), .C2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n235), .B1(G33), .B2(G41), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT65), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n207), .B(KEYINPUT65), .C1(G41), .C2(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n281), .B1(new_n287), .B2(G226), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(G223), .B2(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G222), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(G1698), .ZN(new_n294));
  OR2_X1    g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(KEYINPUT3), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n294), .B1(G77), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(G1), .A3(G13), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT66), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n235), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(KEYINPUT66), .A3(new_n299), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n288), .B1(new_n298), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(G200), .B2(new_n306), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n279), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n279), .A2(new_n312), .A3(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n306), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n269), .A2(new_n272), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT68), .B(G179), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n316), .B(new_n317), .C1(new_n318), .C2(new_n306), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT16), .ZN(new_n321));
  INV_X1    g0121(.A(G68), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n295), .A2(new_n208), .A3(new_n296), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT7), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n291), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n224), .A2(new_n322), .ZN(new_n328));
  OAI21_X1  g0128(.A(G20), .B1(new_n328), .B2(new_n232), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n259), .A2(G159), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n321), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT7), .B1(new_n291), .B2(new_n208), .ZN(new_n333));
  NOR4_X1   g0133(.A1(new_n289), .A2(new_n290), .A3(new_n324), .A4(G20), .ZN(new_n334));
  OAI21_X1  g0134(.A(G68), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n331), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(KEYINPUT16), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n332), .A2(new_n337), .A3(new_n264), .ZN(new_n338));
  INV_X1    g0138(.A(new_n305), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n220), .A2(G1698), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n340), .B1(G223), .B2(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G87), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n281), .B1(new_n287), .B2(G232), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G200), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(new_n345), .A3(G190), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n257), .A2(new_n267), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n271), .B2(new_n257), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n338), .A2(new_n347), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT17), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n318), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n344), .A2(new_n345), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(G169), .B1(new_n344), .B2(new_n345), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n338), .A2(KEYINPUT72), .A3(new_n350), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT72), .B1(new_n338), .B2(new_n350), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT18), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(KEYINPUT18), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n353), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n322), .A2(G20), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n208), .A2(G33), .ZN(new_n366));
  INV_X1    g0166(.A(new_n259), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n365), .B1(new_n366), .B2(new_n221), .C1(new_n367), .C2(new_n219), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n264), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT11), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n271), .A2(G68), .ZN(new_n371));
  INV_X1    g0171(.A(new_n266), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n365), .ZN(new_n373));
  XOR2_X1   g0173(.A(new_n373), .B(KEYINPUT12), .Z(new_n374));
  NAND3_X1  g0174(.A1(new_n370), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT14), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n287), .A2(G238), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n280), .B(KEYINPUT71), .ZN(new_n379));
  INV_X1    g0179(.A(G1698), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n220), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n225), .A2(G1698), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n297), .B1(G33), .B2(G97), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n378), .B(new_n379), .C1(new_n305), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT13), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n297), .A2(new_n381), .A3(new_n382), .ZN(new_n387));
  INV_X1    g0187(.A(G33), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n387), .B1(new_n388), .B2(new_n202), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n339), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT13), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(new_n378), .A4(new_n379), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n377), .B1(new_n393), .B2(G169), .ZN(new_n394));
  AOI211_X1 g0194(.A(KEYINPUT14), .B(new_n315), .C1(new_n386), .C2(new_n392), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G179), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n376), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n376), .B1(new_n393), .B2(new_n307), .ZN(new_n402));
  INV_X1    g0202(.A(G200), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n386), .B2(new_n392), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n380), .A2(G232), .ZN(new_n406));
  INV_X1    g0206(.A(G238), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n297), .B(new_n406), .C1(new_n407), .C2(new_n380), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n339), .B(new_n408), .C1(G107), .C2(new_n297), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n287), .A2(G244), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n280), .A3(new_n410), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n411), .A2(G200), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n307), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT8), .B(G58), .Z(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n415));
  XOR2_X1   g0215(.A(KEYINPUT15), .B(G87), .Z(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n366), .B2(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(new_n264), .B1(new_n221), .B2(new_n268), .ZN(new_n419));
  INV_X1    g0219(.A(new_n271), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(new_n221), .B2(new_n420), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n412), .A2(new_n413), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n364), .A2(new_n401), .A3(new_n405), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n411), .A2(new_n315), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n409), .A2(new_n280), .A3(new_n354), .A4(new_n410), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n421), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n320), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G283), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n208), .C1(G33), .C2(new_n202), .ZN(new_n431));
  INV_X1    g0231(.A(G116), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G20), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n264), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT20), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT76), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n264), .A2(new_n433), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT76), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT20), .A4(new_n431), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n435), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n436), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n266), .A2(G20), .A3(new_n432), .ZN(new_n442));
  INV_X1    g0242(.A(new_n264), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n207), .A2(G33), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n443), .A2(new_n267), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G116), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n441), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT5), .B(G41), .ZN(new_n449));
  INV_X1    g0249(.A(G45), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(G1), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(G274), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n282), .B1(new_n451), .B2(new_n449), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n453), .B1(G270), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n380), .A2(G257), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n297), .B(new_n456), .C1(new_n216), .C2(new_n380), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n339), .B(new_n457), .C1(G303), .C2(new_n297), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G200), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n448), .B(new_n460), .C1(new_n307), .C2(new_n459), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n447), .A2(G169), .A3(new_n459), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT77), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(KEYINPUT21), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n464), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n447), .A2(new_n459), .A3(G169), .A4(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n459), .A2(new_n397), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n447), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT79), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n454), .A2(new_n471), .A3(G264), .ZN(new_n472));
  AND2_X1   g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  NOR2_X1   g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n451), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n300), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT79), .B1(new_n476), .B2(new_n216), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G294), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n297), .B1(G257), .B2(new_n380), .ZN(new_n480));
  NOR2_X1   g0280(.A1(G250), .A2(G1698), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n339), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n478), .A2(new_n483), .A3(G179), .A4(new_n452), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT81), .ZN(new_n485));
  OR2_X1    g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n485), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n478), .A2(new_n483), .A3(new_n452), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT80), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n488), .A2(new_n489), .A3(G169), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n488), .B2(G169), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n486), .B(new_n487), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n266), .A2(G20), .A3(new_n203), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n493), .B(KEYINPUT25), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT23), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(new_n203), .A3(G20), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT78), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT78), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n495), .A2(new_n497), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n208), .B(G87), .C1(new_n289), .C2(new_n290), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT22), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n297), .A2(new_n506), .A3(new_n208), .A4(G87), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n503), .A2(new_n508), .A3(KEYINPUT24), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT24), .B1(new_n503), .B2(new_n508), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n494), .B1(new_n511), .B2(new_n264), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n445), .A2(G107), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n470), .B1(new_n492), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n488), .A2(G200), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n478), .A2(new_n483), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(G190), .A3(new_n452), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n512), .A2(new_n513), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT4), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(G1698), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(G244), .C1(new_n290), .C2(new_n289), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n222), .B1(new_n295), .B2(new_n296), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(KEYINPUT4), .ZN(new_n524));
  OAI21_X1  g0324(.A(G250), .B1(new_n289), .B2(new_n290), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n380), .B1(new_n525), .B2(KEYINPUT4), .ZN(new_n526));
  INV_X1    g0326(.A(new_n430), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT73), .B1(new_n528), .B2(new_n305), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n453), .B1(G257), .B2(new_n454), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n212), .B1(new_n295), .B2(new_n296), .ZN(new_n531));
  OAI21_X1  g0331(.A(G1698), .B1(new_n531), .B2(new_n520), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n520), .B1(new_n291), .B2(new_n222), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n532), .A2(new_n430), .A3(new_n522), .A4(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT73), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n534), .A2(new_n535), .A3(new_n339), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n529), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G200), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n203), .A2(KEYINPUT6), .A3(G97), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n202), .A2(new_n203), .ZN(new_n540));
  NOR2_X1   g0340(.A1(G97), .A2(G107), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n539), .B1(new_n542), .B2(KEYINPUT6), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n544));
  OAI21_X1  g0344(.A(G107), .B1(new_n333), .B2(new_n334), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n443), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n445), .A2(G97), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n267), .A2(G97), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n534), .A2(new_n339), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n530), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G190), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n538), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G274), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n451), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n212), .B1(new_n450), .B2(G1), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n300), .A3(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n295), .A2(new_n296), .B1(new_n222), .B2(G1698), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n407), .A2(new_n380), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n559), .A2(new_n560), .B1(G33), .B2(G116), .ZN(new_n561));
  OAI211_X1 g0361(.A(G190), .B(new_n558), .C1(new_n561), .C2(new_n305), .ZN(new_n562));
  INV_X1    g0362(.A(new_n558), .ZN(new_n563));
  OAI221_X1 g0363(.A(new_n560), .B1(G244), .B2(new_n380), .C1(new_n289), .C2(new_n290), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n388), .B2(new_n432), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n563), .B1(new_n565), .B2(new_n339), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n562), .B1(new_n566), .B2(new_n403), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT19), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n366), .B2(new_n202), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n208), .B(G68), .C1(new_n289), .C2(new_n290), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n211), .A2(KEYINPUT74), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT74), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G87), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n204), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n575), .A2(new_n208), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n569), .B(new_n570), .C1(new_n574), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n264), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n417), .A2(new_n268), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n445), .A2(G87), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n567), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n566), .A2(G169), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n445), .A2(new_n416), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n578), .A2(new_n584), .A3(new_n579), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT75), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT75), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n578), .A2(new_n587), .A3(new_n584), .A4(new_n579), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n583), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n566), .A2(new_n354), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n582), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OR3_X1    g0391(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n551), .A2(new_n315), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n529), .A2(new_n530), .A3(new_n354), .A4(new_n536), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AND4_X1   g0395(.A1(new_n519), .A2(new_n554), .A3(new_n591), .A4(new_n595), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n429), .A2(new_n461), .A3(new_n515), .A4(new_n596), .ZN(G372));
  NOR2_X1   g0397(.A1(new_n402), .A2(new_n404), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n401), .B1(new_n598), .B2(new_n427), .ZN(new_n599));
  INV_X1    g0399(.A(new_n353), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n338), .A2(new_n350), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n357), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n361), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(KEYINPUT18), .A3(new_n357), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n314), .B1(new_n601), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n319), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n589), .A2(new_n590), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n519), .A2(new_n554), .A3(new_n591), .A4(new_n595), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n515), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT82), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n594), .A2(new_n614), .A3(new_n593), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n594), .B2(new_n593), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n591), .B(new_n592), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n617), .A2(KEYINPUT83), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT83), .B1(new_n617), .B2(new_n618), .ZN(new_n620));
  INV_X1    g0420(.A(new_n591), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n621), .A2(new_n618), .A3(new_n595), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n429), .B1(new_n613), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n610), .A2(new_n624), .ZN(G369));
  OR3_X1    g0425(.A1(new_n372), .A2(KEYINPUT27), .A3(G20), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT27), .B1(new_n372), .B2(G20), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(G213), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(G343), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n447), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n470), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n470), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n461), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G330), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n492), .A2(new_n514), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n519), .ZN(new_n638));
  INV_X1    g0438(.A(new_n630), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n512), .B2(new_n513), .ZN(new_n640));
  OAI22_X1  g0440(.A1(new_n638), .A2(new_n640), .B1(new_n637), .B2(new_n639), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n470), .A2(new_n639), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(new_n637), .A3(new_n519), .ZN(new_n645));
  INV_X1    g0445(.A(new_n637), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n639), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT84), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT84), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n645), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n642), .B1(new_n650), .B2(new_n653), .ZN(G399));
  INV_X1    g0454(.A(new_n229), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G41), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G1), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n574), .A2(new_n432), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n658), .A2(new_n659), .B1(new_n234), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT86), .ZN(new_n661));
  XNOR2_X1  g0461(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n621), .A2(new_n595), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n618), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n617), .A2(KEYINPUT26), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI211_X1 g0467(.A(KEYINPUT29), .B(new_n639), .C1(new_n667), .C2(new_n613), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT88), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n617), .A2(new_n618), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT83), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n622), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n617), .A2(KEYINPUT83), .A3(new_n618), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n613), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n630), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n668), .B(new_n669), .C1(new_n677), .C2(KEYINPUT29), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n668), .A2(new_n669), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n596), .A2(new_n461), .A3(new_n515), .A4(new_n639), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT30), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n468), .A2(new_n552), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n517), .A2(new_n566), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n551), .A2(new_n459), .A3(new_n397), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(KEYINPUT30), .A3(new_n517), .A4(new_n566), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n566), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n318), .B1(new_n458), .B2(new_n455), .ZN(new_n690));
  AND4_X1   g0490(.A1(new_n488), .A2(new_n537), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n630), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n630), .B(new_n695), .C1(new_n688), .C2(new_n691), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n681), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n680), .B1(G330), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n663), .B1(new_n698), .B2(G1), .ZN(G364));
  NOR2_X1   g0499(.A1(new_n307), .A2(G200), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n397), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G20), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G97), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n397), .A2(G200), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT95), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G20), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G190), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n703), .B1(new_n708), .B2(new_n203), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n571), .A2(new_n573), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n706), .A2(new_n307), .ZN(new_n711));
  AOI211_X1 g0511(.A(new_n291), .B(new_n709), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n354), .A2(new_n208), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT93), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(KEYINPUT93), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(new_n700), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G58), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n713), .A2(G200), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n307), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n719), .A2(G190), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n219), .A2(new_n721), .B1(new_n723), .B2(new_n322), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G190), .A2(G200), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n714), .A2(new_n715), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n724), .B1(new_n727), .B2(G77), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(G20), .A3(new_n397), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT94), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G159), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT32), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n712), .A2(new_n718), .A3(new_n728), .A4(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n711), .ZN(new_n738));
  INV_X1    g0538(.A(G303), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n720), .A2(G326), .B1(G294), .B2(new_n702), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT96), .Z(new_n742));
  INV_X1    g0542(.A(new_n733), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n740), .B(new_n742), .C1(G329), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n727), .A2(G311), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n717), .A2(G322), .ZN(new_n746));
  XNOR2_X1  g0546(.A(KEYINPUT33), .B(G317), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n297), .B1(new_n722), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n744), .A2(new_n745), .A3(new_n746), .A4(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G283), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n708), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n737), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n235), .B1(G20), .B2(new_n315), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n634), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n655), .A2(new_n291), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G355), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n248), .A2(G45), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT91), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n655), .A2(new_n297), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G45), .B2(new_n234), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n760), .B1(G116), .B2(new_n229), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n757), .A2(new_n753), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT92), .Z(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n208), .A2(G13), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT89), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G45), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G1), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n657), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT90), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n754), .A2(new_n758), .A3(new_n769), .A4(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n636), .ZN(new_n778));
  INV_X1    g0578(.A(new_n776), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n634), .A2(new_n635), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n777), .A2(new_n781), .ZN(G396));
  NOR2_X1   g0582(.A1(new_n753), .A2(new_n755), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT102), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n427), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n421), .A2(new_n425), .A3(KEYINPUT102), .A4(new_n426), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n422), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n421), .A2(new_n630), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n788), .A2(new_n789), .B1(new_n428), .B2(new_n630), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n776), .B1(G77), .B2(new_n784), .C1(new_n791), .C2(new_n756), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n707), .A2(G87), .B1(new_n743), .B2(G311), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT98), .Z(new_n794));
  AOI211_X1 g0594(.A(new_n297), .B(new_n794), .C1(G107), .C2(new_n711), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n727), .A2(G116), .B1(G303), .B2(new_n720), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n750), .B2(new_n723), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT97), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n717), .A2(G294), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n795), .A2(new_n798), .A3(new_n703), .A4(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT99), .B(G143), .Z(new_n801));
  AOI22_X1  g0601(.A1(new_n717), .A2(new_n801), .B1(G150), .B2(new_n722), .ZN(new_n802));
  INV_X1    g0602(.A(G137), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n802), .B1(new_n803), .B2(new_n721), .C1(new_n734), .C2(new_n726), .ZN(new_n804));
  XOR2_X1   g0604(.A(KEYINPUT100), .B(KEYINPUT34), .Z(new_n805));
  XNOR2_X1  g0605(.A(new_n804), .B(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G132), .ZN(new_n807));
  INV_X1    g0607(.A(new_n702), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n733), .A2(new_n807), .B1(new_n224), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G50), .B2(new_n711), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n806), .A2(new_n297), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n708), .A2(new_n322), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n800), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT101), .Z(new_n814));
  AOI21_X1  g0614(.A(new_n792), .B1(new_n814), .B2(new_n753), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n639), .B(new_n788), .C1(new_n623), .C2(new_n613), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n677), .B2(new_n791), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n697), .A2(G330), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT103), .Z(new_n820));
  NOR2_X1   g0620(.A1(new_n817), .A2(new_n818), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n776), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n815), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G384));
  INV_X1    g0624(.A(KEYINPUT38), .ZN(new_n825));
  INV_X1    g0625(.A(new_n628), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n358), .B2(new_n359), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT37), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n351), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n360), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n351), .A2(KEYINPUT106), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n603), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n351), .A2(KEYINPUT106), .ZN(new_n834));
  OAI21_X1  g0634(.A(KEYINPUT107), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n351), .A2(KEYINPUT106), .B1(new_n602), .B2(new_n357), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n338), .A2(new_n350), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT106), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n837), .A2(new_n838), .A3(new_n347), .A4(new_n348), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT107), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n835), .A2(new_n841), .A3(new_n827), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n831), .B1(new_n842), .B2(KEYINPUT37), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n351), .A2(new_n352), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT108), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n351), .A2(new_n352), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n847), .A2(new_n606), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n353), .A2(KEYINPUT108), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n827), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n825), .B1(new_n843), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n602), .A2(new_n826), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n603), .A2(new_n852), .A3(new_n351), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n830), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(KEYINPUT38), .B(new_n855), .C1(new_n364), .C2(new_n852), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n681), .A2(new_n692), .A3(new_n695), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n376), .A2(KEYINPUT105), .A3(new_n639), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT105), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n375), .B2(new_n630), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n400), .B2(new_n598), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n859), .A2(new_n861), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n405), .B(new_n864), .C1(new_n865), .C2(new_n376), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n790), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n692), .A2(KEYINPUT31), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n858), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n857), .A2(KEYINPUT40), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT40), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n855), .B1(new_n364), .B2(new_n852), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n825), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n873), .A2(new_n856), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n858), .A2(new_n867), .A3(new_n868), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n858), .A2(new_n868), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n429), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n877), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(G330), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT109), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n680), .A2(new_n429), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n610), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n882), .B(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n786), .A2(new_n639), .A3(new_n787), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT104), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n816), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n874), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n863), .A2(new_n866), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n607), .A2(new_n628), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n401), .A2(new_n630), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n873), .A2(KEYINPUT39), .A3(new_n856), .ZN(new_n894));
  INV_X1    g0694(.A(new_n856), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n849), .A2(new_n606), .A3(new_n847), .ZN(new_n896));
  INV_X1    g0696(.A(new_n359), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n338), .A2(KEYINPUT72), .A3(new_n350), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n628), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n836), .A2(new_n839), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n899), .B1(new_n901), .B2(KEYINPUT107), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n828), .B1(new_n902), .B2(new_n841), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n900), .B1(new_n903), .B2(new_n831), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n895), .B1(new_n904), .B2(new_n825), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n893), .B(new_n894), .C1(new_n905), .C2(KEYINPUT39), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n891), .A2(new_n892), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n885), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n207), .B2(new_n771), .ZN(new_n909));
  OAI211_X1 g0709(.A(G20), .B(new_n303), .C1(new_n543), .C2(KEYINPUT35), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n432), .B(new_n910), .C1(KEYINPUT35), .C2(new_n543), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT36), .Z(new_n912));
  OAI21_X1  g0712(.A(G77), .B1(new_n224), .B2(new_n322), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n234), .A2(new_n913), .B1(G50), .B2(new_n322), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(G1), .A3(new_n265), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n909), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT110), .ZN(G367));
  INV_X1    g0717(.A(new_n763), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n768), .B1(new_n229), .B2(new_n417), .C1(new_n244), .C2(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n581), .A2(new_n630), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n589), .A2(new_n590), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n621), .B2(new_n920), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n779), .B1(new_n923), .B2(new_n757), .ZN(new_n924));
  AOI22_X1  g0724(.A1(G50), .A2(new_n727), .B1(new_n717), .B2(G150), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n925), .B1(new_n224), .B2(new_n738), .C1(new_n221), .C2(new_n708), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n720), .A2(new_n801), .B1(G68), .B2(new_n702), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n803), .B2(new_n733), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n926), .A2(new_n291), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n734), .B2(new_n723), .ZN(new_n930));
  AOI22_X1  g0730(.A1(G294), .A2(new_n722), .B1(new_n720), .B2(G311), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n707), .A2(G97), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n931), .B(new_n932), .C1(new_n750), .C2(new_n726), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n297), .B(new_n933), .C1(G107), .C2(new_n702), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n711), .A2(KEYINPUT46), .A3(G116), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n717), .A2(G303), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT46), .B1(new_n711), .B2(G116), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(G317), .B2(new_n743), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n930), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT47), .Z(new_n941));
  INV_X1    g0741(.A(new_n753), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n919), .B(new_n924), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT112), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n554), .B(new_n595), .C1(new_n549), .C2(new_n639), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n592), .B(new_n630), .C1(new_n615), .C2(new_n616), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(new_n645), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT42), .Z(new_n950));
  XNOR2_X1  g0750(.A(new_n947), .B(KEYINPUT111), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n646), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n630), .B1(new_n952), .B2(new_n595), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n944), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(new_n923), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT43), .B1(new_n950), .B2(new_n953), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n923), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT43), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n955), .B2(new_n957), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n951), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n642), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n961), .B(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n947), .B1(new_n650), .B2(new_n653), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT45), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n649), .A2(new_n652), .A3(new_n948), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT113), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n966), .A2(KEYINPUT45), .ZN(new_n971));
  XOR2_X1   g0771(.A(KEYINPUT113), .B(KEYINPUT44), .Z(new_n972));
  OR2_X1    g0772(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n967), .A2(new_n970), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(new_n642), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n641), .A2(new_n644), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT114), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT114), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(new_n645), .A3(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(new_n778), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n975), .A2(new_n698), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n698), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n656), .B(KEYINPUT41), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n773), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n943), .B1(new_n965), .B2(new_n985), .ZN(G387));
  OR2_X1    g0786(.A1(new_n981), .A2(new_n698), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n981), .A2(new_n698), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n987), .A2(new_n656), .A3(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n717), .A2(G317), .B1(G311), .B2(new_n722), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n720), .A2(G322), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(new_n739), .C2(new_n726), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT48), .ZN(new_n993));
  INV_X1    g0793(.A(G294), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n993), .B1(new_n750), .B2(new_n808), .C1(new_n994), .C2(new_n738), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT49), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n707), .A2(G116), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n743), .A2(G326), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n996), .A2(new_n291), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n808), .A2(new_n417), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n727), .B2(G68), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n722), .A2(new_n257), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(new_n734), .C2(new_n721), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n711), .A2(G77), .ZN(new_n1004));
  INV_X1    g0804(.A(G150), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n932), .B(new_n1004), .C1(new_n1005), .C2(new_n733), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1003), .A2(new_n291), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n219), .B2(new_n716), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n942), .B1(new_n999), .B2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n641), .A2(G20), .A3(new_n756), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n759), .A2(new_n659), .B1(new_n203), .B2(new_n655), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT115), .Z(new_n1012));
  AOI21_X1  g0812(.A(new_n918), .B1(new_n241), .B2(G45), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n414), .A2(new_n219), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(new_n659), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(G68), .A2(G77), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1016), .A2(new_n450), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1012), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n776), .B1(new_n1020), .B2(new_n767), .ZN(new_n1021));
  OR3_X1    g0821(.A1(new_n1009), .A2(new_n1010), .A3(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n989), .B(new_n1022), .C1(new_n774), .C2(new_n980), .ZN(G393));
  INV_X1    g0823(.A(new_n975), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n657), .B1(new_n1024), .B2(new_n988), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n768), .B1(new_n251), .B2(new_n918), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G97), .B2(new_n655), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n743), .A2(new_n801), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n708), .B2(new_n211), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n702), .A2(G77), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n723), .B2(new_n219), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(G68), .C2(new_n711), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n727), .A2(new_n414), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n734), .A2(new_n716), .B1(new_n721), .B2(new_n1005), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT51), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n291), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1032), .A2(new_n1033), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n717), .A2(G311), .B1(G317), .B2(new_n720), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT52), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n707), .A2(G107), .B1(new_n743), .B2(G322), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1041), .B(new_n291), .C1(new_n750), .C2(new_n738), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT116), .Z(new_n1043));
  AOI211_X1 g0843(.A(new_n1040), .B(new_n1043), .C1(G303), .C2(new_n722), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n432), .B2(new_n808), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n726), .A2(new_n994), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1038), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n779), .B(new_n1027), .C1(new_n1047), .C2(new_n753), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(KEYINPUT117), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(KEYINPUT117), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n962), .A2(new_n757), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1025), .A2(new_n982), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n975), .A2(new_n773), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(G390));
  NOR2_X1   g0855(.A1(new_n808), .A2(new_n734), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n711), .A2(G150), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT120), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT53), .ZN(new_n1059));
  XOR2_X1   g0859(.A(KEYINPUT54), .B(G143), .Z(new_n1060));
  AOI22_X1  g0860(.A1(G132), .A2(new_n717), .B1(new_n727), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n743), .A2(G125), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n708), .B2(new_n219), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n291), .B(new_n1063), .C1(G128), .C2(new_n720), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1059), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1056), .B(new_n1065), .C1(G137), .C2(new_n722), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n733), .A2(new_n994), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n432), .A2(new_n716), .B1(new_n723), .B2(new_n203), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(G97), .C2(new_n727), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1069), .B(new_n1030), .C1(new_n750), .C2(new_n721), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n291), .B1(new_n738), .B2(new_n211), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n1070), .A2(new_n812), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n753), .B1(new_n1066), .B2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1073), .B(new_n776), .C1(new_n257), .C2(new_n784), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n894), .B1(new_n905), .B2(KEYINPUT39), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n755), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n697), .A2(G330), .A3(new_n791), .A4(new_n890), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n893), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n639), .B(new_n788), .C1(new_n667), .C2(new_n613), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1080), .A2(new_n887), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n890), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n857), .B(new_n1079), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n893), .B1(new_n888), .B2(new_n890), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n894), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT39), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n857), .B2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1078), .B(new_n1083), .C1(new_n1084), .C2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1082), .B1(new_n1080), .B2(new_n887), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1089), .A2(new_n905), .A3(new_n893), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n887), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n677), .B2(new_n788), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1079), .B1(new_n1092), .B2(new_n1082), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1090), .B1(new_n1093), .B2(new_n1075), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n858), .A2(new_n867), .A3(G330), .A4(new_n868), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1088), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1076), .B1(new_n1097), .B2(new_n773), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n429), .A2(new_n878), .A3(G330), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n609), .B(new_n1099), .C1(new_n680), .C2(new_n429), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n858), .A2(G330), .A3(new_n791), .A4(new_n868), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n1082), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n1081), .A3(new_n1077), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n697), .A2(G330), .A3(new_n791), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n869), .A2(G330), .B1(new_n1104), .B2(new_n1082), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1105), .A2(KEYINPUT118), .A3(new_n1092), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT118), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1104), .A2(new_n1082), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n1095), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1107), .B1(new_n1109), .B2(new_n888), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1103), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1082), .B1(new_n816), .B2(new_n887), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1075), .B1(new_n1112), .B2(new_n893), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1113), .A2(new_n1078), .A3(new_n1083), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1096), .B1(new_n1113), .B2(new_n1083), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1100), .B(new_n1111), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n788), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n630), .B(new_n1117), .C1(new_n675), .C2(new_n676), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n890), .B1(new_n1118), .B2(new_n1091), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n857), .A2(new_n1086), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1119), .A2(new_n1079), .B1(new_n1120), .B2(new_n894), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1095), .B1(new_n1121), .B2(new_n1090), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1099), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n883), .A2(new_n610), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1103), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT118), .B1(new_n1105), .B2(new_n1092), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1109), .A2(new_n1107), .A3(new_n888), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1122), .B(new_n1088), .C1(new_n1124), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT119), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n656), .B(new_n1116), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1111), .A2(new_n1100), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT119), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1098), .B1(new_n1131), .B2(new_n1134), .ZN(G378));
  OAI21_X1  g0935(.A(new_n1100), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n891), .A2(new_n892), .A3(new_n906), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT122), .Z(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n314), .B2(new_n319), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n274), .A2(new_n275), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n314), .A2(new_n319), .A3(new_n1140), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n826), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n826), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1144), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n1141), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1149), .A2(new_n870), .A3(new_n876), .A4(G330), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n870), .A2(new_n876), .A3(G330), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1149), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1137), .A2(new_n1150), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1137), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1136), .A2(KEYINPUT57), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1124), .B1(new_n1097), .B2(new_n1111), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1153), .A2(new_n1150), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n907), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1154), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1159), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1158), .A2(new_n656), .A3(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n733), .A2(new_n750), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n727), .A2(new_n416), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G41), .B1(new_n702), .B2(G68), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n720), .A2(G116), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1167), .A2(new_n1004), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1166), .B(new_n1170), .C1(G97), .C2(new_n722), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n297), .B1(new_n707), .B2(G58), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n203), .C2(new_n716), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n219), .B1(new_n289), .B2(G41), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n727), .A2(G137), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n717), .A2(G128), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n720), .A2(G125), .B1(G150), .B2(new_n702), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n722), .A2(G132), .B1(new_n711), .B2(new_n1060), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT59), .ZN(new_n1183));
  AOI21_X1  g0983(.A(G33), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(G41), .B1(new_n743), .B2(G124), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n734), .C2(new_n708), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1176), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n753), .B1(new_n1175), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n779), .B1(new_n219), .B2(new_n783), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n1152), .C2(new_n756), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT123), .Z(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1157), .B2(new_n773), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1165), .A2(new_n1193), .ZN(G375));
  NOR2_X1   g0994(.A1(new_n1111), .A2(new_n1100), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(new_n984), .A3(new_n1133), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n773), .B(KEYINPUT124), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1082), .A2(new_n755), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n784), .A2(G68), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n727), .A2(G150), .B1(G50), .B2(new_n702), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n803), .B2(new_n716), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n224), .A2(new_n708), .B1(new_n738), .B2(new_n734), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1060), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n297), .B1(new_n723), .B2(new_n1204), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n743), .A2(G128), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n807), .C2(new_n721), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n717), .A2(G283), .B1(G116), .B2(new_n722), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n739), .B2(new_n733), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1000), .B(new_n1210), .C1(G107), .C2(new_n727), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n221), .B2(new_n708), .C1(new_n994), .C2(new_n721), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n291), .B1(new_n738), .B2(new_n202), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1208), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n779), .B(new_n1200), .C1(new_n1214), .C2(new_n753), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1111), .A2(new_n1198), .B1(new_n1199), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1197), .A2(new_n1216), .ZN(G381));
  INV_X1    g1017(.A(KEYINPUT125), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1134), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1132), .A2(KEYINPUT119), .A3(new_n1133), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1219), .A2(new_n1220), .A3(new_n656), .A4(new_n1116), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1218), .B1(new_n1221), .B2(new_n1098), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(G378), .A2(KEYINPUT125), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1224), .A2(new_n1193), .A3(new_n1165), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1225), .A2(new_n823), .A3(new_n1216), .A4(new_n1197), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n965), .A2(new_n985), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1227), .A2(new_n943), .A3(new_n1228), .ZN(new_n1229));
  OR4_X1    g1029(.A1(G396), .A2(new_n1226), .A3(G393), .A4(new_n1229), .ZN(G407));
  NAND2_X1  g1030(.A1(new_n1225), .A2(new_n629), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(G407), .A2(G213), .A3(new_n1231), .ZN(G409));
  NAND3_X1  g1032(.A1(new_n1165), .A2(G378), .A3(new_n1193), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT126), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1165), .A2(G378), .A3(KEYINPUT126), .A4(new_n1193), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1192), .B1(new_n1157), .B2(new_n1198), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1136), .A2(new_n984), .A3(new_n1157), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n629), .A2(G213), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n657), .B1(new_n1195), .B2(KEYINPUT60), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n1133), .C1(KEYINPUT60), .C2(new_n1195), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1216), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n823), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1246), .A2(new_n823), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1242), .A2(new_n1243), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT62), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1242), .A2(KEYINPUT62), .A3(new_n1243), .A4(new_n1250), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(KEYINPUT127), .A3(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n629), .A2(G213), .A3(G2897), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1250), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1249), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1247), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1256), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT61), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT127), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1251), .A2(new_n1265), .A3(new_n1252), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1255), .A2(new_n1264), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G387), .A2(G390), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1229), .A2(new_n1268), .ZN(new_n1269));
  XOR2_X1   g1069(.A(G393), .B(G396), .Z(new_n1270));
  XNOR2_X1  g1070(.A(new_n1269), .B(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1263), .A2(new_n1257), .A3(new_n1261), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT63), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1251), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1251), .A2(new_n1274), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1277), .A2(new_n1271), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1272), .A2(new_n1279), .ZN(G405));
  NAND2_X1  g1080(.A1(new_n1224), .A2(G375), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1271), .A2(new_n1237), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1270), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1269), .B(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1237), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1282), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1259), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1282), .A2(new_n1286), .A3(new_n1250), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(G402));
endmodule


