//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G141gat), .B(G148gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n203), .B(new_n205), .C1(new_n206), .C2(KEYINPUT2), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n208), .A2(G148gat), .ZN(new_n209));
  XOR2_X1   g008(.A(KEYINPUT81), .B(G148gat), .Z(new_n210));
  AOI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(G141gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n203), .B1(new_n205), .B2(KEYINPUT2), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n207), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT82), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT81), .B(G148gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n212), .B1(new_n218), .B2(new_n209), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(KEYINPUT82), .A3(new_n207), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222));
  XNOR2_X1  g021(.A(G197gat), .B(G204gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT22), .ZN(new_n224));
  INV_X1    g023(.A(G211gat), .ZN(new_n225));
  INV_X1    g024(.A(G218gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n222), .B1(new_n230), .B2(KEYINPUT29), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n202), .B1(new_n221), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n230), .B(KEYINPUT76), .Z(new_n234));
  XOR2_X1   g033(.A(KEYINPUT77), .B(KEYINPUT29), .Z(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT83), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(new_n214), .B2(KEYINPUT3), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n219), .A2(KEYINPUT83), .A3(new_n222), .A4(new_n207), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n236), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n234), .B1(new_n240), .B2(KEYINPUT87), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(KEYINPUT87), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n233), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n230), .ZN(new_n245));
  INV_X1    g044(.A(new_n214), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT3), .B1(new_n245), .B2(new_n235), .ZN(new_n247));
  OAI22_X1  g046(.A1(new_n240), .A2(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n202), .B(KEYINPUT86), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(G22gat), .B1(new_n244), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n234), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n240), .A2(KEYINPUT87), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n232), .B1(new_n255), .B2(new_n242), .ZN(new_n256));
  INV_X1    g055(.A(G22gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(new_n257), .A3(new_n250), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT88), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT89), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT88), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n252), .A2(new_n262), .A3(new_n258), .ZN(new_n263));
  XOR2_X1   g062(.A(G78gat), .B(G106gat), .Z(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT31), .B(G50gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT89), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n259), .A2(KEYINPUT88), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n261), .A2(new_n263), .A3(new_n266), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n263), .A2(new_n266), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n267), .B1(new_n259), .B2(KEYINPUT88), .ZN(new_n271));
  AOI211_X1 g070(.A(new_n262), .B(KEYINPUT89), .C1(new_n252), .C2(new_n258), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  INV_X1    g074(.A(G183gat), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT69), .B1(new_n276), .B2(KEYINPUT27), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT27), .B(G183gat), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n275), .B(new_n277), .C1(new_n278), .C2(KEYINPUT69), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(KEYINPUT28), .A3(new_n275), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n284));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT26), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n289), .A2(KEYINPUT70), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n287), .A2(new_n293), .A3(new_n288), .ZN(new_n294));
  AOI211_X1 g093(.A(new_n284), .B(new_n286), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(KEYINPUT70), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n291), .A2(new_n290), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT71), .B1(new_n298), .B2(new_n285), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n283), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G113gat), .ZN(new_n301));
  INV_X1    g100(.A(G120gat), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT1), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(new_n301), .B2(new_n302), .ZN(new_n304));
  XOR2_X1   g103(.A(G127gat), .B(G134gat), .Z(new_n305));
  AND2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT67), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n309), .A2(KEYINPUT67), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n276), .A2(new_n275), .ZN(new_n313));
  NAND3_X1  g112(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n311), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n318), .A2(new_n288), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n317), .A2(G169gat), .ZN(new_n320));
  INV_X1    g119(.A(G176gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(KEYINPUT25), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT68), .B1(new_n316), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT65), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n309), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n309), .A2(new_n326), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n327), .A2(new_n328), .A3(new_n315), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT66), .B(G176gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n320), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n318), .B(new_n288), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n325), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  OR2_X1    g132(.A1(new_n309), .A2(KEYINPUT67), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n334), .A2(new_n310), .A3(new_n313), .A4(new_n314), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n322), .A2(KEYINPUT25), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT68), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n319), .A4(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n324), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n300), .A2(new_n308), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT72), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n300), .A2(new_n339), .A3(new_n342), .A4(new_n308), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n300), .A2(new_n339), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n304), .B(new_n305), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n341), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g146(.A1(G227gat), .A2(G233gat), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT34), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT32), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT33), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n347), .A2(KEYINPUT73), .A3(new_n348), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT73), .B1(new_n347), .B2(new_n348), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G15gat), .B(G43gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n347), .A2(new_n348), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n347), .A2(KEYINPUT73), .A3(new_n348), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n352), .B1(new_n360), .B2(KEYINPUT33), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n356), .A2(new_n360), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n354), .B2(new_n355), .ZN(new_n369));
  INV_X1    g168(.A(new_n353), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(new_n363), .B2(new_n364), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n369), .B1(new_n371), .B2(new_n359), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n350), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n274), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT35), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n216), .A2(KEYINPUT3), .A3(new_n220), .ZN(new_n377));
  INV_X1    g176(.A(new_n238), .ZN(new_n378));
  INV_X1    g177(.A(new_n239), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n377), .B(new_n345), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n308), .A2(new_n219), .A3(new_n207), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n381), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n380), .B(new_n385), .C1(new_n382), .C2(new_n381), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT5), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n216), .A2(new_n220), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n381), .B1(new_n388), .B2(new_n308), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n389), .B2(new_n384), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n384), .A2(KEYINPUT5), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n382), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT85), .B1(new_n381), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT85), .ZN(new_n396));
  INV_X1    g195(.A(new_n394), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n246), .A2(new_n396), .A3(new_n308), .A4(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(KEYINPUT84), .A2(KEYINPUT4), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n395), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n395), .B2(new_n398), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n380), .B(new_n392), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n391), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT0), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G57gat), .ZN(new_n406));
  INV_X1    g205(.A(G85gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n391), .A2(new_n402), .A3(new_n408), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n403), .A2(KEYINPUT6), .A3(new_n409), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(G226gat), .A2(G233gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n344), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n300), .B2(new_n339), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n418), .B(new_n245), .C1(new_n417), .C2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n418), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n417), .B1(new_n344), .B2(new_n235), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n420), .B1(new_n423), .B2(new_n234), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT78), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(G64gat), .ZN(new_n427));
  INV_X1    g226(.A(G92gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT78), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n431), .B(new_n420), .C1(new_n423), .C2(new_n234), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n425), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n420), .B(new_n429), .C1(new_n423), .C2(new_n234), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT30), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT80), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n437), .B1(new_n434), .B2(new_n438), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n433), .B(new_n436), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n416), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n375), .A2(new_n376), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n441), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n415), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n372), .A2(KEYINPUT74), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT74), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n447), .B(new_n369), .C1(new_n371), .C2(new_n359), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n351), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n368), .ZN(new_n450));
  NOR4_X1   g249(.A1(new_n274), .A2(new_n445), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n443), .B1(new_n451), .B2(new_n376), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n442), .B1(new_n269), .B2(new_n273), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n380), .B1(new_n400), .B2(new_n401), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT39), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n384), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n395), .A2(new_n398), .ZN(new_n458));
  INV_X1    g257(.A(new_n399), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n395), .A2(new_n399), .A3(new_n398), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n383), .B1(new_n462), .B2(new_n380), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT39), .B1(new_n389), .B2(new_n384), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT90), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(KEYINPUT90), .B(KEYINPUT39), .C1(new_n389), .C2(new_n384), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n457), .B(new_n408), .C1(new_n463), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT91), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT40), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n469), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  AND4_X1   g273(.A1(new_n410), .A2(new_n441), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n274), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT37), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(new_n425), .B2(new_n432), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n424), .A2(new_n477), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n430), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT38), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n413), .A2(new_n414), .A3(new_n434), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n423), .A2(new_n234), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n419), .A2(new_n417), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n230), .B1(new_n421), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(KEYINPUT37), .A3(new_n486), .ZN(new_n487));
  AOI211_X1 g286(.A(KEYINPUT38), .B(new_n429), .C1(new_n479), .C2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT92), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n413), .A2(new_n414), .A3(new_n434), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n491), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n482), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n454), .B1(new_n476), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n368), .A2(KEYINPUT36), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT75), .B1(new_n449), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n448), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n356), .A2(new_n360), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n447), .B1(new_n499), .B2(new_n369), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n350), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT75), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n351), .B2(new_n367), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n374), .A2(new_n503), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n497), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n495), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n453), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT11), .ZN(new_n511));
  INV_X1    g310(.A(G169gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G197gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n515), .B(KEYINPUT12), .Z(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT97), .ZN(new_n518));
  INV_X1    g317(.A(G8gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT95), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT16), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(G1gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT96), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(G1gat), .B2(new_n521), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI221_X1 g326(.A(new_n523), .B1(new_n524), .B2(new_n519), .C1(G1gat), .C2(new_n521), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G29gat), .ZN(new_n530));
  INV_X1    g329(.A(G36gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT14), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(G29gat), .B2(G36gat), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n532), .B(new_n534), .C1(new_n530), .C2(new_n531), .ZN(new_n535));
  INV_X1    g334(.A(G50gat), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n536), .A2(G43gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT93), .B(G43gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n537), .B1(new_n538), .B2(G50gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT15), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(G43gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(KEYINPUT15), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n535), .A2(new_n543), .ZN(new_n546));
  OR3_X1    g345(.A1(new_n545), .A2(KEYINPUT94), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT94), .B1(new_n545), .B2(new_n546), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n518), .B1(new_n529), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n547), .A2(new_n548), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n527), .A2(new_n528), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(KEYINPUT97), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n547), .A2(new_n556), .A3(new_n548), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT17), .B1(new_n545), .B2(new_n546), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n529), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT18), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n551), .A2(new_n552), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(new_n550), .B2(new_n553), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n555), .B(KEYINPUT13), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OAI22_X1  g364(.A1(new_n560), .A2(new_n561), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n557), .A2(new_n558), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n550), .A2(new_n553), .B1(new_n567), .B2(new_n529), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT18), .B1(new_n568), .B2(new_n555), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n517), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n560), .A2(new_n561), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(KEYINPUT18), .A3(new_n555), .ZN(new_n572));
  INV_X1    g371(.A(new_n562), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n564), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n571), .A2(new_n572), .A3(new_n575), .A4(new_n516), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n509), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  OR2_X1    g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT9), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G57gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(KEYINPUT98), .A3(G64gat), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(new_n585), .B2(G64gat), .ZN(new_n587));
  INV_X1    g386(.A(G64gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n588), .A2(G57gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(KEYINPUT98), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n584), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n585), .A2(G64gat), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT9), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n582), .A2(new_n581), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n529), .B1(new_n580), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT99), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n580), .ZN(new_n599));
  XNOR2_X1  g398(.A(G127gat), .B(G155gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n598), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n604));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n603), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT7), .ZN(new_n612));
  NAND2_X1  g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  AOI22_X1  g412(.A1(KEYINPUT8), .A2(new_n613), .B1(new_n407), .B2(new_n428), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G99gat), .B(G106gat), .Z(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n567), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n617), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n551), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G190gat), .B(G218gat), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n624));
  AND2_X1   g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n623), .A2(new_n624), .B1(KEYINPUT41), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n623), .A2(new_n624), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n620), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(new_n620), .B2(new_n627), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n633));
  XNOR2_X1  g432(.A(G134gat), .B(G162gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n631), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n627), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n628), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n635), .B1(new_n639), .B2(new_n630), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n610), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n596), .B1(new_n619), .B2(new_n617), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n591), .A2(new_n595), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n612), .A2(new_n614), .ZN(new_n646));
  INV_X1    g445(.A(new_n616), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(new_n648), .A3(new_n618), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n644), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n621), .A2(KEYINPUT10), .A3(new_n645), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n644), .B2(new_n649), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G120gat), .B(G148gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G176gat), .ZN(new_n659));
  INV_X1    g458(.A(G204gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n655), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n654), .B(KEYINPUT101), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n653), .A2(KEYINPUT102), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT102), .B1(new_n653), .B2(new_n663), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n664), .A2(new_n665), .A3(new_n656), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n662), .B1(new_n666), .B2(new_n661), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT103), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n669), .B(new_n662), .C1(new_n666), .C2(new_n661), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n643), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n579), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n415), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n444), .ZN(new_n676));
  OR3_X1    g475(.A1(new_n676), .A2(KEYINPUT104), .A3(new_n519), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT104), .B1(new_n676), .B2(new_n519), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n676), .A2(new_n679), .A3(new_n680), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n677), .B(new_n678), .C1(new_n681), .C2(new_n682), .ZN(G1325gat));
  NAND2_X1  g482(.A1(new_n507), .A2(KEYINPUT105), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n497), .A2(new_n505), .A3(new_n685), .A4(new_n506), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G15gat), .B1(new_n673), .B2(new_n689), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n374), .A2(G15gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n673), .B2(new_n691), .ZN(G1326gat));
  AND2_X1   g491(.A1(new_n269), .A2(new_n273), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n673), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT43), .B(G22gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  INV_X1    g495(.A(new_n610), .ZN(new_n697));
  INV_X1    g496(.A(new_n671), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n642), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n579), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n530), .A3(new_n416), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n684), .A2(new_n495), .A3(new_n686), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n452), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n641), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI211_X1 g508(.A(KEYINPUT44), .B(new_n641), .C1(new_n453), .C2(new_n508), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n699), .A2(new_n578), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n712), .B2(new_n415), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n704), .A2(new_n713), .ZN(G1328gat));
  NOR3_X1   g513(.A1(new_n701), .A2(G36gat), .A3(new_n444), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT46), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n712), .A2(new_n717), .A3(new_n444), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n712), .B2(new_n444), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G36gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n716), .B1(new_n718), .B2(new_n720), .ZN(G1329gat));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722));
  INV_X1    g521(.A(new_n538), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n374), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n722), .B1(new_n702), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n687), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n723), .B1(new_n712), .B2(new_n726), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n725), .A2(KEYINPUT109), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT109), .B1(new_n725), .B2(new_n727), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n712), .A2(new_n689), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n730), .A2(new_n723), .B1(new_n702), .B2(new_n724), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n732));
  OAI22_X1  g531(.A1(new_n728), .A2(new_n729), .B1(new_n731), .B2(new_n732), .ZN(G1330gat));
  NAND3_X1  g532(.A1(new_n702), .A2(new_n536), .A3(new_n274), .ZN(new_n734));
  OAI21_X1  g533(.A(G50gat), .B1(new_n712), .B2(new_n693), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT48), .Z(G1331gat));
  NOR3_X1   g536(.A1(new_n643), .A2(new_n577), .A3(new_n698), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n706), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n415), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(new_n585), .ZN(G1332gat));
  NOR2_X1   g540(.A1(new_n739), .A2(new_n444), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT49), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(new_n588), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT49), .B(G64gat), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT110), .Z(G1333gat));
  INV_X1    g546(.A(G71gat), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n689), .A2(new_n739), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n748), .B1(new_n739), .B2(new_n374), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT50), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n751), .A2(new_n755), .A3(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1334gat));
  NOR2_X1   g556(.A1(new_n739), .A2(new_n693), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(G78gat), .Z(G1335gat));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n610), .A2(new_n577), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n707), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n642), .B1(new_n705), .B2(new_n452), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n764), .A2(KEYINPUT51), .A3(new_n761), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n698), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(new_n407), .A3(new_n416), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n610), .A2(new_n577), .A3(new_n698), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n710), .B(new_n768), .C1(KEYINPUT44), .C2(new_n764), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n415), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(G1336gat));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  OAI21_X1  g571(.A(G92gat), .B1(new_n769), .B2(new_n444), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n444), .A2(G92gat), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n766), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n774), .B1(new_n766), .B2(new_n775), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n772), .B(new_n773), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n444), .A2(new_n698), .A3(G92gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n764), .B2(new_n761), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n765), .B1(new_n782), .B2(KEYINPUT113), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  AOI211_X1 g583(.A(new_n784), .B(new_n781), .C1(new_n764), .C2(new_n761), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n780), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n773), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n779), .B1(new_n787), .B2(KEYINPUT52), .ZN(new_n788));
  AOI211_X1 g587(.A(KEYINPUT114), .B(new_n772), .C1(new_n786), .C2(new_n773), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n778), .B1(new_n788), .B2(new_n789), .ZN(G1337gat));
  INV_X1    g589(.A(G99gat), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n769), .A2(new_n791), .A3(new_n689), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n766), .A2(new_n368), .A3(new_n373), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(new_n791), .ZN(G1338gat));
  OR2_X1    g593(.A1(new_n769), .A2(new_n693), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G106gat), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n763), .A2(new_n765), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n693), .A2(new_n698), .A3(G106gat), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT53), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n783), .A2(new_n785), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n801), .A2(new_n798), .B1(new_n795), .B2(G106gat), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(G1339gat));
  NAND2_X1  g603(.A1(new_n672), .A2(new_n578), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n529), .A2(new_n518), .A3(new_n549), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT97), .B1(new_n551), .B2(new_n552), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n559), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n555), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n808), .A2(new_n809), .B1(new_n563), .B2(new_n565), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n810), .A2(KEYINPUT117), .A3(new_n515), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n573), .B(new_n565), .C1(new_n806), .C2(new_n807), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n568), .B2(new_n555), .ZN(new_n814));
  INV_X1    g613(.A(new_n515), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n576), .A3(new_n641), .ZN(new_n818));
  INV_X1    g617(.A(new_n662), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n664), .B2(new_n665), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n653), .A2(new_n663), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n653), .B2(new_n654), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n661), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n819), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n821), .A2(new_n824), .A3(KEYINPUT55), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n827), .A2(KEYINPUT116), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT116), .B1(new_n827), .B2(new_n828), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n818), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n817), .A2(KEYINPUT118), .A3(new_n576), .A4(new_n671), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n577), .B1(new_n829), .B2(new_n830), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT117), .B1(new_n810), .B2(new_n515), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n814), .A2(new_n812), .A3(new_n815), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n835), .A2(new_n671), .A3(new_n576), .A4(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n833), .A2(new_n834), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n832), .B1(new_n840), .B2(new_n642), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n805), .B1(new_n841), .B2(new_n610), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n416), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n441), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n375), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n845), .A2(new_n301), .A3(new_n578), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n693), .A2(new_n501), .A3(new_n368), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n577), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n846), .B1(new_n301), .B2(new_n851), .ZN(G1340gat));
  NOR3_X1   g651(.A1(new_n845), .A2(new_n302), .A3(new_n698), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n671), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n302), .B2(new_n854), .ZN(G1341gat));
  OAI21_X1  g654(.A(G127gat), .B1(new_n845), .B2(new_n697), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n697), .A2(G127gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n849), .B2(new_n857), .ZN(G1342gat));
  OR3_X1    g657(.A1(new_n849), .A2(G134gat), .A3(new_n642), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n859), .A2(KEYINPUT56), .ZN(new_n860));
  OAI21_X1  g659(.A(G134gat), .B1(new_n845), .B2(new_n642), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(KEYINPUT56), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(G1343gat));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n843), .B(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n693), .A2(new_n441), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n578), .A2(G141gat), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n865), .A2(new_n689), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n687), .A2(new_n415), .A3(new_n441), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n827), .A2(new_n828), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT120), .Z(new_n872));
  OAI21_X1  g671(.A(new_n837), .B1(new_n872), .B2(new_n578), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n642), .ZN(new_n874));
  INV_X1    g673(.A(new_n832), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n610), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n805), .ZN(new_n877));
  OAI211_X1 g676(.A(KEYINPUT57), .B(new_n274), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n842), .B2(new_n274), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI211_X1 g680(.A(KEYINPUT119), .B(KEYINPUT57), .C1(new_n842), .C2(new_n274), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n577), .B(new_n870), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT124), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G141gat), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n883), .A2(KEYINPUT124), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n868), .B(new_n869), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n883), .A2(G141gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n868), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n888), .B1(new_n890), .B2(KEYINPUT58), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT122), .B(new_n892), .C1(new_n889), .C2(new_n868), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n887), .B1(new_n891), .B2(new_n893), .ZN(G1344gat));
  AND3_X1   g693(.A1(new_n865), .A2(new_n689), .A3(new_n866), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n210), .A3(new_n671), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n870), .B1(new_n881), .B2(new_n882), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(new_n698), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n898), .A2(new_n899), .A3(new_n217), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n842), .A2(new_n274), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT125), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n901), .A2(new_n904), .A3(KEYINPUT57), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n874), .B1(new_n871), .B2(new_n818), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n877), .B1(new_n906), .B2(new_n697), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n693), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n903), .B(new_n905), .C1(KEYINPUT57), .C2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n671), .A3(new_n870), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n899), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n896), .B1(new_n900), .B2(new_n911), .ZN(G1345gat));
  NAND2_X1  g711(.A1(new_n610), .A2(G155gat), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n897), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT126), .B1(new_n895), .B2(new_n610), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(G155gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n895), .A2(KEYINPUT126), .A3(new_n610), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(G1346gat));
  INV_X1    g718(.A(G162gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n895), .A2(new_n920), .A3(new_n641), .ZN(new_n921));
  OAI21_X1  g720(.A(G162gat), .B1(new_n897), .B2(new_n642), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n444), .A2(new_n416), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n842), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(new_n848), .ZN(new_n926));
  AOI21_X1  g725(.A(G169gat), .B1(new_n926), .B2(new_n577), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n375), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n928), .A2(new_n512), .A3(new_n578), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n927), .A2(new_n929), .ZN(G1348gat));
  AOI21_X1  g729(.A(G176gat), .B1(new_n926), .B2(new_n671), .ZN(new_n931));
  INV_X1    g730(.A(new_n928), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n671), .A2(new_n330), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n926), .A2(new_n278), .A3(new_n610), .ZN(new_n935));
  OAI21_X1  g734(.A(G183gat), .B1(new_n928), .B2(new_n697), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n926), .A2(new_n275), .A3(new_n641), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT127), .Z(new_n940));
  OAI21_X1  g739(.A(G190gat), .B1(new_n928), .B2(new_n642), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1351gat));
  AND2_X1   g742(.A1(new_n689), .A2(new_n924), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n909), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(G197gat), .B1(new_n945), .B2(new_n578), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n944), .A2(new_n901), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n514), .A3(new_n577), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1352gat));
  NAND3_X1  g748(.A1(new_n947), .A2(new_n660), .A3(new_n671), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n909), .A2(new_n671), .A3(new_n944), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G204gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n947), .A2(new_n225), .A3(new_n610), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n909), .A2(new_n610), .A3(new_n944), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n957), .B2(G211gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1354gat));
  OAI21_X1  g759(.A(G218gat), .B1(new_n945), .B2(new_n642), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n947), .A2(new_n226), .A3(new_n641), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1355gat));
endmodule


