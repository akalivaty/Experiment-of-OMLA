//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G20), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n209), .B1(new_n212), .B2(new_n213), .C1(new_n220), .C2(KEYINPUT1), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0022(.A(G238), .B(G244), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(G232), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT2), .B(G226), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n226), .B(new_n229), .Z(G358));
  XOR2_X1   g0030(.A(G87), .B(G97), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G107), .B(G116), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G68), .B(G77), .Z(new_n235));
  XOR2_X1   g0035(.A(G50), .B(G58), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G351));
  INV_X1    g0038(.A(KEYINPUT66), .ZN(new_n239));
  AND2_X1   g0039(.A1(G33), .A2(G41), .ZN(new_n240));
  OAI21_X1  g0040(.A(new_n239), .B1(new_n240), .B2(new_n210), .ZN(new_n241));
  NAND2_X1  g0041(.A1(G33), .A2(G41), .ZN(new_n242));
  NAND4_X1  g0042(.A1(new_n242), .A2(KEYINPUT66), .A3(G1), .A4(G13), .ZN(new_n243));
  AND2_X1   g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g0044(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n244), .A2(G226), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G222), .A2(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G223), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n247), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n211), .A2(new_n242), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n251), .B(new_n253), .C1(G77), .C2(new_n247), .ZN(new_n254));
  INV_X1    g0054(.A(new_n245), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n241), .A2(new_n255), .A3(G274), .A4(new_n243), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n246), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G169), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n210), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n204), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n262), .A2(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G50), .A2(G58), .ZN(new_n268));
  INV_X1    g0068(.A(G68), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n204), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n261), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(new_n210), .A3(new_n260), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n203), .A2(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G50), .ZN(new_n278));
  INV_X1    g0078(.A(new_n272), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n274), .A2(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n271), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n259), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G179), .ZN(new_n283));
  INV_X1    g0083(.A(new_n257), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n281), .B(KEYINPUT9), .ZN(new_n286));
  XOR2_X1   g0086(.A(KEYINPUT68), .B(G200), .Z(new_n287));
  NAND2_X1  g0087(.A1(new_n257), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(G190), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT10), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT10), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n286), .A2(new_n292), .A3(new_n288), .A4(new_n289), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n285), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT69), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n247), .A2(G232), .A3(new_n249), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n247), .A2(G238), .A3(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G107), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n296), .B(new_n297), .C1(new_n298), .C2(new_n247), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n253), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n244), .A2(G244), .A3(new_n245), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(new_n256), .A3(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n302), .A2(G179), .ZN(new_n303));
  INV_X1    g0103(.A(G77), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n203), .B2(G20), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n274), .A2(new_n305), .B1(new_n304), .B2(new_n279), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT15), .B(G87), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n307), .A2(new_n263), .B1(new_n204), .B2(new_n304), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n262), .A2(new_n266), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n261), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n310), .A2(KEYINPUT67), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(KEYINPUT67), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n306), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n302), .A2(new_n258), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n303), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n299), .A2(new_n253), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n301), .A2(new_n256), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n287), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n300), .A2(G190), .A3(new_n256), .A4(new_n301), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n310), .B(KEYINPUT67), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .A4(new_n306), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n294), .A2(new_n295), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n295), .B1(new_n294), .B2(new_n322), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT79), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n262), .A2(new_n279), .ZN(new_n326));
  INV_X1    g0126(.A(G58), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT8), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT8), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G58), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n275), .ZN(new_n332));
  OAI211_X1 g0132(.A(KEYINPUT78), .B(new_n326), .C1(new_n332), .C2(new_n273), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n260), .A2(new_n210), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n335), .A2(new_n331), .A3(new_n272), .A4(new_n275), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT78), .B1(new_n336), .B2(new_n326), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n325), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n326), .B1(new_n332), .B2(new_n273), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT78), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(KEYINPUT79), .A3(new_n333), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G33), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT3), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G33), .ZN(new_n347));
  AOI21_X1  g0147(.A(G20), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(KEYINPUT7), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  AOI211_X1 g0150(.A(new_n350), .B(G20), .C1(new_n345), .C2(new_n347), .ZN(new_n351));
  OAI21_X1  g0151(.A(G68), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n327), .A2(new_n269), .ZN(new_n353));
  NOR2_X1   g0153(.A1(G58), .A2(G68), .ZN(new_n354));
  OAI21_X1  g0154(.A(G20), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n265), .A2(G159), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(KEYINPUT16), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT76), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n348), .B2(KEYINPUT7), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n346), .A2(KEYINPUT77), .A3(G33), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n345), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT77), .B1(new_n346), .B2(G33), .ZN(new_n364));
  OAI211_X1 g0164(.A(KEYINPUT7), .B(new_n204), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(KEYINPUT76), .B(new_n350), .C1(new_n247), .C2(G20), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n361), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n357), .B1(new_n367), .B2(G68), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n261), .B(new_n359), .C1(new_n368), .C2(KEYINPUT16), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n241), .A2(G232), .A3(new_n245), .A4(new_n243), .ZN(new_n370));
  INV_X1    g0170(.A(G87), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n344), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(G223), .A2(G1698), .ZN(new_n373));
  INV_X1    g0173(.A(G226), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(G1698), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n372), .B1(new_n375), .B2(new_n247), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n256), .B(new_n370), .C1(new_n376), .C2(new_n252), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT80), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n374), .A2(G1698), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(G223), .B2(G1698), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n345), .A2(new_n347), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n253), .B1(new_n383), .B2(new_n372), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n384), .A2(KEYINPUT80), .A3(new_n256), .A4(new_n370), .ZN(new_n385));
  AOI21_X1  g0185(.A(G200), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n377), .A2(G190), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n343), .B(new_n369), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT17), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n338), .A2(new_n342), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n367), .A2(G68), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n358), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n359), .A2(new_n261), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n387), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n379), .A2(new_n385), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(G200), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n400), .A3(KEYINPUT17), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT16), .B1(new_n392), .B2(new_n358), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n359), .A2(new_n261), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n342), .B(new_n338), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n377), .A2(G179), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n379), .A2(new_n385), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(new_n258), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n404), .A2(KEYINPUT18), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT18), .B1(new_n404), .B2(new_n407), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n390), .B(new_n401), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  NOR3_X1   g0210(.A1(new_n323), .A2(new_n324), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n266), .A2(new_n278), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n263), .A2(new_n304), .B1(new_n204), .B2(G68), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n261), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XOR2_X1   g0214(.A(new_n414), .B(KEYINPUT11), .Z(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(KEYINPUT74), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(KEYINPUT74), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT12), .B1(new_n272), .B2(G68), .ZN(new_n418));
  OR3_X1    g0218(.A1(new_n272), .A2(KEYINPUT12), .A3(G68), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n269), .B1(new_n203), .B2(G20), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n418), .A2(new_n419), .B1(new_n274), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n416), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n374), .A2(G1698), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(new_n345), .A3(new_n347), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT70), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G97), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n345), .A2(new_n347), .A3(G232), .A4(G1698), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n424), .A2(new_n345), .A3(new_n347), .A4(KEYINPUT70), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n427), .A2(new_n428), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT71), .B1(new_n431), .B2(new_n253), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(KEYINPUT71), .A3(new_n253), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT73), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT13), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n244), .A2(G238), .A3(new_n245), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n438), .A2(new_n256), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n435), .A2(new_n436), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n431), .A2(KEYINPUT71), .A3(new_n253), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n437), .B(new_n439), .C1(new_n441), .C2(new_n432), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT73), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n439), .B1(new_n441), .B2(new_n432), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT13), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G190), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n423), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(KEYINPUT72), .A3(new_n442), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT72), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n445), .A2(new_n450), .A3(KEYINPUT13), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n449), .A2(G200), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n449), .A2(G169), .A3(new_n451), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT14), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT14), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n449), .A2(new_n456), .A3(G169), .A4(new_n451), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n283), .B1(new_n445), .B2(KEYINPUT13), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(new_n440), .A3(new_n443), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT75), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n458), .A2(new_n440), .A3(new_n443), .A4(KEYINPUT75), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n455), .A2(new_n457), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n453), .B1(new_n463), .B2(new_n422), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n411), .A2(KEYINPUT81), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT81), .B1(new_n411), .B2(new_n464), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n247), .A2(G257), .A3(new_n249), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n382), .A2(G303), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n345), .A2(new_n347), .A3(G264), .A4(G1698), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n253), .ZN(new_n472));
  OR2_X1    g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  NAND2_X1  g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(new_n203), .A3(G45), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n244), .A2(G270), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G45), .ZN(new_n478));
  AOI211_X1 g0278(.A(G1), .B(new_n478), .C1(new_n473), .C2(new_n474), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n244), .A2(G274), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n472), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  OR2_X1    g0281(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(G169), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n472), .A2(new_n477), .A3(new_n480), .A4(G179), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  INV_X1    g0286(.A(G97), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n486), .B(new_n204), .C1(G33), .C2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G116), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G20), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n261), .A2(KEYINPUT84), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT84), .B1(new_n261), .B2(new_n490), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT20), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT85), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n493), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n491), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT85), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT20), .A4(new_n488), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n494), .A2(new_n495), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n496), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n272), .A2(G116), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n273), .B1(new_n203), .B2(G33), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(G116), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n485), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n247), .A2(G257), .A3(G1698), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n345), .A2(new_n347), .A3(G250), .A4(new_n249), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G294), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n253), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n244), .A2(G264), .A3(new_n476), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n480), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n258), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n476), .A2(new_n241), .A3(new_n243), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(G264), .B1(new_n511), .B2(new_n253), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(new_n283), .A3(new_n480), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n345), .A2(new_n347), .A3(new_n204), .A4(G87), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT22), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT22), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n247), .A2(new_n521), .A3(new_n204), .A4(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  OR3_X1    g0324(.A1(new_n524), .A2(KEYINPUT87), .A3(G20), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT87), .B1(new_n524), .B2(G20), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n204), .B2(G107), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n298), .A2(KEYINPUT23), .A3(G20), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n525), .A2(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT24), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT24), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n523), .A2(new_n533), .A3(new_n530), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n335), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n272), .A2(G107), .ZN(new_n536));
  XNOR2_X1  g0336(.A(new_n536), .B(KEYINPUT25), .ZN(new_n537));
  INV_X1    g0337(.A(new_n504), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n298), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n515), .B(new_n518), .C1(new_n535), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n481), .A2(G169), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n502), .B2(new_n505), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n507), .B(new_n540), .C1(new_n482), .C2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT19), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n204), .B1(new_n428), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n371), .A2(new_n487), .A3(new_n298), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n345), .A2(new_n347), .A3(new_n204), .A4(G68), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n544), .B1(new_n263), .B2(new_n487), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(new_n261), .B1(new_n279), .B2(new_n307), .ZN(new_n551));
  INV_X1    g0351(.A(new_n307), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n504), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  OR2_X1    g0354(.A1(G238), .A2(G1698), .ZN(new_n555));
  INV_X1    g0355(.A(G244), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G1698), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n345), .A2(new_n555), .A3(new_n347), .A4(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n252), .B1(new_n558), .B2(new_n524), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  OR3_X1    g0360(.A1(new_n478), .A2(G1), .A3(G274), .ZN(new_n561));
  INV_X1    g0361(.A(G250), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n478), .B2(G1), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n241), .A2(new_n561), .A3(new_n243), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n283), .A3(new_n564), .ZN(new_n565));
  AND4_X1   g0365(.A1(new_n241), .A2(new_n561), .A3(new_n243), .A4(new_n563), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n258), .B1(new_n566), .B2(new_n559), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n554), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n560), .A2(G190), .A3(new_n564), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n287), .B1(new_n566), .B2(new_n559), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n504), .A2(G87), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n551), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G200), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n517), .B2(new_n480), .ZN(new_n575));
  INV_X1    g0375(.A(G190), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n514), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n535), .A2(new_n539), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n573), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n272), .A2(G97), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n504), .B2(G97), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT6), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n583), .A2(new_n487), .A3(G107), .ZN(new_n584));
  XNOR2_X1  g0384(.A(G97), .B(G107), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n586), .A2(new_n204), .B1(new_n304), .B2(new_n266), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(G107), .B2(new_n367), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n582), .B1(new_n588), .B2(new_n335), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n345), .A2(new_n347), .A3(G250), .A4(G1698), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n486), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n556), .A2(G1698), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT4), .B1(new_n247), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n592), .A2(new_n345), .A3(new_n347), .A4(KEYINPUT4), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT82), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n247), .A2(KEYINPUT82), .A3(KEYINPUT4), .A4(new_n592), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n252), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n244), .A2(G257), .A3(new_n476), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n480), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n600), .A2(new_n602), .A3(new_n576), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n589), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n594), .A2(new_n599), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n253), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n601), .A2(new_n480), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT83), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT83), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n600), .B2(new_n602), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n610), .A3(G200), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n604), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n606), .A2(new_n607), .A3(new_n283), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n258), .B1(new_n600), .B2(new_n602), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n589), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n481), .A2(new_n576), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n481), .A2(G200), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n616), .A2(new_n502), .A3(new_n505), .A4(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n580), .A2(new_n612), .A3(new_n615), .A4(new_n618), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n467), .A2(new_n543), .A3(new_n619), .ZN(G372));
  INV_X1    g0420(.A(KEYINPUT88), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n408), .B2(new_n409), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT18), .ZN(new_n623));
  INV_X1    g0423(.A(new_n405), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n399), .B2(G169), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n623), .B1(new_n397), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n404), .A2(KEYINPUT18), .A3(new_n407), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(KEYINPUT88), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n453), .A2(new_n315), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n422), .B2(new_n463), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT17), .B1(new_n397), .B2(new_n400), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n387), .B1(new_n406), .B2(new_n574), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n404), .A2(new_n634), .A3(new_n389), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n630), .B1(new_n632), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n291), .A2(new_n293), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n285), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n613), .A2(new_n614), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n611), .A2(new_n604), .B1(new_n641), .B2(new_n589), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n543), .A3(new_n580), .ZN(new_n643));
  INV_X1    g0443(.A(new_n568), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n615), .B2(new_n573), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n568), .A2(new_n572), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n641), .A2(new_n647), .A3(KEYINPUT26), .A4(new_n589), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n640), .B1(new_n467), .B2(new_n650), .ZN(G369));
  OAI21_X1  g0451(.A(new_n507), .B1(new_n482), .B2(new_n542), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n506), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g0459(.A(new_n652), .B(new_n659), .Z(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n618), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n540), .A2(new_n658), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n578), .A2(new_n579), .ZN(new_n666));
  INV_X1    g0466(.A(new_n658), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n579), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n665), .B1(new_n668), .B2(new_n540), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n665), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n652), .A2(new_n667), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n207), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n546), .A2(G116), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n213), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n658), .B1(new_n643), .B2(new_n649), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT29), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT89), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n642), .B(new_n580), .C1(new_n543), .C2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n543), .A2(new_n685), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n649), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n688), .A2(new_n667), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n684), .B1(new_n689), .B2(new_n683), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n566), .A2(new_n559), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n512), .A3(new_n513), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n484), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n600), .A2(new_n602), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n695), .A2(KEYINPUT30), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT30), .B1(new_n695), .B2(new_n696), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n693), .A2(G179), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n481), .A3(new_n514), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n696), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n697), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n692), .B1(new_n702), .B2(new_n667), .ZN(new_n703));
  INV_X1    g0503(.A(new_n698), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n695), .A2(KEYINPUT30), .A3(new_n696), .ZN(new_n705));
  INV_X1    g0505(.A(new_n701), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n619), .A2(new_n543), .A3(new_n658), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G330), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n691), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n681), .B1(new_n714), .B2(G1), .ZN(G364));
  INV_X1    g0515(.A(G13), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G20), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n203), .B1(new_n717), .B2(G45), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n677), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n662), .A2(G330), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n664), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n661), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n210), .B1(G20), .B2(new_n258), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n204), .A2(new_n283), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G190), .A2(G200), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n247), .B1(new_n732), .B2(G311), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n204), .A2(G179), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n730), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n574), .A2(G190), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n737), .A2(new_n204), .A3(new_n283), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n736), .A2(G329), .B1(new_n738), .B2(G322), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n287), .A2(new_n734), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G190), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G283), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n733), .B(new_n739), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n740), .A2(new_n576), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n744), .B1(G303), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n729), .A2(new_n576), .A3(G200), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n747), .A2(KEYINPUT91), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(KEYINPUT91), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT33), .B(G317), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n729), .A2(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n576), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT93), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G326), .ZN(new_n758));
  OAI21_X1  g0558(.A(G20), .B1(new_n737), .B2(G179), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT92), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G294), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n746), .A2(new_n753), .A3(new_n758), .A4(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G159), .ZN(new_n767));
  OR3_X1    g0567(.A1(new_n735), .A2(KEYINPUT32), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(KEYINPUT32), .B1(new_n735), .B2(new_n767), .ZN(new_n769));
  INV_X1    g0569(.A(new_n755), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n768), .B(new_n769), .C1(new_n770), .C2(new_n278), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n751), .B2(G68), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n741), .A2(G107), .ZN(new_n773));
  INV_X1    g0573(.A(new_n738), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n247), .B1(new_n304), .B2(new_n731), .C1(new_n774), .C2(new_n327), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G87), .B2(new_n745), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n763), .A2(new_n487), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n772), .A2(new_n773), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n728), .B1(new_n766), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n725), .A2(new_n727), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n675), .A2(new_n382), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G355), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G116), .B2(new_n207), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT90), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n237), .A2(G45), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n675), .A2(new_n247), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(G45), .C2(new_n213), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n784), .A2(KEYINPUT90), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n785), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n719), .B(new_n780), .C1(new_n781), .C2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n722), .B1(new_n726), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  NAND2_X1  g0593(.A1(new_n313), .A2(new_n658), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n321), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n315), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n303), .A2(new_n313), .A3(new_n314), .A4(new_n667), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  OR3_X1    g0599(.A1(new_n799), .A2(new_n682), .A3(KEYINPUT96), .ZN(new_n800));
  OAI21_X1  g0600(.A(KEYINPUT96), .B1(new_n799), .B2(new_n682), .ZN(new_n801));
  INV_X1    g0601(.A(new_n798), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n682), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n712), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT97), .Z(new_n806));
  AOI21_X1  g0606(.A(new_n720), .B1(new_n804), .B2(new_n712), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G311), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n382), .B1(new_n735), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G294), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n774), .A2(new_n811), .B1(new_n731), .B2(new_n489), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n810), .B(new_n812), .C1(G303), .C2(new_n755), .ZN(new_n813));
  INV_X1    g0613(.A(new_n745), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n371), .B2(new_n742), .C1(new_n298), .C2(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n777), .B(new_n815), .C1(G283), .C2(new_n751), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT94), .ZN(new_n817));
  INV_X1    g0617(.A(G132), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n247), .B1(new_n735), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n742), .A2(new_n269), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n819), .B(new_n820), .C1(G50), .C2(new_n745), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n732), .A2(G159), .B1(new_n738), .B2(G143), .ZN(new_n822));
  INV_X1    g0622(.A(G137), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n822), .B1(new_n823), .B2(new_n770), .C1(new_n750), .C2(new_n264), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(KEYINPUT34), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n764), .A2(G58), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n821), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT34), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n828), .B1(new_n829), .B2(new_n824), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n727), .B1(new_n817), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n727), .A2(new_n723), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n719), .B1(new_n304), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n831), .B(new_n833), .C1(new_n724), .C2(new_n802), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n808), .A2(new_n834), .ZN(G384));
  INV_X1    g0635(.A(new_n586), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n489), .B(new_n212), .C1(new_n836), .C2(KEYINPUT35), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(KEYINPUT35), .B2(new_n836), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT36), .ZN(new_n839));
  OAI21_X1  g0639(.A(G77), .B1(new_n327), .B2(new_n269), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n840), .A2(new_n213), .B1(G50), .B2(new_n269), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n841), .A2(G1), .A3(new_n716), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT98), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n690), .B1(new_n465), .B2(new_n466), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n640), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT103), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n463), .A2(new_n422), .A3(new_n667), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT38), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n350), .B1(new_n247), .B2(G20), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n382), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n269), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n394), .B1(new_n852), .B2(new_n357), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n359), .A2(new_n853), .A3(new_n261), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n334), .A2(new_n337), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n656), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n407), .A2(new_n856), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n388), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT101), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n397), .A2(new_n400), .B1(new_n407), .B2(new_n856), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT101), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n404), .A2(new_n407), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n404), .A2(new_n857), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n388), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n863), .A2(new_n865), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n626), .A2(new_n627), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n858), .B1(new_n636), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n870), .B1(new_n872), .B2(KEYINPUT100), .ZN(new_n873));
  INV_X1    g0673(.A(new_n858), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n410), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT100), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n849), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT100), .B1(new_n410), .B2(new_n874), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n872), .A2(KEYINPUT100), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT38), .A4(new_n870), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n878), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT39), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n622), .A2(new_n636), .A3(new_n628), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT102), .ZN(new_n886));
  INV_X1    g0686(.A(new_n868), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n885), .B2(new_n887), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n868), .A2(new_n621), .A3(new_n388), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n869), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n868), .A2(new_n388), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(KEYINPUT88), .A3(KEYINPUT37), .A4(new_n867), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n888), .A2(new_n889), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n882), .B1(new_n896), .B2(KEYINPUT38), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n848), .B(new_n883), .C1(new_n884), .C2(new_n897), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n658), .B(new_n798), .C1(new_n643), .C2(new_n649), .ZN(new_n899));
  INV_X1    g0699(.A(new_n797), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT99), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT99), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n803), .A2(new_n902), .A3(new_n797), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n461), .A2(new_n457), .A3(new_n462), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n454), .A2(KEYINPUT14), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n422), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n453), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n422), .A2(new_n658), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n422), .B(new_n658), .C1(new_n463), .C2(new_n453), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n904), .A2(new_n912), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n873), .A2(new_n877), .A3(new_n849), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n869), .A2(new_n866), .ZN(new_n915));
  INV_X1    g0715(.A(new_n859), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n864), .B2(KEYINPUT101), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n861), .A2(new_n862), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n879), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n920), .B2(new_n881), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n914), .A2(new_n921), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n913), .A2(new_n922), .B1(new_n630), .B2(new_n857), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n898), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n847), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n802), .B1(new_n709), .B2(new_n710), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n910), .B2(new_n911), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n927), .A2(KEYINPUT40), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n927), .B1(new_n914), .B2(new_n921), .ZN(new_n929));
  XNOR2_X1  g0729(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n928), .A2(new_n897), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n467), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n932), .A3(new_n711), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(G330), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n932), .B2(new_n711), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n925), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n203), .B2(new_n717), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n925), .A2(new_n936), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n844), .B1(new_n938), .B2(new_n939), .ZN(G367));
  NAND2_X1  g0740(.A1(new_n787), .A2(new_n229), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n725), .B(new_n727), .C1(new_n675), .C2(new_n552), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n719), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n667), .B1(new_n551), .B2(new_n571), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n644), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n573), .B2(new_n944), .ZN(new_n946));
  INV_X1    g0746(.A(new_n725), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n757), .A2(G143), .B1(G159), .B2(new_n751), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n745), .A2(G58), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n731), .A2(new_n278), .B1(new_n735), .B2(new_n823), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n247), .B1(new_n774), .B2(new_n264), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n950), .B(new_n951), .C1(G77), .C2(new_n741), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n763), .A2(new_n269), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n948), .A2(new_n949), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n247), .B1(new_n736), .B2(G317), .ZN(new_n956));
  INV_X1    g0756(.A(G303), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n956), .B1(new_n957), .B2(new_n774), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n742), .A2(new_n487), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n958), .B(new_n959), .C1(G311), .C2(new_n757), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT109), .B1(new_n745), .B2(G116), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT46), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n960), .B(new_n962), .C1(new_n811), .C2(new_n750), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n763), .A2(new_n298), .B1(new_n743), .B2(new_n731), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT108), .Z(new_n965));
  OAI21_X1  g0765(.A(new_n955), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT47), .Z(new_n967));
  OAI221_X1 g0767(.A(new_n943), .B1(new_n946), .B2(new_n947), .C1(new_n967), .C2(new_n728), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT106), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n589), .A2(new_n658), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n642), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n641), .A2(new_n589), .A3(new_n658), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT105), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n615), .B1(new_n976), .B2(new_n540), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n977), .A2(new_n667), .ZN(new_n978));
  INV_X1    g0778(.A(new_n974), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n979), .A2(new_n673), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT42), .Z(new_n981));
  OAI21_X1  g0781(.A(new_n970), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n982), .B(new_n983), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n670), .A2(new_n976), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n718), .B(KEYINPUT107), .Z(new_n987));
  NAND2_X1  g0787(.A1(new_n673), .A2(new_n671), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n979), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT44), .Z(new_n990));
  NOR2_X1   g0790(.A1(new_n988), .A2(new_n979), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(new_n670), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n669), .B(new_n672), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n663), .B(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n714), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n676), .B(KEYINPUT41), .Z(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n987), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n968), .B1(new_n986), .B2(new_n1001), .ZN(G387));
  NOR2_X1   g0802(.A1(new_n997), .A2(new_n713), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n677), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n997), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n714), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n959), .B1(G77), .B2(new_n745), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n731), .A2(new_n269), .B1(new_n735), .B2(new_n264), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n247), .B1(new_n774), .B2(new_n278), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(G159), .C2(new_n755), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n751), .A2(new_n331), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n764), .A2(new_n552), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n247), .B1(new_n736), .B2(G326), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n814), .A2(new_n811), .B1(new_n763), .B2(new_n743), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n732), .A2(G303), .B1(new_n738), .B2(G317), .ZN(new_n1016));
  INV_X1    g0816(.A(G322), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1016), .B1(new_n750), .B2(new_n809), .C1(new_n756), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT48), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1015), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n1019), .B2(new_n1018), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT49), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1014), .B1(new_n489), .B2(new_n742), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1013), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n727), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n678), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n782), .A2(new_n1027), .B1(new_n298), .B2(new_n675), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n226), .A2(new_n478), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n331), .A2(new_n278), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT50), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n678), .B(new_n478), .C1(new_n269), .C2(new_n304), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n787), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1028), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n719), .B1(new_n1034), .B2(new_n781), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1026), .B(new_n1035), .C1(new_n669), .C2(new_n947), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n987), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1006), .B(new_n1036), .C1(new_n997), .C2(new_n1037), .ZN(G393));
  AOI21_X1  g0838(.A(new_n677), .B1(new_n994), .B2(new_n1003), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n1003), .B2(new_n994), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n976), .A2(new_n725), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n234), .A2(new_n787), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n781), .B1(new_n487), .B2(new_n207), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n720), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n755), .A2(G150), .B1(G159), .B2(new_n738), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1045), .A2(KEYINPUT51), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G50), .B2(new_n751), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n745), .A2(G68), .ZN(new_n1048));
  INV_X1    g0848(.A(G143), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n247), .B1(new_n735), .B2(new_n1049), .C1(new_n262), .C2(new_n731), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G87), .B2(new_n741), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n764), .A2(G77), .B1(KEYINPUT51), .B2(new_n1045), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1047), .A2(new_n1048), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n755), .A2(G317), .B1(G311), .B2(new_n738), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT52), .Z(new_n1055));
  NAND2_X1  g0855(.A1(new_n745), .A2(G283), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n382), .B1(new_n735), .B2(new_n1017), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G294), .B2(new_n732), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1055), .A2(new_n773), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n750), .A2(new_n957), .B1(new_n763), .B2(new_n489), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT110), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1053), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT111), .Z(new_n1063));
  AOI21_X1  g0863(.A(new_n1044), .B1(new_n1063), .B2(new_n727), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n994), .A2(new_n987), .B1(new_n1041), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1040), .A2(new_n1065), .ZN(G390));
  OAI211_X1 g0866(.A(G330), .B(new_n802), .C1(new_n709), .C2(new_n710), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n910), .B2(new_n911), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n848), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n904), .B2(new_n912), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n885), .A2(new_n887), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n895), .B1(new_n1071), .B2(KEYINPUT102), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT38), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n884), .B1(new_n1074), .B2(new_n914), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n878), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1070), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n688), .A2(new_n667), .A3(new_n796), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n797), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n912), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1080), .B(new_n848), .C1(new_n1074), .C2(new_n914), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1068), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1068), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n883), .B1(new_n897), .B2(new_n884), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1081), .C1(new_n1085), .C2(new_n1070), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1083), .A2(new_n1086), .A3(new_n987), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT113), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n910), .A2(new_n911), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1090), .A2(new_n1067), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n904), .B1(new_n1091), .B2(new_n1068), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n799), .B(G330), .C1(new_n710), .C2(new_n709), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1093), .A2(new_n910), .A3(new_n911), .ZN(new_n1094));
  NOR4_X1   g0894(.A1(new_n1094), .A2(new_n1068), .A3(KEYINPUT112), .A4(new_n1079), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT112), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1068), .A2(new_n1079), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1092), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(G330), .B(new_n711), .C1(new_n465), .C2(new_n466), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n640), .A2(new_n845), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1089), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1083), .A2(new_n1086), .A3(new_n1103), .A4(new_n1100), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n676), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n832), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n720), .B1(new_n331), .B2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT114), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n820), .B1(G87), .B2(new_n745), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n774), .A2(new_n489), .B1(new_n735), .B2(new_n811), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n247), .B(new_n1112), .C1(G97), .C2(new_n732), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1111), .B(new_n1113), .C1(new_n743), .C2(new_n770), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n750), .A2(new_n298), .B1(new_n763), .B2(new_n304), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n755), .A2(G128), .B1(G132), .B2(new_n738), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT115), .ZN(new_n1117));
  INV_X1    g0917(.A(G125), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n247), .B1(new_n735), .B2(new_n1118), .C1(new_n731), .C2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G50), .B2(new_n741), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1117), .B(new_n1121), .C1(new_n767), .C2(new_n763), .ZN(new_n1122));
  OR3_X1    g0922(.A1(new_n814), .A2(KEYINPUT53), .A3(new_n264), .ZN(new_n1123));
  OAI21_X1  g0923(.A(KEYINPUT53), .B1(new_n814), .B2(new_n264), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(new_n750), .C2(new_n823), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1114), .A2(new_n1115), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1110), .B1(new_n1126), .B2(new_n727), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1085), .B2(new_n724), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1088), .A2(new_n1107), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(G378));
  NAND2_X1  g0930(.A1(new_n281), .A2(new_n857), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n294), .B(new_n1131), .Z(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1132), .B(new_n1133), .Z(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n723), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n720), .B1(G50), .B2(new_n1108), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n732), .A2(G137), .B1(new_n738), .B2(G128), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n1118), .B2(new_n770), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1119), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n745), .B2(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(new_n818), .B2(new_n750), .C1(new_n264), .C2(new_n763), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n741), .A2(G159), .ZN(new_n1143));
  AOI211_X1 g0943(.A(G33), .B(G41), .C1(new_n736), .C2(G124), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n247), .A2(G41), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G283), .B2(new_n736), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n742), .B2(new_n327), .C1(new_n304), .C2(new_n814), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT116), .Z(new_n1150));
  AOI22_X1  g0950(.A1(new_n732), .A2(new_n552), .B1(new_n738), .B2(G107), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n489), .B2(new_n770), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1152), .B(new_n953), .C1(G97), .C2(new_n751), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1145), .A2(new_n1146), .B1(new_n1154), .B2(KEYINPUT58), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1147), .B(new_n278), .C1(G33), .C2(G41), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(KEYINPUT58), .C2(new_n1154), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1136), .B1(new_n1157), .B2(new_n727), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1135), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT118), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n929), .A2(new_n930), .ZN(new_n1162));
  OAI211_X1 g0962(.A(KEYINPUT40), .B(new_n927), .C1(new_n1074), .C2(new_n914), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(G330), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT117), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT117), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1162), .A2(new_n1163), .A3(new_n1166), .A4(G330), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1167), .A3(new_n1134), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1134), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(KEYINPUT117), .A3(new_n1169), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1168), .A2(new_n924), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n924), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1161), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n924), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1166), .B1(new_n931), .B2(G330), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1167), .A2(new_n1134), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1170), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1174), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1168), .A2(new_n924), .A3(new_n1170), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(KEYINPUT118), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1173), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1160), .B1(new_n1182), .B2(new_n987), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1106), .A2(new_n1103), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1179), .A2(KEYINPUT57), .A3(new_n1184), .A4(new_n1180), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n676), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT119), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT119), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1185), .A2(new_n1188), .A3(new_n676), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1184), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n1173), .B2(new_n1181), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1192), .A2(KEYINPUT57), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1183), .B1(new_n1190), .B2(new_n1193), .ZN(G375));
  OAI211_X1 g0994(.A(new_n1102), .B(new_n1092), .C1(new_n1095), .C2(new_n1099), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1104), .A2(new_n1000), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n720), .B1(G68), .B2(new_n1108), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n912), .A2(new_n724), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n382), .B1(new_n736), .B2(G128), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n823), .B2(new_n774), .C1(new_n264), .C2(new_n731), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n327), .A2(new_n742), .B1(new_n814), .B2(new_n767), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(G132), .C2(new_n755), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n278), .B2(new_n763), .C1(new_n750), .C2(new_n1119), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n382), .B1(new_n735), .B2(new_n957), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n774), .A2(new_n743), .B1(new_n731), .B2(new_n298), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(G294), .C2(new_n755), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G77), .A2(new_n741), .B1(new_n745), .B2(G97), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n751), .A2(G116), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1206), .A2(new_n1012), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1203), .A2(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(KEYINPUT120), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n728), .B1(new_n1210), .B2(KEYINPUT120), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1197), .B(new_n1198), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1100), .B2(new_n987), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1196), .A2(new_n1214), .ZN(G381));
  NAND2_X1  g1015(.A1(new_n1182), .A2(new_n987), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1159), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1192), .A2(KEYINPUT57), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1185), .A2(new_n1188), .A3(new_n676), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1188), .B1(new_n1185), .B2(new_n676), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1217), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1129), .ZN(new_n1223));
  INV_X1    g1023(.A(G390), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1224), .B(new_n968), .C1(new_n986), .C2(new_n1001), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(G393), .A2(G396), .ZN(new_n1226));
  INV_X1    g1026(.A(G384), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  OR4_X1    g1028(.A1(G381), .A2(new_n1223), .A3(new_n1225), .A4(new_n1228), .ZN(G407));
  OAI211_X1 g1029(.A(G407), .B(G213), .C1(G343), .C2(new_n1223), .ZN(G409));
  AND2_X1   g1030(.A1(G387), .A2(G390), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1225), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AND2_X1   g1033(.A1(G393), .A2(G396), .ZN(new_n1234));
  OR3_X1    g1034(.A1(new_n1234), .A2(new_n1226), .A3(KEYINPUT125), .ZN(new_n1235));
  OAI21_X1  g1035(.A(KEYINPUT125), .B1(new_n1234), .B2(new_n1226), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1235), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT62), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n657), .A2(G213), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1171), .A2(new_n1172), .A3(new_n1037), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT121), .B1(new_n1243), .B2(new_n1160), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1179), .A2(new_n987), .A3(new_n1180), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT121), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n1246), .A3(new_n1159), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1244), .A2(new_n1129), .A3(new_n1247), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n999), .B(new_n1191), .C1(new_n1173), .C2(new_n1181), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1242), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G378), .B2(G375), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1104), .A2(KEYINPUT60), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT122), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1195), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT60), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1195), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT122), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n677), .B1(new_n1257), .B2(KEYINPUT60), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1254), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(G384), .A3(new_n1214), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G384), .B1(new_n1260), .B2(new_n1214), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1241), .B1(new_n1251), .B2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1187), .B(new_n1189), .C1(KEYINPUT57), .C2(new_n1192), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1129), .B1(new_n1266), .B2(new_n1183), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1264), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(new_n1267), .A2(new_n1250), .A3(KEYINPUT62), .A4(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1265), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1242), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT123), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(G2897), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1274), .B(KEYINPUT124), .Z(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1264), .A2(new_n1273), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1260), .A2(new_n1214), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1227), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(new_n1261), .A3(new_n1273), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1275), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G375), .A2(G378), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1244), .A2(new_n1129), .A3(new_n1247), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1249), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1272), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1282), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1271), .B1(new_n1287), .B2(KEYINPUT61), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1240), .B1(new_n1270), .B2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1238), .A2(new_n1239), .A3(new_n1271), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1277), .B(new_n1281), .C1(new_n1267), .C2(new_n1250), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT61), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1286), .B(new_n1264), .C1(new_n1222), .C2(new_n1129), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1251), .A2(KEYINPUT63), .A3(new_n1264), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1293), .B1(new_n1298), .B2(new_n1240), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT127), .B1(new_n1289), .B2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT63), .B1(new_n1251), .B2(new_n1264), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1240), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1293), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1240), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1294), .A2(KEYINPUT62), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1251), .A2(new_n1241), .A3(new_n1264), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT126), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1307), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1305), .A2(new_n1306), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1300), .A2(new_n1313), .ZN(G405));
  NAND2_X1  g1114(.A1(new_n1223), .A2(new_n1283), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1315), .B(new_n1268), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1316), .B(new_n1307), .ZN(G402));
endmodule


