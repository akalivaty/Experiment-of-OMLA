//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(G58), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n204), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT64), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n209), .B(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XOR2_X1   g0036(.A(G50), .B(G58), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  OR2_X1    g0042(.A1(KEYINPUT3), .A2(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(KEYINPUT3), .A2(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G223), .A3(G1698), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G222), .ZN(new_n250));
  OAI221_X1 g0050(.A(new_n246), .B1(new_n247), .B2(new_n245), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n215), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT65), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(KEYINPUT65), .A2(G33), .A3(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n252), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n260), .A2(new_n261), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n265), .B1(G226), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n256), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n269), .A2(G190), .B1(new_n270), .B2(KEYINPUT10), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(G200), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n204), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G150), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n204), .A2(new_n277), .ZN(new_n278));
  OAI22_X1  g0078(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G50), .A2(G58), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n204), .B1(new_n280), .B2(new_n211), .ZN(new_n281));
  OR2_X1    g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n215), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT66), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT66), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(new_n286), .A3(new_n215), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G50), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n290), .A2(new_n204), .A3(G1), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n282), .A2(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n203), .A2(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G50), .ZN(new_n294));
  XOR2_X1   g0094(.A(new_n294), .B(KEYINPUT67), .Z(new_n295));
  INV_X1    g0095(.A(new_n291), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(new_n285), .A3(new_n287), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n299), .A2(KEYINPUT9), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(KEYINPUT9), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n273), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n270), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT15), .B(G87), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n277), .A2(G20), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n308), .A2(new_n309), .B1(G20), .B2(G77), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n278), .B2(new_n274), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n311), .A2(new_n284), .B1(new_n247), .B2(new_n291), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n291), .A2(new_n284), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(G77), .A3(new_n293), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT68), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n245), .A2(G238), .A3(G1698), .ZN(new_n317));
  INV_X1    g0117(.A(G107), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n317), .B1(new_n318), .B2(new_n245), .C1(new_n249), .C2(new_n228), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n255), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n265), .B1(G244), .B2(new_n266), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n316), .B1(new_n323), .B2(G190), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n323), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(new_n322), .B1(new_n312), .B2(new_n315), .ZN(new_n328));
  INV_X1    g0128(.A(G179), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n304), .B1(new_n273), .B2(new_n302), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n268), .A2(new_n327), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n334), .B(new_n299), .C1(G179), .C2(new_n268), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n306), .A2(new_n332), .A3(new_n333), .A4(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n274), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n293), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n297), .A2(new_n338), .B1(new_n296), .B2(new_n337), .ZN(new_n339));
  INV_X1    g0139(.A(new_n284), .ZN(new_n340));
  AND2_X1   g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  NOR2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT7), .B1(new_n343), .B2(new_n204), .ZN(new_n344));
  AND4_X1   g0144(.A1(KEYINPUT7), .A2(new_n243), .A3(new_n204), .A4(new_n244), .ZN(new_n345));
  OAI21_X1  g0145(.A(G68), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G159), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n278), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G58), .A2(G68), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT78), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT78), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(G58), .A3(G68), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n352), .A3(new_n212), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n348), .B1(new_n353), .B2(G20), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n346), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n340), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n354), .A2(KEYINPUT79), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT79), .ZN(new_n359));
  AOI211_X1 g0159(.A(new_n359), .B(new_n348), .C1(new_n353), .C2(G20), .ZN(new_n360));
  OAI211_X1 g0160(.A(KEYINPUT16), .B(new_n346), .C1(new_n358), .C2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n339), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT81), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n260), .A2(G232), .A3(new_n261), .ZN(new_n364));
  MUX2_X1   g0164(.A(G223), .B(G226), .S(G1698), .Z(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(new_n245), .B1(G33), .B2(G87), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n264), .B(new_n364), .C1(new_n366), .C2(new_n254), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n367), .A2(G200), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n362), .A2(new_n363), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT17), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT17), .A4(new_n371), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n357), .A2(new_n361), .ZN(new_n377));
  INV_X1    g0177(.A(new_n339), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n365), .A2(new_n245), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G87), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n265), .B1(new_n255), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT80), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n383), .A2(new_n384), .A3(new_n329), .A4(new_n364), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT80), .B1(new_n367), .B2(G179), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n367), .A2(new_n327), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n379), .A2(new_n389), .A3(KEYINPUT18), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n362), .B2(new_n388), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n336), .A2(new_n376), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n264), .A2(KEYINPUT71), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT71), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n260), .A2(new_n263), .A3(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n396), .A2(new_n398), .B1(new_n266), .B2(G238), .ZN(new_n399));
  OAI211_X1 g0199(.A(G232), .B(G1698), .C1(new_n341), .C2(new_n342), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT70), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT70), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n245), .A2(new_n402), .A3(G232), .A4(G1698), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G97), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n245), .A2(G226), .A3(new_n248), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n401), .A2(new_n403), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n255), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n399), .A2(new_n407), .ZN(new_n408));
  XOR2_X1   g0208(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n399), .A2(new_n407), .A3(new_n409), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(KEYINPUT73), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT73), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(new_n414), .A3(new_n410), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G200), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n309), .A2(G77), .B1(G20), .B2(new_n211), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n289), .B2(new_n278), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n288), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT11), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(KEYINPUT11), .A3(new_n288), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n291), .A2(new_n211), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT12), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n313), .A2(G68), .A3(new_n293), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n422), .A2(new_n423), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT74), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n408), .A2(KEYINPUT13), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n429), .A2(new_n412), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n428), .B1(new_n430), .B2(G190), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n417), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT76), .B(KEYINPUT14), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n416), .A2(KEYINPUT77), .A3(G169), .A4(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n413), .A2(G169), .A3(new_n415), .A4(new_n433), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT77), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n435), .A2(new_n436), .B1(new_n430), .B2(G179), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n413), .A2(G169), .A3(new_n415), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n438), .A2(KEYINPUT75), .A3(KEYINPUT14), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT75), .B1(new_n438), .B2(KEYINPUT14), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n434), .B(new_n437), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n432), .B1(new_n441), .B2(new_n428), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n395), .A2(new_n442), .ZN(new_n443));
  AND2_X1   g0243(.A1(KEYINPUT4), .A2(G244), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n248), .B(new_n444), .C1(new_n341), .C2(new_n342), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G283), .ZN(new_n446));
  INV_X1    g0246(.A(G244), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n447), .B1(new_n243), .B2(new_n244), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n445), .B(new_n446), .C1(new_n448), .C2(KEYINPUT4), .ZN(new_n449));
  OAI21_X1  g0249(.A(G250), .B1(new_n341), .B2(new_n342), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n248), .B1(new_n450), .B2(KEYINPUT4), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n255), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g0252(.A1(KEYINPUT65), .A2(G33), .A3(G41), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT65), .B1(G33), .B2(G41), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n453), .A2(new_n454), .A3(new_n215), .ZN(new_n455));
  INV_X1    g0255(.A(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G1), .ZN(new_n457));
  NOR2_X1   g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  AND2_X1   g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(G274), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT84), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n203), .A2(G45), .ZN(new_n462));
  OR2_X1    g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  NAND2_X1  g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT84), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n465), .A2(new_n260), .A3(new_n466), .A4(G274), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n455), .A2(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G257), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n452), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G169), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n452), .A2(new_n468), .A3(G179), .A4(new_n470), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT6), .ZN(new_n474));
  AND2_X1   g0274(.A1(G97), .A2(G107), .ZN(new_n475));
  NOR2_X1   g0275(.A1(G97), .A2(G107), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n318), .A2(KEYINPUT6), .A3(G97), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n204), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n278), .A2(new_n247), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT82), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT82), .ZN(new_n482));
  INV_X1    g0282(.A(new_n480), .ZN(new_n483));
  NAND2_X1  g0283(.A1(KEYINPUT6), .A2(G97), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G107), .ZN(new_n485));
  XNOR2_X1  g0285(.A(G97), .B(G107), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(new_n474), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n482), .B(new_n483), .C1(new_n487), .C2(new_n204), .ZN(new_n488));
  OAI21_X1  g0288(.A(G107), .B1(new_n344), .B2(new_n345), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n481), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n284), .ZN(new_n491));
  INV_X1    g0291(.A(G97), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n291), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n203), .A2(G33), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n296), .A2(new_n285), .A3(new_n287), .A4(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n495), .B2(new_n492), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n472), .A2(new_n473), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT83), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n491), .B2(new_n497), .ZN(new_n500));
  AOI211_X1 g0300(.A(KEYINPUT83), .B(new_n496), .C1(new_n490), .C2(new_n284), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n471), .A2(new_n369), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(G200), .B2(new_n471), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n498), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(G257), .B(G1698), .C1(new_n341), .C2(new_n342), .ZN(new_n506));
  OAI211_X1 g0306(.A(G250), .B(new_n248), .C1(new_n341), .C2(new_n342), .ZN(new_n507));
  INV_X1    g0307(.A(G294), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n506), .B(new_n507), .C1(new_n277), .C2(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n255), .A2(new_n509), .B1(new_n469), .B2(G264), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n329), .A3(new_n468), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n255), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n469), .A2(G264), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n461), .A2(new_n467), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n327), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT23), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n204), .B2(G107), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n318), .A2(KEYINPUT23), .A3(G20), .ZN(new_n519));
  INV_X1    g0319(.A(G116), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n277), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n518), .A2(new_n519), .B1(new_n521), .B2(new_n204), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT22), .ZN(new_n523));
  AOI21_X1  g0323(.A(G20), .B1(new_n243), .B2(new_n244), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(G87), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n204), .B(G87), .C1(new_n341), .C2(new_n342), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(KEYINPUT22), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n522), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT24), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n526), .A2(KEYINPUT22), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n245), .A2(new_n523), .A3(new_n204), .A4(G87), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT24), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(new_n533), .A3(new_n522), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n340), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n495), .A2(new_n318), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n291), .A2(new_n318), .ZN(new_n537));
  XNOR2_X1  g0337(.A(new_n537), .B(KEYINPUT25), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n511), .B(new_n516), .C1(new_n535), .C2(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n532), .A2(new_n533), .A3(new_n522), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n533), .B1(new_n532), .B2(new_n522), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n284), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AND4_X1   g0344(.A1(new_n369), .A2(new_n468), .A3(new_n513), .A4(new_n512), .ZN(new_n545));
  AOI21_X1  g0345(.A(G200), .B1(new_n510), .B2(new_n468), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n544), .B(new_n539), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n245), .A2(new_n204), .A3(G68), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT19), .ZN(new_n550));
  INV_X1    g0350(.A(G87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n476), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n404), .A2(new_n204), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n275), .A2(KEYINPUT19), .A3(new_n492), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n549), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n340), .B1(new_n556), .B2(KEYINPUT85), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT85), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n549), .B(new_n558), .C1(new_n554), .C2(new_n555), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n495), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n308), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n307), .A2(new_n291), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n521), .B1(new_n448), .B2(G1698), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n245), .A2(G238), .A3(new_n248), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n255), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n457), .A2(G250), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n262), .B2(new_n457), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n260), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n327), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n567), .A2(new_n255), .B1(new_n570), .B2(new_n260), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n329), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n564), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(G200), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n557), .A2(new_n559), .B1(new_n291), .B2(new_n307), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n561), .A2(G87), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(G190), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(G264), .B(G1698), .C1(new_n341), .C2(new_n342), .ZN(new_n583));
  INV_X1    g0383(.A(G257), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(G1698), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n341), .B2(new_n342), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n243), .A2(G303), .A3(new_n244), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n255), .ZN(new_n589));
  INV_X1    g0389(.A(new_n465), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(G270), .A3(new_n260), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(G200), .B1(new_n515), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n446), .B(new_n204), .C1(G33), .C2(new_n492), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n520), .A2(G20), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n284), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n594), .A2(KEYINPUT20), .A3(new_n284), .A4(new_n595), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n595), .A2(G1), .A3(new_n290), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n520), .B1(new_n203), .B2(G33), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n601), .B1(new_n313), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n468), .A2(G190), .A3(new_n591), .A4(new_n589), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n593), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n468), .A2(new_n591), .A3(new_n589), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(G179), .A3(new_n604), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n327), .B1(new_n600), .B2(new_n603), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT21), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n608), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n608), .B2(new_n611), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n607), .B(new_n610), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n548), .A2(new_n582), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n443), .A2(new_n505), .A3(new_n616), .ZN(G372));
  OR2_X1    g0417(.A1(new_n613), .A2(new_n614), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(new_n610), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n541), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n578), .A2(new_n579), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(G190), .B2(new_n574), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT86), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n568), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n567), .A2(KEYINPUT86), .A3(new_n255), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n570), .A2(KEYINPUT87), .A3(new_n260), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT87), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n571), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n624), .A2(new_n625), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G200), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n564), .A2(new_n575), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n327), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n622), .A2(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n620), .A2(new_n505), .A3(new_n547), .A4(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n468), .A2(new_n470), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n327), .B1(new_n635), .B2(new_n452), .ZN(new_n636));
  INV_X1    g0436(.A(new_n473), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n638), .B(KEYINPUT88), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  INV_X1    g0440(.A(new_n502), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n639), .A2(new_n633), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n631), .A2(new_n632), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n582), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n498), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n644), .B1(new_n646), .B2(KEYINPUT26), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n634), .A2(new_n642), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n443), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n306), .A2(new_n333), .ZN(new_n650));
  INV_X1    g0450(.A(new_n432), .ZN(new_n651));
  INV_X1    g0451(.A(new_n331), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n441), .A2(new_n428), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n376), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT89), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n393), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n390), .A2(KEYINPUT89), .A3(new_n392), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n650), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n649), .A2(new_n661), .A3(new_n335), .ZN(G369));
  NOR2_X1   g0462(.A1(new_n290), .A2(G1), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n204), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT27), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n665), .A2(KEYINPUT90), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT90), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n664), .B2(KEYINPUT27), .ZN(new_n669));
  OAI221_X1 g0469(.A(G213), .B1(KEYINPUT27), .B2(new_n664), .C1(new_n667), .C2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n604), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n673), .B(KEYINPUT91), .Z(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n619), .A3(new_n607), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n619), .B2(new_n674), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n541), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n672), .B1(new_n535), .B2(new_n540), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n547), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n541), .A2(new_n672), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n619), .A2(new_n672), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n682), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(G41), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n207), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n552), .A2(G116), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n213), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  INV_X1    g0495(.A(new_n672), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n648), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(KEYINPUT29), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n639), .A2(new_n641), .A3(new_n633), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT26), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n643), .A2(KEYINPUT93), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n645), .A2(new_n640), .A3(new_n498), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n643), .A2(KEYINPUT93), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n701), .A2(new_n705), .A3(new_n634), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n699), .B1(new_n706), .B2(new_n696), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n548), .A2(new_n615), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n505), .A3(new_n645), .A4(new_n696), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT92), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n616), .A2(KEYINPUT92), .A3(new_n505), .A4(new_n696), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n572), .A2(new_n608), .A3(new_n514), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n637), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n609), .A2(G179), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n510), .A2(new_n468), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(new_n629), .A3(new_n471), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n715), .A2(new_n637), .A3(KEYINPUT30), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n718), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT31), .B1(new_n723), .B2(new_n672), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n708), .B1(new_n714), .B2(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n698), .A2(new_n707), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n695), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n290), .A2(G20), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT94), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G45), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G1), .ZN(new_n733));
  INV_X1    g0533(.A(new_n691), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n677), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G330), .B2(new_n676), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n207), .A2(new_n245), .ZN(new_n738));
  INV_X1    g0538(.A(G355), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n738), .A2(new_n739), .B1(G116), .B2(new_n207), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n238), .A2(G45), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n207), .A2(new_n343), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n456), .B2(new_n214), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n740), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n215), .B1(G20), .B2(new_n327), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n735), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n204), .A2(new_n329), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n369), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n204), .A2(G190), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G179), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n347), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n755), .A2(new_n289), .B1(new_n760), .B2(KEYINPUT32), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n204), .B1(new_n757), .B2(G190), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n492), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n325), .A2(G179), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n756), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n318), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n765), .A2(G20), .A3(G190), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n343), .B(new_n767), .C1(G87), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n753), .A2(G190), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n760), .A2(KEYINPUT32), .B1(new_n771), .B2(G68), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n764), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n752), .ZN(new_n774));
  AOI21_X1  g0574(.A(G200), .B1(new_n774), .B2(KEYINPUT95), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(KEYINPUT95), .B2(new_n774), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n369), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n776), .A2(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n210), .A2(new_n778), .B1(new_n780), .B2(new_n247), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  INV_X1    g0582(.A(G322), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n780), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT33), .B(G317), .ZN(new_n785));
  INV_X1    g0585(.A(new_n762), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n771), .A2(new_n785), .B1(G294), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n758), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n769), .A2(G303), .B1(new_n788), .B2(G329), .ZN(new_n789));
  INV_X1    g0589(.A(new_n766), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n245), .B1(new_n790), .B2(G283), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n754), .A2(G326), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n787), .A2(new_n789), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n773), .A2(new_n781), .B1(new_n784), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n751), .B1(new_n794), .B2(new_n748), .ZN(new_n795));
  INV_X1    g0595(.A(new_n747), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n676), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n737), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(G396));
  NAND2_X1  g0599(.A1(new_n316), .A2(new_n672), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n326), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n331), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n652), .A2(new_n696), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n697), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n804), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n648), .A2(new_n696), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n727), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n735), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n805), .A2(new_n727), .A3(new_n807), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n748), .A2(new_n745), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n735), .B1(G77), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G303), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n755), .A2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n763), .B(new_n816), .C1(G283), .C2(new_n771), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n768), .A2(new_n318), .B1(new_n758), .B2(new_n782), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n245), .B(new_n818), .C1(G87), .C2(new_n790), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G116), .A2(new_n779), .B1(new_n777), .B2(G294), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n768), .A2(new_n289), .B1(new_n766), .B2(new_n211), .ZN(new_n822));
  INV_X1    g0622(.A(G132), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n245), .B1(new_n758), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT96), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n822), .B(new_n825), .C1(G58), .C2(new_n786), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT97), .Z(new_n827));
  AOI22_X1  g0627(.A1(G137), .A2(new_n754), .B1(new_n771), .B2(G150), .ZN(new_n828));
  INV_X1    g0628(.A(G143), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n778), .B2(new_n829), .C1(new_n347), .C2(new_n780), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT34), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n830), .A2(new_n831), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n821), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n814), .B1(new_n835), .B2(new_n748), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n746), .B2(new_n806), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n811), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G384));
  NOR2_X1   g0639(.A1(new_n731), .A2(new_n203), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n346), .B1(new_n358), .B2(new_n360), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n356), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(new_n288), .A3(new_n361), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n378), .ZN(new_n844));
  INV_X1    g0644(.A(new_n670), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n394), .B2(new_n376), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n389), .A2(new_n379), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n379), .A2(new_n845), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n362), .A2(new_n371), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n844), .A2(new_n389), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n846), .A2(new_n855), .A3(KEYINPUT37), .A4(new_n851), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n848), .A2(KEYINPUT38), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n851), .B(new_n656), .C1(new_n362), .C2(new_n670), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n852), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n362), .A2(new_n670), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n362), .B2(new_n371), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n862), .A2(KEYINPUT89), .A3(KEYINPUT37), .A4(new_n849), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n374), .A2(new_n375), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n657), .A2(new_n865), .A3(new_n658), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n864), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n857), .B1(new_n867), .B2(KEYINPUT38), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n654), .A2(new_n672), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n846), .B1(new_n865), .B2(new_n393), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n854), .A2(new_n856), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n857), .A3(KEYINPUT39), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n870), .A2(new_n871), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n660), .A2(new_n670), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n807), .A2(new_n803), .ZN(new_n880));
  INV_X1    g0680(.A(new_n428), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n437), .A2(new_n434), .ZN(new_n882));
  INV_X1    g0682(.A(new_n440), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n438), .A2(KEYINPUT75), .A3(KEYINPUT14), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n881), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n672), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n881), .A2(new_n696), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n654), .A2(new_n651), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n880), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT100), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n807), .A2(new_n803), .B1(new_n887), .B2(new_n890), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT100), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n875), .A2(new_n857), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n879), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n443), .B1(new_n698), .B2(new_n707), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(new_n335), .A3(new_n661), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n899), .B(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n804), .B1(new_n714), .B2(new_n726), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n888), .B(new_n432), .C1(new_n441), .C2(new_n428), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n654), .A2(new_n696), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n903), .B(new_n897), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT40), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n868), .A2(new_n891), .A3(KEYINPUT40), .A4(new_n903), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n714), .A2(new_n726), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n443), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n708), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n910), .B2(new_n912), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n840), .B1(new_n902), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n902), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n214), .A2(G77), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n350), .A2(new_n352), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n917), .A2(new_n918), .B1(G50), .B2(new_n211), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(G1), .A3(new_n290), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT98), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT36), .ZN(new_n922));
  INV_X1    g0722(.A(new_n487), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n923), .A2(KEYINPUT35), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(KEYINPUT35), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n924), .A2(new_n925), .A3(G116), .A4(new_n216), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n921), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n922), .B2(new_n926), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT99), .Z(new_n929));
  NAND2_X1  g0729(.A1(new_n916), .A2(new_n929), .ZN(G367));
  OAI221_X1 g0730(.A(new_n749), .B1(new_n207), .B2(new_n307), .C1(new_n234), .C2(new_n742), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n735), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n762), .A2(new_n211), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n755), .A2(new_n829), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n933), .B(new_n934), .C1(G159), .C2(new_n771), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n768), .A2(new_n210), .B1(new_n766), .B2(new_n247), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n343), .B(new_n936), .C1(G137), .C2(new_n788), .ZN(new_n937));
  AOI22_X1  g0737(.A1(G50), .A2(new_n779), .B1(new_n777), .B2(G150), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT107), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n768), .A2(new_n520), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(KEYINPUT46), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT104), .Z(new_n943));
  AOI22_X1  g0743(.A1(KEYINPUT46), .A2(new_n941), .B1(new_n771), .B2(G294), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT105), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT105), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n777), .A2(G303), .ZN(new_n948));
  XNOR2_X1  g0748(.A(KEYINPUT106), .B(G317), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n343), .B1(new_n758), .B2(new_n949), .C1(new_n492), .C2(new_n766), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n755), .A2(new_n782), .B1(new_n762), .B2(new_n318), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n950), .B(new_n951), .C1(G283), .C2(new_n779), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n946), .A2(new_n947), .A3(new_n948), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n940), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT47), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n932), .B1(new_n955), .B2(new_n748), .ZN(new_n956));
  INV_X1    g0756(.A(new_n633), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n621), .A2(new_n672), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT101), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n644), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(new_n747), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n956), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n639), .A2(new_n641), .A3(new_n672), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n505), .B1(new_n502), .B2(new_n696), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n687), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT42), .Z(new_n968));
  INV_X1    g0768(.A(new_n966), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(new_n541), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n696), .B1(new_n970), .B2(new_n498), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n960), .A2(new_n961), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n975), .B(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n685), .A2(new_n969), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT102), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n978), .A2(KEYINPUT102), .A3(new_n979), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(new_n979), .C2(new_n978), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n688), .A2(new_n966), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT45), .Z(new_n986));
  NOR2_X1   g0786(.A1(new_n688), .A2(new_n966), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT44), .ZN(new_n988));
  AND3_X1   g0788(.A1(new_n986), .A2(new_n685), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n685), .B1(new_n986), .B2(new_n988), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n683), .B(new_n686), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT103), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(new_n678), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n677), .B(KEYINPUT103), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n995), .B1(new_n996), .B2(new_n993), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n728), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n728), .B1(new_n992), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n691), .B(KEYINPUT41), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n733), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n963), .B1(new_n984), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT108), .ZN(G387));
  INV_X1    g0804(.A(new_n998), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(new_n691), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n728), .B2(new_n997), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n683), .A2(new_n747), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n738), .A2(new_n692), .B1(G107), .B2(new_n207), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n231), .A2(new_n456), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT109), .Z(new_n1011));
  INV_X1    g0811(.A(new_n692), .ZN(new_n1012));
  AOI211_X1 g0812(.A(G45), .B(new_n1012), .C1(G68), .C2(G77), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n274), .A2(G50), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT50), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n742), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1009), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n735), .B1(new_n1017), .B2(new_n750), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G311), .A2(new_n771), .B1(new_n754), .B2(G322), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n778), .B2(new_n949), .C1(new_n815), .C2(new_n780), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT48), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n769), .A2(G294), .B1(new_n786), .B2(G283), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT49), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n766), .A2(new_n520), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n245), .B(new_n1029), .C1(G326), .C2(new_n788), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n786), .A2(new_n308), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n771), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1032), .B1(new_n755), .B2(new_n347), .C1(new_n274), .C2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n245), .B1(new_n766), .B2(new_n492), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n768), .A2(new_n247), .B1(new_n758), .B2(new_n276), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n289), .B2(new_n778), .C1(new_n211), .C2(new_n780), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1031), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1018), .B1(new_n1039), .B2(new_n748), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n997), .A2(new_n733), .B1(new_n1008), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1007), .A2(new_n1041), .ZN(G393));
  NAND2_X1  g0842(.A1(new_n969), .A2(new_n747), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT110), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n777), .A2(G159), .B1(G150), .B2(new_n754), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT51), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n780), .A2(new_n274), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n769), .A2(G68), .B1(new_n788), .B2(G143), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n245), .C1(new_n551), .C2(new_n766), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1033), .A2(new_n289), .B1(new_n762), .B2(new_n247), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT111), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(KEYINPUT111), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n777), .A2(G311), .B1(G317), .B2(new_n754), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT52), .Z(new_n1055));
  OAI22_X1  g0855(.A1(new_n1033), .A2(new_n815), .B1(new_n762), .B2(new_n520), .ZN(new_n1056));
  INV_X1    g0856(.A(G283), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n768), .A2(new_n1057), .B1(new_n758), .B2(new_n783), .ZN(new_n1058));
  NOR4_X1   g0858(.A1(new_n1056), .A2(new_n1058), .A3(new_n245), .A4(new_n767), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1055), .B(new_n1059), .C1(new_n508), .C2(new_n780), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1052), .A2(new_n1053), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n748), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n749), .B1(new_n492), .B2(new_n207), .C1(new_n241), .C2(new_n742), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1044), .A2(new_n735), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n733), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n734), .B1(new_n992), .B2(new_n998), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n991), .A2(new_n1005), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1064), .B1(new_n1065), .B2(new_n992), .C1(new_n1066), .C2(new_n1067), .ZN(G390));
  OAI21_X1  g0868(.A(new_n735), .B1(new_n337), .B2(new_n813), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n762), .A2(new_n247), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n755), .A2(new_n1057), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(G107), .C2(new_n771), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n766), .A2(new_n211), .B1(new_n758), .B2(new_n508), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n245), .B(new_n1073), .C1(G87), .C2(new_n769), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G97), .A2(new_n779), .B1(new_n777), .B2(G116), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n245), .B1(new_n766), .B2(new_n289), .ZN(new_n1077));
  INV_X1    g0877(.A(G128), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n755), .A2(new_n1078), .B1(new_n762), .B2(new_n347), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1077), .B(new_n1079), .C1(G125), .C2(new_n788), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n769), .A2(G150), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1081), .A2(KEYINPUT53), .B1(new_n771), .B2(G137), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1080), .B(new_n1082), .C1(KEYINPUT53), .C2(new_n1081), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(KEYINPUT54), .B(G143), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n823), .A2(new_n778), .B1(new_n780), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1076), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1069), .B1(new_n1086), .B2(new_n748), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n870), .A2(new_n876), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1087), .B1(new_n1089), .B2(new_n746), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n903), .A2(G330), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n442), .A2(new_n889), .B1(new_n886), .B2(new_n672), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n871), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n868), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT112), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n891), .A2(KEYINPUT112), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n706), .A2(new_n696), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n802), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n803), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1095), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n892), .A2(new_n1094), .B1(new_n870), .B2(new_n876), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1093), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1093), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n892), .A2(new_n1094), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1088), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1100), .A2(new_n802), .B1(new_n652), .B2(new_n696), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n1098), .B2(new_n1097), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1106), .B(new_n1108), .C1(new_n1110), .C2(new_n1095), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1105), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1090), .B1(new_n1112), .B2(new_n1065), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n443), .A2(new_n727), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT113), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1115), .A2(new_n901), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1109), .B1(new_n1092), .B2(new_n1091), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n804), .B1(new_n727), .B2(KEYINPUT114), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(KEYINPUT114), .B2(new_n727), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1117), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1106), .A2(new_n1122), .B1(new_n803), .B2(new_n807), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1116), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1124), .A2(new_n1112), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n691), .B1(new_n1124), .B2(new_n1112), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1113), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(G378));
  NOR2_X1   g0928(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1116), .B1(new_n1112), .B2(new_n1129), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n879), .A2(new_n898), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n650), .A2(new_n335), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1132), .A2(new_n299), .A3(new_n845), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n299), .A2(new_n845), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n650), .A2(new_n335), .A3(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT117), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n866), .A2(new_n861), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n859), .A2(new_n852), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n862), .A2(new_n849), .B1(new_n858), .B2(KEYINPUT37), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n872), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n907), .B1(new_n1148), .B2(new_n857), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n708), .B1(new_n1142), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1140), .B1(new_n1150), .B2(new_n908), .ZN(new_n1151));
  AND4_X1   g0951(.A1(new_n1140), .A2(new_n908), .A3(G330), .A4(new_n909), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1139), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n908), .A2(new_n909), .A3(G330), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1139), .B1(new_n1154), .B2(KEYINPUT117), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1131), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1139), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n906), .A2(new_n907), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT38), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n857), .ZN(new_n1161));
  OAI21_X1  g0961(.A(KEYINPUT40), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(G330), .B1(new_n1141), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT117), .B1(new_n1159), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n908), .A2(new_n909), .A3(new_n1140), .A4(G330), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1158), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1166), .A2(new_n899), .A3(new_n1155), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1130), .B1(new_n1157), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT57), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n691), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1153), .A2(new_n1131), .A3(new_n1156), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n899), .B1(new_n1166), .B2(new_n1155), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n1172), .A3(KEYINPUT118), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT118), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1174), .B(new_n899), .C1(new_n1166), .C2(new_n1155), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1173), .A2(new_n1175), .A3(KEYINPUT57), .A4(new_n1130), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1170), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n733), .B1(new_n1157), .B2(new_n1167), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1139), .A2(new_n745), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n754), .A2(G125), .B1(G150), .B2(new_n786), .ZN(new_n1180));
  OR3_X1    g0980(.A1(new_n768), .A2(new_n1084), .A3(KEYINPUT116), .ZN(new_n1181));
  OAI21_X1  g0981(.A(KEYINPUT116), .B1(new_n768), .B2(new_n1084), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n771), .A2(G132), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n778), .A2(new_n1078), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(G137), .C2(new_n779), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n790), .A2(G159), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G33), .B(G41), .C1(new_n788), .C2(G124), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n755), .A2(new_n520), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n933), .B(new_n1193), .C1(G97), .C2(new_n771), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n343), .A2(new_n690), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n768), .A2(new_n247), .B1(new_n766), .B2(new_n210), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(G283), .C2(new_n788), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G107), .A2(new_n777), .B1(new_n779), .B2(new_n308), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1194), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT115), .Z(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT58), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1195), .B(new_n289), .C1(G33), .C2(G41), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(KEYINPUT58), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1192), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n748), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n812), .A2(new_n289), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1179), .A2(new_n735), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1178), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1177), .A2(new_n1209), .ZN(G375));
  OAI21_X1  g1010(.A(new_n733), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT121), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1118), .A2(new_n745), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n735), .B1(G68), .B2(new_n813), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G107), .A2(new_n779), .B1(new_n777), .B2(G283), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n343), .B1(new_n766), .B2(new_n247), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n768), .A2(new_n492), .B1(new_n758), .B2(new_n815), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1032), .B1(new_n755), .B2(new_n508), .C1(new_n520), .C2(new_n1033), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1220), .A2(KEYINPUT119), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(KEYINPUT119), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n245), .B1(new_n766), .B2(new_n210), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n1033), .A2(new_n1084), .B1(new_n289), .B2(new_n762), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(G132), .C2(new_n754), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n779), .A2(G150), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n768), .A2(new_n347), .B1(new_n758), .B2(new_n1078), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT120), .Z(new_n1228));
  NAND2_X1  g1028(.A1(new_n777), .A2(G137), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1225), .A2(new_n1226), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1221), .A2(new_n1222), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1214), .B1(new_n1231), .B2(new_n748), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1213), .A2(new_n1232), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1211), .A2(new_n1212), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1212), .B1(new_n1211), .B2(new_n1233), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1123), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(new_n901), .C2(new_n1115), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n1001), .A3(new_n1124), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1237), .A2(new_n1242), .ZN(G381));
  NAND3_X1  g1043(.A1(new_n1007), .A2(new_n798), .A3(new_n1041), .ZN(new_n1244));
  OR3_X1    g1044(.A1(G390), .A2(G384), .A3(new_n1244), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(G387), .A2(G381), .A3(new_n1245), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1246), .A2(new_n1127), .A3(new_n1177), .A4(new_n1209), .ZN(G407));
  INV_X1    g1047(.A(G213), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(G343), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1127), .A2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(G375), .C2(new_n1250), .ZN(G409));
  NAND2_X1  g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1244), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G390), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT108), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1252), .B2(new_n1244), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1256), .B2(G390), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1003), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1254), .B(new_n1003), .C1(G390), .C2(new_n1256), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1241), .A2(KEYINPUT123), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1263), .B1(new_n1241), .B2(KEYINPUT123), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1124), .A2(new_n734), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n838), .B1(new_n1267), .B2(new_n1236), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G384), .B(new_n1237), .C1(new_n1269), .C2(new_n1264), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1249), .A2(G2897), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1271), .B(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1173), .A2(new_n733), .A3(new_n1175), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(KEYINPUT122), .A3(new_n1207), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1168), .A2(new_n1000), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT122), .B1(new_n1275), .B2(new_n1207), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1127), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1177), .A2(G378), .A3(new_n1209), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1249), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1262), .B1(new_n1274), .B2(new_n1282), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1249), .B(new_n1271), .C1(new_n1280), .C2(new_n1281), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(KEYINPUT63), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n1127), .B(new_n1208), .C1(new_n1170), .C2(new_n1176), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1275), .A2(new_n1207), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT122), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n1277), .A3(new_n1276), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1287), .B1(new_n1127), .B2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT124), .B1(new_n1292), .B2(new_n1249), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT124), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1249), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1271), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1293), .A2(KEYINPUT63), .A3(new_n1297), .A4(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1286), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1274), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1295), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1302));
  AOI211_X1 g1102(.A(KEYINPUT124), .B(new_n1249), .C1(new_n1280), .C2(new_n1281), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1301), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1260), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1293), .A2(KEYINPUT62), .A3(new_n1297), .A4(new_n1298), .ZN(new_n1306));
  AOI211_X1 g1106(.A(KEYINPUT125), .B(KEYINPUT62), .C1(new_n1282), .C2(new_n1298), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT125), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1294), .A2(new_n1296), .A3(new_n1298), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1308), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1307), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1305), .B1(new_n1306), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1314));
  XOR2_X1   g1114(.A(new_n1314), .B(KEYINPUT126), .Z(new_n1315));
  OAI211_X1 g1115(.A(KEYINPUT127), .B(new_n1300), .C1(new_n1313), .C2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT127), .ZN(new_n1317));
  OAI21_X1  g1117(.A(KEYINPUT125), .B1(new_n1284), .B2(KEYINPUT62), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1309), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1306), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1293), .A2(new_n1297), .ZN(new_n1321));
  AOI21_X1  g1121(.A(KEYINPUT61), .B1(new_n1321), .B2(new_n1301), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1315), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1286), .A2(new_n1299), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1317), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1316), .A2(new_n1325), .ZN(G405));
  NAND2_X1  g1126(.A1(G375), .A2(new_n1127), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1281), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(new_n1271), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1315), .B(new_n1329), .ZN(G402));
endmodule


