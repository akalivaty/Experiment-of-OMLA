//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109;
  INV_X1    g000(.A(G224), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G953), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT67), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n192), .B(KEYINPUT1), .C1(new_n189), .C2(G146), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(G128), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n189), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(new_n196), .A3(new_n197), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(new_n200), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n194), .A2(new_n198), .B1(new_n202), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  OR2_X1    g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n196), .A2(new_n197), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n196), .A2(new_n197), .A3(new_n209), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G125), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n188), .B1(new_n207), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n202), .A2(new_n205), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n193), .A2(G128), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n192), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n198), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n213), .ZN(new_n221));
  INV_X1    g035(.A(new_n188), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n221), .B(new_n222), .C1(new_n213), .C2(new_n212), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G110), .B(G122), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G107), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G107), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(G104), .B2(new_n228), .ZN(new_n229));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G107), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT84), .ZN(new_n231));
  INV_X1    g045(.A(G104), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT84), .A2(G104), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT85), .B(G101), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n229), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G101), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(G104), .B2(G107), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n234), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(G107), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  XOR2_X1   g056(.A(KEYINPUT2), .B(G113), .Z(new_n243));
  XNOR2_X1  g057(.A(G116), .B(G119), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT5), .ZN(new_n246));
  INV_X1    g060(.A(G119), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(G116), .ZN(new_n248));
  XOR2_X1   g062(.A(G116), .B(G119), .Z(new_n249));
  OAI211_X1 g063(.A(G113), .B(new_n248), .C1(new_n249), .C2(new_n246), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n242), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n230), .A2(new_n233), .A3(new_n234), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT3), .A2(G107), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n230), .B2(new_n232), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n252), .B(G101), .C1(new_n253), .C2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(KEYINPUT86), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n238), .B1(new_n229), .B2(new_n235), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n252), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT2), .B(G113), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n249), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n245), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n237), .A2(KEYINPUT4), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(new_n259), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n251), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT89), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n226), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n250), .A2(new_n245), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n237), .A2(new_n241), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n263), .A2(new_n245), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n237), .A2(KEYINPUT4), .ZN(new_n274));
  INV_X1    g088(.A(new_n259), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n256), .A2(KEYINPUT86), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n259), .A2(new_n258), .A3(new_n252), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n272), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT89), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n251), .B(new_n226), .C1(new_n261), .C2(new_n266), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n269), .A2(new_n281), .B1(KEYINPUT6), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n226), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n280), .B2(KEYINPUT89), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n268), .B(new_n272), .C1(new_n276), .C2(new_n279), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n225), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G210), .B1(G237), .B2(G902), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n215), .B(new_n223), .C1(KEYINPUT7), .C2(new_n188), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n207), .A2(new_n214), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT7), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n222), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n270), .A2(new_n271), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT90), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n226), .B(KEYINPUT8), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n251), .A2(KEYINPUT90), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n297), .B(new_n298), .C1(new_n299), .C2(new_n295), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n291), .A2(new_n294), .A3(new_n300), .A4(new_n282), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n289), .A2(new_n290), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n290), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n282), .A2(KEYINPUT6), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n307), .B1(new_n285), .B2(new_n287), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n267), .A2(new_n268), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n309), .A2(new_n281), .A3(KEYINPUT6), .A4(new_n284), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n224), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n306), .B1(new_n311), .B2(new_n303), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n305), .A2(new_n312), .A3(KEYINPUT91), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT80), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n213), .A2(G140), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT16), .ZN(new_n318));
  OR3_X1    g132(.A1(new_n213), .A2(KEYINPUT16), .A3(G140), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n314), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n213), .A2(KEYINPUT16), .A3(G140), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(KEYINPUT80), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n195), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n322), .ZN(new_n324));
  XNOR2_X1  g138(.A(G125), .B(G140), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n321), .B1(new_n325), .B2(KEYINPUT16), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n324), .B(G146), .C1(new_n326), .C2(new_n314), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G953), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT72), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G953), .ZN(new_n332));
  INV_X1    g146(.A(G237), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n330), .A2(new_n332), .A3(G214), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n189), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT72), .B(G953), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n336), .A2(G143), .A3(G214), .A4(new_n333), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G131), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT17), .ZN(new_n340));
  INV_X1    g154(.A(G131), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n335), .A2(new_n337), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n341), .B1(new_n335), .B2(new_n337), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT17), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n328), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  XOR2_X1   g160(.A(G113), .B(G122), .Z(new_n347));
  XOR2_X1   g161(.A(KEYINPUT94), .B(G104), .Z(new_n348));
  XOR2_X1   g162(.A(new_n347), .B(new_n348), .Z(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT18), .A2(G131), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n335), .A2(new_n337), .A3(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n325), .B(new_n195), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT92), .ZN(new_n353));
  INV_X1    g167(.A(new_n350), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(new_n338), .B2(new_n354), .ZN(new_n355));
  AOI211_X1 g169(.A(KEYINPUT92), .B(new_n350), .C1(new_n335), .C2(new_n337), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n351), .B(new_n352), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n346), .A2(new_n349), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n349), .B1(new_n346), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n302), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G475), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n362));
  INV_X1    g176(.A(new_n349), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n351), .A2(new_n352), .ZN(new_n364));
  INV_X1    g178(.A(new_n355), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n338), .A2(new_n353), .A3(new_n354), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT19), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT93), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n370));
  MUX2_X1   g184(.A(new_n369), .B(new_n370), .S(new_n325), .Z(new_n371));
  OAI21_X1  g185(.A(new_n327), .B1(new_n371), .B2(G146), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n335), .A2(new_n337), .A3(new_n341), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(new_n344), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n363), .B1(new_n367), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n346), .A2(new_n349), .A3(new_n357), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(G475), .A2(G902), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n362), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n379), .ZN(new_n381));
  AOI211_X1 g195(.A(KEYINPUT20), .B(new_n381), .C1(new_n376), .C2(new_n377), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n361), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G952), .ZN(new_n384));
  AOI211_X1 g198(.A(G953), .B(new_n384), .C1(G234), .C2(G237), .ZN(new_n385));
  AOI211_X1 g199(.A(new_n302), .B(new_n336), .C1(G234), .C2(G237), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT21), .B(G898), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G134), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n189), .A2(G128), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n199), .A2(G143), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT96), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(new_n390), .B2(new_n391), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n391), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT96), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(G134), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G116), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(G122), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n403));
  INV_X1    g217(.A(G122), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(G116), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n402), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n401), .A2(G122), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT97), .B1(new_n407), .B2(KEYINPUT14), .ZN(new_n408));
  OAI211_X1 g222(.A(KEYINPUT97), .B(KEYINPUT14), .C1(new_n404), .C2(G116), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n406), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G107), .ZN(new_n412));
  OR3_X1    g226(.A1(new_n402), .A2(new_n405), .A3(G107), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n400), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G107), .B1(new_n402), .B2(new_n405), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT13), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n391), .B1(new_n390), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n390), .A2(new_n417), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT95), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT95), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n390), .A2(new_n421), .A3(new_n417), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n418), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n416), .B(new_n395), .C1(new_n423), .C2(new_n389), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n414), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT9), .B(G234), .ZN(new_n426));
  INV_X1    g240(.A(G217), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n426), .A2(new_n427), .A3(G953), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT98), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n414), .A2(new_n429), .A3(new_n424), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n302), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G478), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT15), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n433), .B(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n383), .A2(new_n388), .A3(new_n436), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n311), .A2(new_n306), .A3(new_n303), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT91), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(G214), .B1(G237), .B2(G902), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n313), .A2(new_n437), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(new_n302), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n190), .A2(G128), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n198), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n204), .B1(new_n203), .B2(new_n200), .ZN(new_n447));
  AND4_X1   g261(.A1(new_n204), .A2(new_n200), .A3(new_n196), .A4(new_n197), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT87), .B1(new_n242), .B2(new_n449), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n202), .A2(new_n205), .B1(new_n198), .B2(new_n445), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n451), .A2(new_n271), .A3(new_n452), .ZN(new_n453));
  OAI22_X1  g267(.A1(new_n450), .A2(new_n453), .B1(new_n220), .B2(new_n242), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT11), .B1(new_n389), .B2(G137), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT11), .ZN(new_n456));
  INV_X1    g270(.A(G137), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(G134), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT64), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n457), .B2(G134), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n389), .A2(KEYINPUT64), .A3(G137), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(KEYINPUT65), .A2(G131), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n461), .A2(new_n462), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n464), .A3(new_n459), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n454), .A2(KEYINPUT12), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT12), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n242), .A2(KEYINPUT87), .A3(new_n449), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n452), .B1(new_n451), .B2(new_n271), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n472), .A2(new_n473), .B1(new_n206), .B2(new_n271), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n455), .A2(new_n458), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n461), .A2(new_n462), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n475), .A2(new_n465), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n464), .B1(new_n467), .B2(new_n459), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n471), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT10), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n450), .B2(new_n453), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT69), .B1(new_n210), .B2(new_n211), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n196), .A2(new_n197), .A3(new_n209), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT69), .ZN(new_n486));
  INV_X1    g300(.A(new_n209), .ZN(new_n487));
  NOR2_X1   g301(.A1(KEYINPUT0), .A2(G128), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n485), .B(new_n486), .C1(new_n489), .C2(new_n203), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n484), .B(new_n490), .C1(new_n265), .C2(new_n259), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n279), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n469), .B(KEYINPUT88), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n242), .A2(new_n220), .A3(KEYINPUT10), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n483), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n481), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n336), .A2(G227), .ZN(new_n498));
  XOR2_X1   g312(.A(G110), .B(G140), .Z(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n495), .B1(new_n261), .B2(new_n491), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT10), .B1(new_n472), .B2(new_n473), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n469), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n501), .A2(new_n502), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n500), .B1(new_n504), .B2(new_n494), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n497), .A2(new_n500), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n444), .B1(new_n506), .B2(G469), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n481), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n503), .A2(new_n496), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n500), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n443), .A3(new_n302), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G221), .B1(new_n426), .B2(G902), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n442), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(G221), .A2(G234), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n336), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT81), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT81), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n336), .A2(new_n520), .A3(new_n517), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT22), .B(G137), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n519), .A2(new_n521), .A3(new_n523), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT79), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT23), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT23), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT79), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n199), .A2(G119), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G110), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n247), .A2(G128), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n533), .A2(new_n529), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n535), .A2(new_n536), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT78), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n533), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n540), .B1(new_n533), .B2(new_n537), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT24), .B(G110), .Z(new_n545));
  OAI21_X1  g359(.A(new_n539), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n325), .A2(new_n195), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n327), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n543), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n541), .A3(new_n545), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n538), .A2(new_n537), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n533), .B1(new_n529), .B2(new_n531), .ZN(new_n553));
  OAI21_X1  g367(.A(G110), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n323), .B2(new_n327), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n527), .B1(new_n549), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n323), .A2(new_n327), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(new_n551), .A3(new_n554), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n559), .A2(new_n548), .A3(new_n526), .A4(new_n525), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n427), .B1(G234), .B2(new_n302), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(G902), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT25), .ZN(new_n567));
  AOI21_X1  g381(.A(G902), .B1(new_n567), .B2(KEYINPUT82), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n557), .A2(new_n560), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n567), .A2(KEYINPUT82), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n570), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n557), .A2(new_n560), .A3(new_n572), .A4(new_n568), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(new_n573), .A3(new_n562), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n561), .A2(KEYINPUT83), .A3(new_n563), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n566), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n336), .A2(G210), .A3(new_n333), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT26), .B(G101), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT28), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT68), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n389), .A2(G137), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n457), .A2(G134), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n585), .A2(new_n586), .A3(new_n341), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n463), .B2(new_n341), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n584), .B1(new_n206), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n341), .B1(new_n475), .B2(new_n476), .ZN(new_n590));
  INV_X1    g404(.A(new_n587), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(new_n220), .A3(KEYINPUT68), .ZN(new_n593));
  OAI22_X1  g407(.A1(new_n477), .A2(new_n478), .B1(new_n210), .B2(new_n211), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n589), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n264), .ZN(new_n596));
  INV_X1    g410(.A(new_n490), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT0), .B(G128), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n198), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n486), .B1(new_n599), .B2(new_n485), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n601), .A2(new_n469), .B1(new_n592), .B2(new_n220), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n264), .B(KEYINPUT71), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n583), .B1(new_n596), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT71), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n264), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n484), .A2(new_n490), .ZN(new_n608));
  OAI22_X1  g422(.A1(new_n479), .A2(new_n608), .B1(new_n206), .B2(new_n588), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT75), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n602), .A2(KEYINPUT75), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT28), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n582), .B1(new_n605), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n604), .A2(KEYINPUT74), .A3(new_n581), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(KEYINPUT31), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT30), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n595), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT70), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n602), .B2(KEYINPUT30), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n592), .A2(new_n220), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n484), .B(new_n490), .C1(new_n477), .C2(new_n478), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n619), .A4(KEYINPUT30), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n618), .B(new_n264), .C1(new_n620), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n616), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT70), .B1(new_n609), .B2(new_n617), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n627), .A2(new_n623), .B1(new_n617), .B2(new_n595), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n615), .B1(new_n628), .B2(new_n264), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT31), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n614), .B(new_n626), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(G472), .A2(G902), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT76), .Z(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT32), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT32), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n631), .A2(new_n637), .A3(new_n634), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n603), .B1(new_n602), .B2(KEYINPUT75), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n609), .A2(new_n610), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n583), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n602), .A2(new_n603), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n609), .A2(new_n607), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT28), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n581), .A2(KEYINPUT29), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n642), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT77), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT77), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n642), .A2(new_n645), .A3(new_n649), .A4(new_n646), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n302), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n581), .B1(new_n605), .B2(new_n613), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n625), .A2(new_n604), .A3(new_n582), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT29), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(G472), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n576), .B1(new_n639), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n516), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(new_n236), .Z(G3));
  INV_X1    g472(.A(new_n514), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n507), .B2(new_n512), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n631), .A2(new_n302), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n661), .B2(KEYINPUT99), .ZN(new_n662));
  INV_X1    g476(.A(new_n615), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n625), .A2(new_n663), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n664), .A2(KEYINPUT31), .B1(new_n625), .B2(new_n616), .ZN(new_n665));
  AOI21_X1  g479(.A(G902), .B1(new_n665), .B2(new_n614), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n660), .B(new_n635), .C1(new_n662), .C2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n576), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n290), .B1(new_n289), .B2(new_n304), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n441), .B1(new_n672), .B2(new_n438), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n434), .A2(G902), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT33), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n414), .A2(new_n429), .A3(new_n424), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n429), .B1(new_n414), .B2(new_n424), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n431), .A2(KEYINPUT33), .A3(new_n432), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT100), .B1(new_n433), .B2(new_n434), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI211_X1 g497(.A(KEYINPUT100), .B(new_n675), .C1(new_n679), .C2(new_n680), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT101), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n679), .A2(new_n680), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n687), .A3(new_n674), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n688), .B(new_n689), .C1(new_n681), .C2(new_n682), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n685), .A2(new_n383), .A3(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n673), .A2(new_n388), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n670), .A2(new_n671), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT34), .B(G104), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G6));
  INV_X1    g509(.A(new_n441), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n305), .B2(new_n312), .ZN(new_n697));
  INV_X1    g511(.A(new_n388), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n361), .B(new_n436), .C1(new_n380), .C2(new_n382), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n670), .A2(new_n671), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT35), .B(G107), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G9));
  INV_X1    g518(.A(new_n442), .ZN(new_n705));
  INV_X1    g519(.A(new_n635), .ZN(new_n706));
  INV_X1    g520(.A(G472), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n666), .B2(new_n667), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n661), .A2(KEYINPUT99), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI22_X1  g524(.A1(new_n549), .A2(new_n556), .B1(KEYINPUT36), .B2(new_n527), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n527), .A2(KEYINPUT36), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n559), .A3(new_n548), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n711), .A2(new_n713), .A3(new_n563), .ZN(new_n714));
  INV_X1    g528(.A(new_n562), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n569), .B2(new_n570), .ZN(new_n716));
  AOI211_X1 g530(.A(KEYINPUT102), .B(new_n714), .C1(new_n716), .C2(new_n573), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n718));
  INV_X1    g532(.A(new_n714), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n718), .B1(new_n574), .B2(new_n719), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n705), .A2(new_n710), .A3(new_n660), .A4(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT37), .B(G110), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G12));
  AND3_X1   g538(.A1(new_n631), .A2(new_n637), .A3(new_n634), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n637), .B1(new_n631), .B2(new_n634), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n655), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n727), .A2(new_n660), .A3(new_n721), .ZN(new_n728));
  INV_X1    g542(.A(G900), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n386), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n385), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n700), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT103), .B1(new_n673), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT103), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n699), .A2(new_n731), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n697), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n728), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G128), .ZN(G30));
  XOR2_X1   g554(.A(new_n731), .B(KEYINPUT39), .Z(new_n741));
  NAND2_X1  g555(.A1(new_n660), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(KEYINPUT40), .Z(new_n743));
  NAND2_X1  g557(.A1(new_n313), .A2(new_n440), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT38), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT38), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n313), .A2(new_n746), .A3(new_n440), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n625), .A2(new_n604), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n581), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n643), .A2(new_n644), .ZN(new_n752));
  AOI21_X1  g566(.A(G902), .B1(new_n752), .B2(new_n582), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n707), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n754), .B1(new_n636), .B2(new_n638), .ZN(new_n755));
  OAI221_X1 g569(.A(new_n327), .B1(new_n371), .B2(G146), .C1(new_n344), .C2(new_n373), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n349), .B1(new_n756), .B2(new_n357), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n379), .B1(new_n358), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT20), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n378), .A2(new_n362), .A3(new_n379), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n759), .A2(new_n760), .B1(G475), .B2(new_n360), .ZN(new_n761));
  INV_X1    g575(.A(new_n436), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n755), .A2(new_n696), .A3(new_n721), .A4(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n743), .A2(new_n749), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G143), .ZN(G45));
  NAND4_X1  g581(.A1(new_n685), .A2(new_n383), .A3(new_n690), .A4(new_n732), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n673), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n727), .A3(new_n660), .A4(new_n721), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G146), .ZN(G48));
  AOI22_X1  g585(.A1(new_n481), .A2(new_n505), .B1(new_n509), .B2(new_n500), .ZN(new_n772));
  OAI21_X1  g586(.A(G469), .B1(new_n772), .B2(G902), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n512), .A3(new_n514), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n692), .A2(new_n727), .A3(new_n671), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(KEYINPUT41), .B(G113), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT104), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n776), .B(new_n778), .ZN(G15));
  NAND4_X1  g593(.A1(new_n701), .A2(new_n727), .A3(new_n671), .A4(new_n775), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G116), .ZN(G18));
  NOR2_X1   g595(.A1(new_n717), .A2(new_n720), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n639), .B2(new_n655), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT105), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n673), .A2(new_n774), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n437), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n727), .A2(new_n721), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n775), .A2(new_n437), .A3(new_n697), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT105), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G119), .ZN(G21));
  NAND2_X1  g605(.A1(new_n642), .A2(new_n645), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n582), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n665), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n634), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n795), .B(new_n671), .C1(new_n666), .C2(new_n707), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n305), .A2(new_n312), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n763), .A3(new_n441), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n773), .A2(new_n512), .A3(new_n514), .A4(new_n698), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n404), .ZN(G24));
  AOI21_X1  g615(.A(new_n707), .B1(new_n631), .B2(new_n302), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n633), .B1(new_n665), .B2(new_n793), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n782), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n768), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n785), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G125), .ZN(G27));
  INV_X1    g621(.A(KEYINPUT42), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n768), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n727), .A2(new_n809), .A3(new_n671), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n744), .A2(new_n660), .A3(new_n441), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT106), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n744), .A2(new_n660), .A3(new_n441), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT106), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n656), .A3(new_n814), .A4(new_n809), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n656), .A3(new_n805), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n812), .A2(new_n815), .B1(new_n816), .B2(new_n808), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(new_n341), .ZN(G33));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n656), .A3(new_n736), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G134), .ZN(G36));
  INV_X1    g634(.A(new_n512), .ZN(new_n821));
  INV_X1    g635(.A(new_n444), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n506), .A2(KEYINPUT45), .ZN(new_n823));
  INV_X1    g637(.A(new_n500), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n503), .A2(new_n496), .A3(new_n824), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n470), .A2(new_n480), .B1(new_n504), .B2(new_n494), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n825), .B1(new_n826), .B2(new_n824), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT45), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n443), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT107), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n823), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI211_X1 g645(.A(KEYINPUT107), .B(new_n443), .C1(new_n827), .C2(new_n828), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n822), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT46), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n821), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(KEYINPUT46), .B(new_n822), .C1(new_n831), .C2(new_n832), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n659), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n685), .A2(new_n761), .A3(new_n690), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT43), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT43), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n685), .A2(new_n761), .A3(new_n840), .A4(new_n690), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n839), .A2(new_n721), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT44), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n635), .B1(new_n662), .B2(new_n668), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n839), .A2(new_n721), .A3(new_n841), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT44), .B1(new_n710), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n696), .B1(new_n313), .B2(new_n440), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT108), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n837), .A2(new_n848), .A3(new_n741), .A4(new_n850), .ZN(new_n851));
  XOR2_X1   g665(.A(KEYINPUT109), .B(G137), .Z(new_n852));
  XNOR2_X1  g666(.A(new_n851), .B(new_n852), .ZN(G39));
  INV_X1    g667(.A(new_n849), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n854), .A2(new_n727), .A3(new_n671), .A4(new_n768), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT47), .ZN(new_n856));
  AOI211_X1 g670(.A(new_n856), .B(new_n659), .C1(new_n835), .C2(new_n836), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n833), .A2(new_n834), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n512), .A3(new_n836), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT47), .B1(new_n859), .B2(new_n514), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n855), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(G140), .ZN(G42));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n802), .A2(new_n803), .A3(new_n576), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n385), .A3(new_n839), .A4(new_n841), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n850), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n857), .A2(new_n860), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n773), .A2(new_n512), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n659), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT114), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n867), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n755), .A2(new_n671), .A3(new_n385), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n849), .A2(new_n775), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n685), .A2(new_n690), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n873), .A2(new_n874), .A3(new_n383), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n839), .A2(new_n385), .A3(new_n841), .ZN(new_n877));
  OR3_X1    g691(.A1(new_n874), .A2(new_n877), .A3(KEYINPUT116), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT116), .B1(new_n874), .B2(new_n877), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n876), .B1(new_n880), .B2(new_n804), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n775), .A2(new_n696), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT115), .B1(new_n749), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n882), .B1(new_n745), .B2(new_n747), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n865), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n883), .A2(new_n886), .A3(KEYINPUT50), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT50), .B1(new_n883), .B2(new_n886), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n881), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n863), .B1(new_n872), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n859), .A2(new_n514), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n856), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n837), .A2(KEYINPUT47), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n893), .A3(new_n870), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(new_n850), .A3(new_n866), .ZN(new_n895));
  INV_X1    g709(.A(new_n888), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n883), .A2(new_n886), .A3(KEYINPUT50), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n895), .A2(new_n898), .A3(KEYINPUT51), .A4(new_n881), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n384), .B(G953), .C1(new_n866), .C2(new_n785), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n873), .A2(new_n874), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n900), .B1(new_n691), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n880), .A2(new_n656), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n903), .A2(KEYINPUT48), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(KEYINPUT48), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n890), .A2(new_n899), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n908));
  INV_X1    g722(.A(new_n798), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n698), .A3(new_n775), .A4(new_n864), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n776), .A2(new_n780), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n786), .B2(new_n789), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n722), .A2(new_n657), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n804), .A2(new_n849), .A3(new_n660), .A4(new_n805), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n849), .A2(new_n727), .A3(new_n671), .A4(new_n660), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n733), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n708), .A2(new_n709), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n917), .A2(new_n635), .A3(new_n671), .A4(new_n660), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n388), .B1(new_n691), .B2(new_n699), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n919), .A2(new_n441), .A3(new_n440), .A4(new_n313), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n913), .A2(new_n916), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n815), .A2(new_n812), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n816), .A2(new_n808), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n727), .A2(new_n660), .A3(new_n721), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n761), .A2(new_n762), .A3(new_n732), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n849), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT111), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n696), .B(new_n927), .C1(new_n313), .C2(new_n440), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT111), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n931), .A2(new_n783), .A3(new_n932), .A4(new_n660), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n912), .A2(new_n922), .A3(new_n925), .A4(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT52), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n735), .A2(new_n797), .A3(new_n736), .A4(new_n441), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n735), .B1(new_n697), .B2(new_n736), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n770), .B(new_n806), .C1(new_n939), .C2(new_n926), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n574), .A2(new_n719), .A3(new_n732), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n515), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n755), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n943), .A3(new_n909), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n936), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  NOR4_X1   g760(.A1(new_n768), .A2(new_n782), .A3(new_n802), .A4(new_n803), .ZN(new_n947));
  AOI22_X1  g761(.A1(new_n728), .A2(new_n738), .B1(new_n947), .B2(new_n785), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n948), .A2(KEYINPUT52), .A3(new_n770), .A4(new_n944), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n908), .B1(new_n935), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n442), .A2(new_n782), .ZN(new_n952));
  AOI22_X1  g766(.A1(new_n670), .A2(new_n952), .B1(new_n516), .B2(new_n656), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n691), .A2(new_n699), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n698), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n313), .A2(new_n441), .A3(new_n440), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n670), .A2(new_n957), .A3(new_n671), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n953), .A2(new_n819), .A3(new_n958), .A4(new_n914), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n930), .A2(new_n933), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(new_n908), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n727), .A2(new_n775), .A3(new_n671), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n800), .B1(new_n962), .B2(new_n692), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n790), .A2(new_n963), .A3(new_n780), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT112), .B1(new_n964), .B2(new_n817), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT112), .ZN(new_n966));
  INV_X1    g780(.A(new_n911), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n925), .A2(new_n966), .A3(new_n790), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n946), .A2(new_n949), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n961), .A2(new_n965), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT54), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n951), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT113), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n964), .A2(new_n817), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n959), .A2(new_n960), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n974), .A2(new_n975), .A3(new_n969), .A4(KEYINPUT53), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n971), .B1(new_n951), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT113), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n951), .A2(new_n970), .A3(new_n979), .A4(new_n971), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n907), .A2(new_n973), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT117), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n951), .A2(new_n971), .A3(new_n970), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n977), .B1(new_n983), .B2(new_n979), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT117), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n984), .A2(new_n985), .A3(new_n973), .A4(new_n907), .ZN(new_n986));
  NOR2_X1   g800(.A1(G952), .A2(G953), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT118), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n982), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n869), .A2(KEYINPUT49), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n869), .A2(KEYINPUT49), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n838), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n576), .A2(new_n659), .A3(new_n696), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT110), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n992), .A2(new_n748), .A3(new_n755), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n989), .A2(new_n995), .ZN(G75));
  NOR2_X1   g810(.A1(new_n336), .A2(G952), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n302), .B1(new_n951), .B2(new_n970), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(G210), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n308), .A2(new_n310), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT119), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT55), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(new_n224), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n1005), .A2(KEYINPUT56), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n998), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(KEYINPUT56), .B1(new_n1000), .B2(KEYINPUT120), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(KEYINPUT120), .B2(new_n1000), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1007), .B1(new_n1009), .B2(new_n1005), .ZN(G51));
  NAND2_X1  g824(.A1(new_n951), .A2(new_n970), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(KEYINPUT54), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n972), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n444), .B(KEYINPUT57), .Z(new_n1015));
  OAI21_X1  g829(.A(new_n511), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n829), .A2(new_n830), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n827), .A2(new_n828), .ZN(new_n1018));
  OAI21_X1  g832(.A(G469), .B1(new_n506), .B2(KEYINPUT45), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(KEYINPUT107), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n999), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n997), .B1(new_n1016), .B2(new_n1021), .ZN(G54));
  AND2_X1   g836(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n999), .A2(new_n378), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT121), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n378), .B1(new_n999), .B2(new_n1023), .ZN(new_n1028));
  NOR4_X1   g842(.A1(new_n1026), .A2(new_n1027), .A3(new_n997), .A4(new_n1028), .ZN(G60));
  INV_X1    g843(.A(KEYINPUT122), .ZN(new_n1030));
  NAND2_X1  g844(.A1(G478), .A2(G902), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1031), .B(KEYINPUT59), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n686), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1030), .B1(new_n1013), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n971), .B1(new_n951), .B2(new_n970), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n1030), .B(new_n1033), .C1(new_n983), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n998), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n984), .A2(new_n973), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n686), .B1(new_n1039), .B2(new_n1032), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1038), .A2(new_n1040), .ZN(G63));
  NAND2_X1  g855(.A1(G217), .A2(G902), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(KEYINPUT123), .Z(new_n1043));
  XNOR2_X1  g857(.A(new_n1043), .B(KEYINPUT60), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1044), .B1(new_n951), .B2(new_n970), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1045), .A2(new_n713), .A3(new_n711), .ZN(new_n1046));
  OAI211_X1 g860(.A(new_n1046), .B(new_n998), .C1(new_n561), .C2(new_n1045), .ZN(new_n1047));
  INV_X1    g861(.A(KEYINPUT61), .ZN(new_n1048));
  XNOR2_X1  g862(.A(new_n1047), .B(new_n1048), .ZN(G66));
  OAI21_X1  g863(.A(G953), .B1(new_n387), .B2(new_n187), .ZN(new_n1050));
  NOR3_X1   g864(.A1(new_n964), .A2(new_n921), .A3(new_n913), .ZN(new_n1051));
  INV_X1    g865(.A(new_n336), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1003), .B1(G898), .B2(new_n336), .ZN(new_n1054));
  XNOR2_X1  g868(.A(new_n1053), .B(new_n1054), .ZN(G69));
  XOR2_X1   g869(.A(new_n628), .B(new_n371), .Z(new_n1056));
  INV_X1    g870(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g871(.A(G227), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1052), .A2(G900), .ZN(new_n1059));
  INV_X1    g873(.A(new_n940), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n766), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g875(.A(new_n1061), .B(KEYINPUT62), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n727), .A2(new_n671), .ZN(new_n1063));
  NAND4_X1  g877(.A1(new_n849), .A2(new_n660), .A3(new_n741), .A4(new_n954), .ZN(new_n1064));
  OAI211_X1 g878(.A(new_n861), .B(new_n851), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  OR2_X1    g879(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  OAI221_X1 g880(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .C1(new_n1066), .C2(new_n1052), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n843), .B1(new_n842), .B2(new_n844), .ZN(new_n1068));
  NOR3_X1   g882(.A1(new_n710), .A2(new_n846), .A3(KEYINPUT44), .ZN(new_n1069));
  OAI21_X1  g883(.A(new_n850), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n444), .B1(new_n1020), .B2(new_n1017), .ZN(new_n1071));
  OAI21_X1  g885(.A(new_n512), .B1(new_n1071), .B2(KEYINPUT46), .ZN(new_n1072));
  INV_X1    g886(.A(new_n836), .ZN(new_n1073));
  OAI211_X1 g887(.A(new_n514), .B(new_n741), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g888(.A(KEYINPUT124), .B(new_n1060), .C1(new_n1070), .C2(new_n1074), .ZN(new_n1075));
  INV_X1    g889(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g890(.A(KEYINPUT124), .B1(new_n851), .B2(new_n1060), .ZN(new_n1077));
  NOR2_X1   g891(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g892(.A1(new_n1063), .A2(new_n798), .ZN(new_n1079));
  NAND4_X1  g893(.A1(new_n859), .A2(new_n514), .A3(new_n741), .A4(new_n1079), .ZN(new_n1080));
  NAND4_X1  g894(.A1(new_n861), .A2(new_n925), .A3(new_n819), .A4(new_n1080), .ZN(new_n1081));
  OAI21_X1  g895(.A(KEYINPUT125), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g896(.A(new_n855), .ZN(new_n1083));
  AOI21_X1  g897(.A(new_n1083), .B1(new_n892), .B2(new_n893), .ZN(new_n1084));
  NAND3_X1  g898(.A1(new_n925), .A2(new_n819), .A3(new_n1080), .ZN(new_n1085));
  NOR2_X1   g899(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g900(.A(KEYINPUT125), .ZN(new_n1087));
  OAI211_X1 g901(.A(new_n1086), .B(new_n1087), .C1(new_n1077), .C2(new_n1076), .ZN(new_n1088));
  AOI21_X1  g902(.A(new_n1052), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g903(.A(new_n1056), .B1(G227), .B2(new_n1059), .ZN(new_n1090));
  OAI21_X1  g904(.A(new_n1067), .B1(new_n1089), .B2(new_n1090), .ZN(G72));
  NAND2_X1  g905(.A1(G472), .A2(G902), .ZN(new_n1092));
  XOR2_X1   g906(.A(new_n1092), .B(KEYINPUT63), .Z(new_n1093));
  INV_X1    g907(.A(new_n1051), .ZN(new_n1094));
  OAI21_X1  g908(.A(new_n1093), .B1(new_n1066), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g909(.A(new_n751), .ZN(new_n1096));
  NAND2_X1  g910(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g911(.A1(new_n951), .A2(new_n976), .ZN(new_n1098));
  NAND4_X1  g912(.A1(new_n1098), .A2(new_n653), .A3(new_n751), .A4(new_n1093), .ZN(new_n1099));
  NAND2_X1  g913(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g914(.A1(new_n1082), .A2(new_n1051), .A3(new_n1088), .ZN(new_n1101));
  NAND2_X1  g915(.A1(new_n1101), .A2(new_n1093), .ZN(new_n1102));
  XNOR2_X1  g916(.A(new_n653), .B(KEYINPUT126), .ZN(new_n1103));
  NAND2_X1  g917(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g918(.A(KEYINPUT127), .ZN(new_n1105));
  NAND3_X1  g919(.A1(new_n1104), .A2(new_n1105), .A3(new_n998), .ZN(new_n1106));
  INV_X1    g920(.A(new_n1103), .ZN(new_n1107));
  AOI21_X1  g921(.A(new_n1107), .B1(new_n1101), .B2(new_n1093), .ZN(new_n1108));
  OAI21_X1  g922(.A(KEYINPUT127), .B1(new_n1108), .B2(new_n997), .ZN(new_n1109));
  AOI21_X1  g923(.A(new_n1100), .B1(new_n1106), .B2(new_n1109), .ZN(G57));
endmodule


