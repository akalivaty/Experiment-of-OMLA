//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  OR2_X1    g000(.A1(KEYINPUT72), .A2(G953), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT72), .A2(G953), .ZN(new_n189));
  NAND4_X1  g003(.A1(new_n187), .A2(G214), .A3(new_n188), .A4(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT72), .A2(G953), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT72), .A2(G953), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n195), .A2(G143), .A3(G214), .A4(new_n188), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT18), .A2(G131), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n197), .B(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n204), .A2(KEYINPUT90), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(KEYINPUT90), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(G146), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n204), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n199), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT91), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n197), .A2(new_n198), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n197), .A2(new_n198), .ZN(new_n216));
  OAI211_X1 g030(.A(KEYINPUT91), .B(new_n211), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G113), .B(G122), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n219), .B(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT92), .B1(new_n197), .B2(G131), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT92), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  AOI211_X1 g038(.A(new_n223), .B(new_n224), .C1(new_n192), .C2(new_n196), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT17), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT16), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n200), .A3(G125), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n228), .B1(new_n204), .B2(new_n227), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n209), .ZN(new_n230));
  OAI211_X1 g044(.A(G146), .B(new_n228), .C1(new_n204), .C2(new_n227), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n226), .A2(KEYINPUT93), .A3(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n222), .A2(new_n225), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT17), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n192), .A2(new_n196), .A3(new_n224), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT93), .B1(new_n226), .B2(new_n233), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n218), .B(new_n221), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n221), .ZN(new_n242));
  INV_X1    g056(.A(new_n217), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT91), .B1(new_n199), .B2(new_n211), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n205), .A2(KEYINPUT19), .A3(new_n206), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(KEYINPUT19), .B2(new_n204), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n231), .B1(new_n247), .B2(G146), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n235), .B2(new_n237), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n242), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n241), .A2(KEYINPUT94), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT94), .B1(new_n241), .B2(new_n250), .ZN(new_n252));
  NOR2_X1   g066(.A1(G475), .A2(G902), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT20), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT95), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n252), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n241), .A2(KEYINPUT94), .A3(new_n250), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n253), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT95), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT20), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n241), .A2(new_n250), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n254), .A2(KEYINPUT20), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n257), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G902), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n218), .B1(new_n239), .B2(new_n240), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n242), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT96), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n241), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n267), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G475), .ZN(new_n274));
  XNOR2_X1  g088(.A(G128), .B(G143), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT98), .ZN(new_n276));
  INV_X1    g090(.A(G134), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT97), .B(KEYINPUT13), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(G128), .A3(new_n191), .ZN(new_n280));
  INV_X1    g094(.A(new_n275), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n280), .B(G134), .C1(new_n281), .C2(new_n279), .ZN(new_n282));
  XOR2_X1   g096(.A(G116), .B(G122), .Z(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(G107), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n278), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G107), .ZN(new_n287));
  INV_X1    g101(.A(G116), .ZN(new_n288));
  OR2_X1    g102(.A1(new_n288), .A2(G122), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n287), .B1(new_n289), .B2(KEYINPUT14), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n290), .B(new_n283), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT98), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n275), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G134), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n291), .B1(new_n278), .B2(new_n294), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n286), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  INV_X1    g111(.A(G217), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n297), .A2(new_n298), .A3(G953), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(KEYINPUT100), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n300), .B1(new_n286), .B2(new_n295), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT100), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n286), .A2(new_n295), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n305), .A2(KEYINPUT99), .A3(new_n299), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT99), .B1(new_n305), .B2(new_n299), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n301), .B(new_n304), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n267), .ZN(new_n309));
  INV_X1    g123(.A(G478), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT15), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n311), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(new_n308), .B2(new_n267), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G953), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n316), .A2(G952), .ZN(new_n317));
  INV_X1    g131(.A(G234), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(new_n188), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI211_X1 g134(.A(new_n267), .B(new_n195), .C1(G234), .C2(G237), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT21), .B(G898), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AND4_X1   g138(.A1(new_n266), .A2(new_n274), .A3(new_n315), .A4(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G469), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n195), .A2(G227), .ZN(new_n327));
  XOR2_X1   g141(.A(G110), .B(G140), .Z(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT86), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n191), .A2(G146), .ZN(new_n333));
  OAI21_X1  g147(.A(G128), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT64), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n209), .A3(G143), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT64), .B1(new_n191), .B2(G146), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(new_n333), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT1), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT68), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT68), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT1), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n341), .A2(new_n343), .A3(G128), .ZN(new_n344));
  XNOR2_X1  g158(.A(G143), .B(G146), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT71), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n334), .A2(new_n338), .B1(new_n345), .B2(new_n344), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT71), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n352));
  XNOR2_X1  g166(.A(G104), .B(G107), .ZN(new_n353));
  INV_X1    g167(.A(G101), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT3), .B1(new_n220), .B2(G107), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(new_n287), .A3(G104), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n220), .A2(G107), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n356), .A2(new_n358), .A3(new_n354), .A4(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n220), .A2(G107), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n287), .A2(G104), .ZN(new_n362));
  OAI211_X1 g176(.A(KEYINPUT82), .B(G101), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n355), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n349), .A2(new_n351), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G101), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT4), .A3(new_n360), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT65), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n191), .A2(KEYINPUT64), .A3(G146), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n209), .A2(G143), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n335), .B1(new_n209), .B2(G143), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AND2_X1   g191(.A1(KEYINPUT0), .A2(G128), .ZN(new_n378));
  NOR2_X1   g192(.A1(KEYINPUT0), .A2(G128), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n373), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n338), .A2(KEYINPUT65), .A3(new_n380), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n345), .A2(new_n378), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n369), .A2(KEYINPUT4), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n367), .B1(new_n372), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n191), .A2(G146), .ZN(new_n389));
  AOI21_X1  g203(.A(G128), .B1(new_n375), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n191), .A2(KEYINPUT1), .A3(G146), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT83), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n394), .B(new_n391), .C1(new_n345), .C2(G128), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n346), .A3(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n355), .A2(new_n360), .A3(new_n363), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT84), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT84), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT10), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n331), .B1(new_n388), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT11), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n404), .B1(new_n277), .B2(G137), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n277), .A2(G137), .ZN(new_n406));
  INV_X1    g220(.A(G137), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT11), .A3(G134), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G131), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n405), .A2(new_n408), .A3(new_n224), .A4(new_n406), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n396), .A2(new_n397), .A3(new_n400), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n400), .B1(new_n396), .B2(new_n397), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n365), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n382), .A2(new_n383), .B1(new_n345), .B2(new_n378), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n370), .A2(KEYINPUT81), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n370), .A2(KEYINPUT81), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n416), .B(new_n386), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n415), .A2(new_n419), .A3(KEYINPUT86), .A4(new_n367), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n403), .A2(new_n412), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT87), .ZN(new_n422));
  INV_X1    g236(.A(new_n412), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n415), .A2(new_n419), .A3(new_n367), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n424), .B2(new_n331), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT87), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(new_n420), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n412), .B(KEYINPUT85), .Z(new_n429));
  OR2_X1    g243(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n330), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI22_X1  g245(.A1(new_n413), .A2(new_n414), .B1(new_n347), .B2(new_n397), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n412), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT12), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n435), .A2(new_n430), .A3(new_n330), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n326), .B(new_n267), .C1(new_n431), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n430), .A2(new_n330), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n428), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n330), .B1(new_n435), .B2(new_n430), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n442), .A3(G469), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n326), .A2(new_n267), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n437), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G210), .B1(G237), .B2(G902), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT69), .B1(new_n288), .B2(G119), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT69), .ZN(new_n451));
  INV_X1    g265(.A(G119), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(G116), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT70), .B1(new_n452), .B2(G116), .ZN(new_n455));
  OR3_X1    g269(.A1(new_n452), .A2(KEYINPUT70), .A3(G116), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT2), .B(G113), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n458), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n460), .A2(new_n454), .A3(new_n455), .A4(new_n456), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n462), .B(new_n386), .C1(new_n417), .C2(new_n418), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G122), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n288), .A2(KEYINPUT5), .A3(G119), .ZN(new_n465));
  INV_X1    g279(.A(G113), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT5), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n467), .B1(new_n457), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n397), .A2(new_n469), .A3(new_n461), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT88), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n470), .A2(new_n471), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n463), .B(new_n464), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n469), .A2(new_n461), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n364), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n470), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(KEYINPUT89), .A3(new_n364), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n464), .B(KEYINPUT8), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n350), .A2(new_n202), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n416), .B2(new_n202), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n316), .A2(G224), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n474), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n485), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n482), .B(new_n485), .C1(new_n416), .C2(new_n202), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI22_X1  g305(.A1(new_n489), .A2(new_n491), .B1(KEYINPUT7), .B2(new_n488), .ZN(new_n492));
  AOI21_X1  g306(.A(G902), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n463), .B1(new_n472), .B2(new_n473), .ZN(new_n494));
  INV_X1    g308(.A(new_n464), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT6), .A3(new_n474), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n489), .A2(new_n491), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(new_n499), .A3(new_n495), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n449), .B1(new_n493), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n493), .A2(new_n501), .A3(new_n449), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n448), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G221), .B1(new_n297), .B2(G902), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n446), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n298), .B1(G234), .B2(new_n267), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT79), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(KEYINPUT25), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT22), .B(G137), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n452), .A2(G128), .ZN(new_n516));
  INV_X1    g330(.A(G128), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G119), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT24), .B(G110), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(KEYINPUT23), .A3(G119), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n452), .A2(G128), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(new_n516), .C1(new_n523), .C2(KEYINPUT23), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n521), .B1(new_n524), .B2(G110), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(new_n210), .A3(new_n231), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT77), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G110), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT76), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n529), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n530), .B2(new_n524), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n532), .B(new_n232), .C1(new_n519), .C2(new_n520), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT78), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n528), .A2(KEYINPUT78), .A3(new_n533), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n515), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n515), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n511), .B1(new_n541), .B2(new_n267), .ZN(new_n542));
  INV_X1    g356(.A(new_n537), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT78), .B1(new_n528), .B2(new_n533), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n514), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n539), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n546), .A2(G902), .A3(new_n510), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n508), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n546), .A2(KEYINPUT80), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(KEYINPUT80), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n508), .A2(G902), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G472), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n195), .A2(G210), .A3(new_n188), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT26), .B(G101), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n407), .A2(KEYINPUT67), .A3(G134), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n406), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT67), .B1(new_n407), .B2(G134), .ZN(new_n563));
  OAI21_X1  g377(.A(G131), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n564), .A2(new_n411), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n349), .A2(new_n351), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n462), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n338), .A2(KEYINPUT65), .A3(new_n380), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT65), .B1(new_n338), .B2(new_n380), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n385), .B(new_n412), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n571), .A2(KEYINPUT28), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(KEYINPUT28), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(KEYINPUT66), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT66), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n384), .A2(new_n576), .A3(new_n385), .A4(new_n412), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n347), .A2(new_n565), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n462), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n560), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT30), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n566), .A2(KEYINPUT30), .A3(new_n570), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n462), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT31), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n571), .A4(new_n560), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n588), .A2(KEYINPUT75), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(KEYINPUT75), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n582), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n586), .A2(new_n571), .A3(new_n560), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n592), .A2(KEYINPUT74), .A3(KEYINPUT31), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT74), .B1(new_n592), .B2(KEYINPUT31), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n554), .B(new_n267), .C1(new_n591), .C2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT32), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n571), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n570), .A2(KEYINPUT66), .B1(new_n347), .B2(new_n565), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT30), .B1(new_n600), .B2(new_n577), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n566), .A2(KEYINPUT30), .A3(new_n570), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n599), .B1(new_n603), .B2(new_n462), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT75), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n587), .A4(new_n560), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n588), .A2(KEYINPUT75), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n581), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n592), .A2(KEYINPUT31), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT74), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n592), .A2(KEYINPUT74), .A3(KEYINPUT31), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n554), .A2(new_n267), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n597), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n567), .B1(new_n566), .B2(new_n570), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n572), .B2(new_n573), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT29), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n559), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(G902), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n574), .A2(new_n560), .A3(new_n580), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n619), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n604), .A2(new_n560), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n614), .A2(new_n616), .B1(G472), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n553), .B1(new_n598), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n325), .A2(new_n507), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  AND3_X1   g443(.A1(new_n493), .A2(new_n501), .A3(new_n449), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n447), .B(new_n324), .C1(new_n630), .C2(new_n502), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n553), .A2(new_n631), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n632), .A2(new_n446), .A3(new_n506), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n267), .B1(new_n591), .B2(new_n595), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(G472), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n635), .A2(new_n596), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n296), .A2(new_n300), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n638), .A2(KEYINPUT102), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(KEYINPUT102), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n302), .B(KEYINPUT101), .Z(new_n643));
  AOI22_X1  g457(.A1(new_n642), .A2(new_n643), .B1(new_n641), .B2(new_n308), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n310), .A2(G902), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT103), .B(G478), .Z(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n644), .A2(new_n645), .B1(new_n309), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n266), .B2(new_n274), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n637), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT34), .B(G104), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  NOR2_X1   g467(.A1(new_n251), .A2(new_n252), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n264), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n257), .A2(new_n262), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n315), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n656), .A2(new_n274), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n633), .A2(new_n636), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT35), .B(G107), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NOR2_X1   g475(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n534), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n551), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n548), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n635), .A2(new_n596), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n325), .A2(new_n507), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n320), .B1(new_n321), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n656), .A2(new_n274), .A3(new_n657), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n510), .B1(new_n546), .B2(G902), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n541), .A2(new_n267), .A3(new_n511), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n677), .A2(new_n508), .B1(new_n551), .B2(new_n663), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n598), .B2(new_n626), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n674), .A2(new_n507), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  OAI21_X1  g495(.A(new_n616), .B1(new_n591), .B2(new_n595), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n559), .B1(new_n599), .B2(new_n617), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT104), .Z(new_n684));
  INV_X1    g498(.A(new_n592), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n267), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(G472), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n598), .A2(new_n682), .A3(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n446), .A2(new_n506), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n671), .B(KEYINPUT39), .Z(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT40), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n266), .A2(new_n274), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n630), .A2(new_n502), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n695), .A2(KEYINPUT38), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(KEYINPUT38), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n696), .A2(new_n447), .A3(new_n678), .A4(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n694), .A2(new_n698), .A3(new_n315), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT40), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n689), .A2(new_n700), .A3(new_n690), .ZN(new_n701));
  AND4_X1   g515(.A1(new_n688), .A2(new_n692), .A3(new_n699), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n191), .ZN(G45));
  AOI211_X1 g517(.A(new_n648), .B(new_n671), .C1(new_n266), .C2(new_n274), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n507), .A3(new_n679), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  INV_X1    g520(.A(new_n631), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n649), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n426), .B1(new_n425), .B2(new_n420), .ZN(new_n711));
  AND4_X1   g525(.A1(new_n426), .A2(new_n403), .A3(new_n412), .A4(new_n420), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n430), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n436), .B1(new_n713), .B2(new_n329), .ZN(new_n714));
  OAI21_X1  g528(.A(G469), .B1(new_n714), .B2(G902), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n715), .A2(new_n506), .A3(new_n437), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n709), .A2(new_n710), .A3(new_n627), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n627), .A2(new_n716), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT105), .B1(new_n718), .B2(new_n708), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  NAND4_X1  g536(.A1(new_n658), .A2(new_n627), .A3(new_n707), .A4(new_n716), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G116), .ZN(G18));
  NAND4_X1  g538(.A1(new_n715), .A2(new_n505), .A3(new_n506), .A4(new_n437), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n325), .A2(new_n679), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  AOI21_X1  g542(.A(G902), .B1(new_n608), .B2(new_n613), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n554), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n606), .A2(new_n607), .ZN(new_n731));
  INV_X1    g545(.A(new_n618), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n732), .A2(new_n559), .B1(new_n592), .B2(KEYINPUT31), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n615), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n730), .A2(new_n553), .A3(new_n734), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n506), .A2(new_n715), .A3(new_n437), .A4(new_n324), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n315), .B1(new_n266), .B2(new_n274), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n735), .A2(new_n736), .A3(new_n737), .A4(new_n505), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  INV_X1    g553(.A(new_n734), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n665), .B(new_n740), .C1(new_n729), .C2(new_n554), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n725), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n704), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n598), .A2(new_n626), .ZN(new_n746));
  INV_X1    g560(.A(new_n553), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n443), .A2(KEYINPUT106), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n438), .B1(new_n422), .B2(new_n427), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n441), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n751), .A3(G469), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n748), .A2(new_n437), .A3(new_n752), .A4(new_n445), .ZN(new_n753));
  INV_X1    g567(.A(new_n506), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n630), .A2(new_n502), .A3(new_n448), .A4(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n746), .A2(new_n747), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n649), .A2(new_n672), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n745), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n753), .A2(new_n755), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n704), .A2(new_n759), .A3(KEYINPUT42), .A4(new_n627), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n756), .B2(new_n673), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n674), .A2(new_n759), .A3(KEYINPUT107), .A4(new_n627), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT108), .B(G134), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G36));
  INV_X1    g582(.A(new_n648), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n694), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT43), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n693), .A2(KEYINPUT43), .A3(new_n648), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n636), .A2(new_n678), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n750), .A2(KEYINPUT45), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n750), .A2(KEYINPUT45), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(G469), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n445), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n713), .A2(new_n329), .ZN(new_n782));
  INV_X1    g596(.A(new_n436), .ZN(new_n783));
  AOI21_X1  g597(.A(G902), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI22_X1  g598(.A1(new_n780), .A2(new_n781), .B1(new_n326), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n445), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n754), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n695), .A2(new_n447), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n787), .A2(new_n690), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n774), .A2(new_n775), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n776), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  XOR2_X1   g606(.A(KEYINPUT109), .B(G137), .Z(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(G39));
  NAND2_X1  g608(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n757), .A2(new_n746), .A3(new_n747), .A4(new_n788), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n798));
  OAI211_X1 g612(.A(new_n796), .B(new_n797), .C1(new_n787), .C2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  NAND3_X1  g614(.A1(new_n771), .A2(new_n320), .A3(new_n772), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT113), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n771), .A2(new_n803), .A3(new_n320), .A4(new_n772), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n726), .A3(new_n735), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n716), .A2(new_n320), .A3(new_n747), .A4(new_n789), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n688), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(KEYINPUT117), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(KEYINPUT117), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n806), .B(new_n317), .C1(new_n650), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n716), .A2(new_n789), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n802), .B2(new_n804), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n627), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(KEYINPUT48), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(KEYINPUT48), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n812), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n696), .A2(new_n697), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n716), .A2(new_n448), .ZN(new_n821));
  OAI221_X1 g635(.A(new_n820), .B1(KEYINPUT116), .B2(KEYINPUT50), .C1(new_n821), .C2(KEYINPUT115), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(KEYINPUT115), .B2(new_n821), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n805), .A2(new_n735), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n827), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n805), .A2(new_n735), .A3(new_n829), .A4(new_n823), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n805), .A2(new_n735), .A3(new_n789), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n796), .B1(new_n787), .B2(new_n798), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n715), .A2(new_n437), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n754), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n832), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n741), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n814), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n693), .A2(new_n769), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n839), .B(new_n840), .C1(new_n811), .C2(new_n842), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n741), .B(new_n813), .C1(new_n802), .C2(new_n804), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n811), .A2(new_n842), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT118), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n819), .B1(new_n837), .B2(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT51), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n787), .A2(new_n795), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n787), .A2(new_n798), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT114), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n796), .B(new_n853), .C1(new_n787), .C2(new_n798), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n852), .A2(new_n835), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n849), .B1(new_n832), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n831), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n818), .B1(new_n848), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n266), .A2(new_n274), .A3(new_n657), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n633), .B(new_n636), .C1(new_n860), .C2(new_n649), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n325), .B(new_n507), .C1(new_n627), .C2(new_n666), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n723), .A2(new_n727), .A3(new_n738), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT111), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n865), .A2(new_n720), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n312), .A2(new_n314), .A3(new_n671), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n870), .A2(new_n695), .A3(new_n447), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n446), .A2(new_n871), .A3(new_n506), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n656), .A2(new_n274), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n873), .A3(new_n679), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT112), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT112), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n872), .A2(new_n876), .A3(new_n873), .A4(new_n679), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n704), .A2(new_n759), .A3(new_n838), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n761), .A3(new_n766), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n869), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n678), .A2(new_n506), .A3(new_n672), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n444), .B1(new_n784), .B2(new_n326), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n751), .B1(new_n750), .B2(G469), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n749), .A2(new_n441), .A3(KEYINPUT106), .A4(new_n326), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n882), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n505), .A3(new_n688), .A4(new_n737), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n705), .A2(new_n680), .A3(new_n888), .A4(new_n743), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT52), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT32), .B1(new_n729), .B2(new_n554), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n625), .A2(G472), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n682), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n665), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n446), .A2(new_n505), .A3(new_n506), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI22_X1  g710(.A1(new_n896), .A2(new_n674), .B1(new_n704), .B2(new_n742), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT52), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n898), .A3(new_n705), .A4(new_n888), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n890), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT53), .B1(new_n881), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT53), .ZN(new_n903));
  NOR4_X1   g717(.A1(new_n869), .A2(new_n900), .A3(new_n880), .A4(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n859), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n878), .A2(new_n761), .A3(new_n879), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT111), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT111), .B1(new_n861), .B2(new_n862), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n866), .B1(new_n717), .B2(new_n719), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n906), .A2(new_n909), .A3(new_n766), .A4(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n903), .B1(new_n911), .B2(new_n900), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n881), .A2(KEYINPUT53), .A3(new_n901), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(KEYINPUT54), .A3(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n905), .A2(new_n914), .ZN(new_n915));
  OAI22_X1  g729(.A1(new_n858), .A2(new_n915), .B1(G952), .B2(G953), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n820), .A2(new_n447), .A3(new_n506), .A4(new_n747), .ZN(new_n917));
  INV_X1    g731(.A(new_n834), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(KEYINPUT49), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(KEYINPUT49), .B2(new_n918), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n920), .A2(new_n688), .A3(new_n770), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n916), .A2(new_n921), .ZN(G75));
  AOI21_X1  g736(.A(new_n267), .B1(new_n912), .B2(new_n913), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(G210), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT56), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n497), .A2(new_n500), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT119), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(new_n498), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n924), .A2(new_n925), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n924), .B2(new_n925), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n195), .A2(G952), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(G51));
  XNOR2_X1  g747(.A(new_n444), .B(KEYINPUT57), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n905), .A2(new_n914), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n714), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI211_X1 g751(.A(new_n267), .B(new_n779), .C1(new_n912), .C2(new_n913), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n941));
  INV_X1    g755(.A(new_n932), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n938), .B1(new_n935), .B2(new_n936), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT120), .B1(new_n944), .B2(new_n932), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(G54));
  NAND3_X1  g760(.A1(new_n923), .A2(KEYINPUT58), .A3(G475), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n252), .B2(new_n251), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n923), .A2(KEYINPUT58), .A3(G475), .A4(new_n654), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n948), .A2(new_n942), .A3(new_n949), .ZN(G60));
  NAND2_X1  g764(.A1(G478), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT59), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n905), .A2(new_n914), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n644), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n955), .A2(new_n956), .A3(new_n932), .ZN(G63));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT121), .Z(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT60), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n912), .B2(new_n913), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n663), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n549), .A2(new_n550), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n962), .B(new_n942), .C1(new_n963), .C2(new_n961), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT122), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT61), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n964), .B(new_n966), .ZN(G66));
  INV_X1    g781(.A(new_n322), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n316), .B1(new_n968), .B2(G224), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n869), .B2(new_n195), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n927), .B1(G898), .B2(new_n195), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT123), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n970), .B(new_n972), .ZN(G69));
  XOR2_X1   g787(.A(new_n603), .B(new_n247), .Z(new_n974));
  INV_X1    g788(.A(KEYINPUT124), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n897), .A2(new_n705), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n977));
  OR3_X1    g791(.A1(new_n702), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n702), .B2(new_n976), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n691), .A2(new_n788), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n981), .B(new_n627), .C1(new_n649), .C2(new_n860), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n792), .A2(new_n799), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n975), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n792), .A2(new_n799), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n978), .A2(new_n979), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT124), .A4(new_n982), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n974), .B1(new_n988), .B2(new_n195), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n627), .A2(new_n737), .A3(new_n505), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n787), .A2(new_n690), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n992), .A2(new_n761), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n976), .B1(new_n764), .B2(new_n765), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n792), .A2(new_n993), .A3(new_n799), .A4(new_n994), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n995), .A2(new_n194), .A3(new_n193), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n974), .B1(new_n670), .B2(new_n195), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OR3_X1    g812(.A1(new_n989), .A2(new_n990), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n990), .B1(new_n989), .B2(new_n998), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(G72));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  OAI221_X1 g817(.A(new_n1003), .B1(new_n685), .B2(new_n624), .C1(new_n902), .C2(new_n904), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1003), .B(KEYINPUT125), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(new_n995), .B2(new_n869), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n604), .A2(new_n559), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1005), .B1(new_n1009), .B2(new_n942), .ZN(new_n1010));
  AOI211_X1 g824(.A(KEYINPUT127), .B(new_n932), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1004), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n869), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n984), .A2(new_n987), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n1006), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n604), .A2(new_n559), .ZN(new_n1016));
  AOI21_X1  g830(.A(KEYINPUT126), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT126), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1016), .ZN(new_n1019));
  AOI211_X1 g833(.A(new_n1018), .B(new_n1019), .C1(new_n1014), .C2(new_n1006), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n1012), .A2(new_n1017), .A3(new_n1020), .ZN(G57));
endmodule


