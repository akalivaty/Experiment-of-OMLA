//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT64), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n206));
  INV_X1    g005(.A(G127gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(G134gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G127gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G113gat), .ZN(new_n212));
  INV_X1    g011(.A(G120gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n215));
  NAND2_X1  g014(.A1(G113gat), .A2(G120gat), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n209), .A2(G127gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n207), .A2(G134gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT68), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n211), .A2(new_n217), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n223), .A2(KEYINPUT68), .A3(new_n218), .A4(new_n219), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n222), .B1(new_n221), .B2(new_n224), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228));
  NOR2_X1   g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  AND2_X1   g028(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n231), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G169gat), .ZN(new_n240));
  INV_X1    g039(.A(G176gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(KEYINPUT23), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT23), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(G169gat), .B2(G176gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT25), .B1(new_n239), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(G183gat), .B2(G190gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(new_n237), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n252));
  NOR3_X1   g051(.A1(new_n251), .A2(new_n252), .A3(new_n246), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n228), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n234), .B(new_n249), .C1(G183gat), .C2(G190gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n247), .A2(KEYINPUT25), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT65), .B1(new_n232), .B2(new_n233), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n246), .B1(new_n258), .B2(new_n238), .ZN(new_n259));
  OAI211_X1 g058(.A(KEYINPUT66), .B(new_n256), .C1(new_n259), .C2(KEYINPUT25), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT26), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n262), .A2(KEYINPUT26), .ZN(new_n264));
  INV_X1    g063(.A(new_n245), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n263), .B(new_n232), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n267));
  INV_X1    g066(.A(G183gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT27), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT67), .ZN(new_n270));
  INV_X1    g069(.A(G190gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT27), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G183gat), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT67), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n267), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n269), .A2(new_n274), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(KEYINPUT28), .A3(new_n271), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n266), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n227), .B1(new_n261), .B2(new_n280), .ZN(new_n281));
  AOI211_X1 g080(.A(new_n279), .B(new_n225), .C1(new_n254), .C2(new_n260), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n205), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT33), .ZN(new_n284));
  XNOR2_X1  g083(.A(G15gat), .B(G43gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(G71gat), .B(G99gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n283), .B(KEYINPUT32), .C1(new_n284), .C2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n283), .B2(KEYINPUT32), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n283), .A2(new_n284), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n290), .B1(new_n289), .B2(new_n291), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n288), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n281), .A2(new_n282), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n202), .B2(new_n203), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT34), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n205), .A2(KEYINPUT34), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n302));
  INV_X1    g101(.A(new_n300), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n303), .B(new_n288), .C1(new_n292), .C2(new_n293), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n301), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT36), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n294), .A2(KEYINPUT72), .A3(new_n300), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n305), .A2(KEYINPUT73), .A3(new_n306), .A4(new_n307), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n294), .A2(KEYINPUT71), .A3(new_n300), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n312), .A2(new_n304), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n301), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(KEYINPUT36), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n310), .A2(new_n311), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G197gat), .B(G204gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT22), .ZN(new_n319));
  INV_X1    g118(.A(G211gat), .ZN(new_n320));
  INV_X1    g119(.A(G218gat), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G211gat), .B(G218gat), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n323), .B(new_n324), .Z(new_n325));
  XOR2_X1   g124(.A(G155gat), .B(G162gat), .Z(new_n326));
  INV_X1    g125(.A(KEYINPUT78), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G148gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT77), .B1(new_n329), .B2(G141gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n331));
  INV_X1    g130(.A(G141gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n332), .A3(G148gat), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n330), .B(new_n333), .C1(new_n332), .C2(G148gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT2), .ZN(new_n336));
  XNOR2_X1  g135(.A(G155gat), .B(G162gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT78), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n328), .A2(new_n334), .A3(new_n336), .A4(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G141gat), .B(G148gat), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n326), .B1(KEYINPUT2), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n325), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(KEYINPUT81), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT81), .ZN(new_n348));
  AOI211_X1 g147(.A(new_n348), .B(new_n325), .C1(new_n344), .C2(new_n345), .ZN(new_n349));
  INV_X1    g148(.A(G228gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(new_n203), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT3), .B1(new_n325), .B2(new_n345), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(new_n342), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n347), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n324), .A2(new_n318), .A3(new_n355), .A4(new_n322), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n345), .B(new_n356), .C1(new_n325), .C2(new_n355), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n342), .B1(new_n357), .B2(new_n343), .ZN(new_n358));
  OAI22_X1  g157(.A1(new_n358), .A2(new_n346), .B1(new_n350), .B2(new_n203), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(G22gat), .B1(new_n354), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G22gat), .ZN(new_n362));
  OAI221_X1 g161(.A(new_n351), .B1(new_n342), .B2(new_n352), .C1(new_n346), .C2(KEYINPUT81), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n362), .B(new_n359), .C1(new_n363), .C2(new_n349), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT82), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT83), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT31), .B(G50gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n365), .B2(new_n366), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT83), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n361), .A2(KEYINPUT82), .A3(new_n364), .A4(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n367), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n372), .B1(new_n367), .B2(new_n374), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT6), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n221), .A2(new_n224), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n339), .A2(new_n341), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n381), .B2(KEYINPUT3), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n344), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n342), .A2(new_n380), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n342), .A2(KEYINPUT4), .A3(new_n380), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n383), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT5), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n381), .A2(new_n224), .A3(new_n221), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n387), .B1(new_n384), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n389), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G1gat), .B(G29gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(KEYINPUT0), .ZN(new_n396));
  XNOR2_X1  g195(.A(G57gat), .B(G85gat), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n396), .B(new_n397), .Z(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n391), .A2(new_n394), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n391), .B2(new_n394), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n379), .B(new_n400), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n401), .A2(new_n402), .ZN(new_n404));
  OAI22_X1  g203(.A1(new_n403), .A2(new_n404), .B1(new_n379), .B2(new_n400), .ZN(new_n405));
  INV_X1    g204(.A(new_n325), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n256), .B1(new_n259), .B2(KEYINPUT25), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n280), .A2(KEYINPUT74), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT74), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n248), .A2(new_n253), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(new_n279), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n408), .A2(new_n411), .A3(new_n345), .ZN(new_n412));
  NAND2_X1  g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n261), .A2(new_n280), .ZN(new_n416));
  INV_X1    g215(.A(new_n413), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n412), .A2(new_n415), .A3(new_n413), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n406), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n416), .A2(new_n345), .A3(new_n413), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n408), .A2(new_n411), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n422), .B1(new_n423), .B2(new_n413), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(new_n325), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT76), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n429), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n421), .A2(new_n425), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT30), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n433), .A2(KEYINPUT30), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n405), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n378), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n317), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n317), .A2(KEYINPUT84), .A3(new_n437), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT37), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n419), .A2(new_n420), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n406), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n445), .B(KEYINPUT37), .C1(new_n406), .C2(new_n424), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT87), .B(KEYINPUT38), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n430), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n443), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n449), .B(KEYINPUT88), .Z(new_n450));
  INV_X1    g249(.A(new_n443), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n432), .B1(new_n426), .B2(new_n442), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n447), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n405), .A2(new_n433), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n435), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n383), .A2(new_n386), .A3(new_n388), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(G225gat), .A3(G233gat), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n458), .A2(KEYINPUT39), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n384), .A2(new_n387), .A3(new_n392), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT39), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n461), .A2(KEYINPUT85), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(KEYINPUT85), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n458), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n459), .A2(new_n464), .A3(new_n398), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT40), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n467), .A2(new_n400), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT40), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n469), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n466), .A2(KEYINPUT86), .A3(KEYINPUT40), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n456), .B(new_n468), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n377), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n440), .A2(new_n441), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT35), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n436), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n405), .A2(new_n434), .A3(KEYINPUT89), .A4(new_n435), .ZN(new_n479));
  AND4_X1   g278(.A1(new_n476), .A2(new_n478), .A3(new_n377), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n305), .A2(new_n307), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n436), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n377), .A2(new_n483), .A3(new_n315), .A4(new_n313), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n475), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(G29gat), .A2(G36gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT14), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G36gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT91), .B(G29gat), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT15), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n494), .ZN(new_n496));
  XNOR2_X1  g295(.A(G43gat), .B(G50gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OR3_X1    g297(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT17), .ZN(new_n501));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT16), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n502), .B1(new_n503), .B2(G1gat), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(G1gat), .B2(new_n502), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(G8gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT92), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n501), .A2(new_n507), .B1(new_n506), .B2(new_n500), .ZN(new_n508));
  NAND2_X1  g307(.A1(G229gat), .A2(G233gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT93), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT18), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n508), .A2(KEYINPUT18), .A3(new_n511), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT94), .B1(new_n500), .B2(new_n506), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n506), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n510), .B(KEYINPUT13), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n514), .A2(new_n515), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT90), .B(G197gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(KEYINPUT11), .B(G169gat), .Z(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT12), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n514), .A2(new_n515), .A3(new_n520), .A4(new_n527), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(G71gat), .A2(G78gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT95), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT9), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G64gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n538), .A2(G57gat), .ZN(new_n539));
  INV_X1    g338(.A(G57gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n540), .A2(G64gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n539), .A2(KEYINPUT96), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n539), .A2(KEYINPUT96), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n544), .B(new_n545), .C1(new_n540), .C2(G64gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n533), .B1(new_n532), .B2(new_n536), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n549), .A2(KEYINPUT21), .ZN(new_n550));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G127gat), .B(G155gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT20), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n552), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G183gat), .B(G211gat), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n506), .B1(new_n549), .B2(KEYINPUT21), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n558), .B(KEYINPUT98), .Z(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n556), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n555), .B(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n561), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT101), .B(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G99gat), .ZN(new_n571));
  INV_X1    g370(.A(G106gat), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT8), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT102), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G85gat), .A2(G92gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT7), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G99gat), .B(G106gat), .Z(new_n580));
  OR2_X1    g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n501), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n581), .A2(new_n582), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n500), .ZN(new_n586));
  NAND3_X1  g385(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT103), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n584), .A2(new_n586), .A3(new_n587), .A4(new_n589), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT99), .ZN(new_n595));
  XOR2_X1   g394(.A(G134gat), .B(G162gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT100), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n591), .A2(new_n592), .A3(new_n593), .A4(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n591), .A2(new_n593), .A3(new_n598), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT103), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n597), .B1(new_n591), .B2(new_n593), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n567), .A2(KEYINPUT104), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT104), .B1(new_n567), .B2(new_n603), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n585), .A2(new_n549), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(KEYINPUT105), .A3(KEYINPUT10), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g410(.A(new_n549), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n583), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT105), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G230gat), .A2(G233gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n583), .A2(new_n612), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n610), .A2(new_n615), .A3(new_n616), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n609), .A2(new_n617), .ZN(new_n619));
  INV_X1    g418(.A(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT107), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT106), .ZN(new_n625));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n622), .A2(KEYINPUT107), .A3(new_n627), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n608), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n487), .A2(new_n531), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT108), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n487), .A2(KEYINPUT108), .A3(new_n531), .A4(new_n632), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n405), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G1gat), .ZN(G1324gat));
  INV_X1    g439(.A(new_n456), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT16), .B(G8gat), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AOI211_X1 g442(.A(new_n641), .B(new_n643), .C1(new_n635), .C2(new_n636), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n644), .A2(KEYINPUT42), .ZN(new_n645));
  INV_X1    g444(.A(G8gat), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n646), .B1(new_n637), .B2(new_n456), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT42), .B1(new_n647), .B2(new_n644), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(G1325gat));
  INV_X1    g448(.A(new_n317), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(G15gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT110), .Z(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n635), .B2(new_n636), .ZN(new_n653));
  INV_X1    g452(.A(new_n481), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n654), .B1(new_n635), .B2(new_n636), .ZN(new_n655));
  OR3_X1    g454(.A1(new_n655), .A2(KEYINPUT109), .A3(G15gat), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT109), .B1(new_n655), .B2(G15gat), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(G1326gat));
  NAND2_X1  g457(.A1(new_n637), .A2(new_n378), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT43), .B(G22gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  AOI21_X1  g460(.A(new_n603), .B1(new_n475), .B2(new_n486), .ZN(new_n662));
  INV_X1    g461(.A(new_n531), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n567), .A2(new_n663), .A3(new_n631), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n665), .A2(new_n638), .A3(new_n492), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT45), .ZN(new_n667));
  INV_X1    g466(.A(new_n603), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n317), .A2(KEYINPUT84), .A3(new_n437), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT84), .B1(new_n317), .B2(new_n437), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n455), .A2(new_n377), .A3(new_n473), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n480), .A2(new_n481), .B1(new_n484), .B2(KEYINPUT35), .ZN(new_n673));
  OAI211_X1 g472(.A(KEYINPUT44), .B(new_n668), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  INV_X1    g474(.A(new_n438), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n673), .B1(new_n676), .B2(new_n474), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n677), .B2(new_n603), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n674), .A2(new_n664), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT111), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n674), .A2(new_n678), .A3(KEYINPUT111), .A4(new_n664), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n681), .A2(new_n638), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n667), .B1(new_n492), .B2(new_n683), .ZN(G1328gat));
  NAND3_X1  g483(.A1(new_n665), .A2(new_n491), .A3(new_n456), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT46), .Z(new_n686));
  NAND3_X1  g485(.A1(new_n681), .A2(new_n456), .A3(new_n682), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G36gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(G1329gat));
  INV_X1    g488(.A(KEYINPUT113), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n679), .B2(new_n317), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n474), .A2(new_n437), .A3(new_n317), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n486), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT44), .B1(new_n693), .B2(new_n668), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n662), .B2(KEYINPUT44), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n695), .A2(KEYINPUT113), .A3(new_n650), .A4(new_n664), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n691), .A2(new_n696), .A3(G43gat), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n654), .A2(G43gat), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n662), .A2(new_n664), .A3(new_n698), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n699), .A2(KEYINPUT47), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(KEYINPUT112), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT112), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n662), .A2(new_n703), .A3(new_n664), .A4(new_n698), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n681), .A2(new_n650), .A3(new_n682), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(G43gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n701), .B1(new_n707), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g507(.A(G50gat), .B1(new_n679), .B2(new_n377), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n377), .A2(G50gat), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT114), .Z(new_n711));
  NAND2_X1  g510(.A1(new_n665), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(KEYINPUT48), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n712), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n681), .A2(new_n378), .A3(new_n682), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(G50gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n713), .B1(new_n716), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g516(.A(new_n631), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n608), .A2(new_n531), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n693), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n405), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(new_n540), .ZN(G1332gat));
  INV_X1    g521(.A(KEYINPUT115), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n720), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n456), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT49), .B(G64gat), .Z(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n725), .B2(new_n727), .ZN(G1333gat));
  NAND3_X1  g527(.A1(new_n724), .A2(G71gat), .A3(new_n650), .ZN(new_n729));
  INV_X1    g528(.A(G71gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n720), .B2(new_n654), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g532(.A1(new_n724), .A2(new_n378), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT116), .B(G78gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1335gat));
  NOR3_X1   g535(.A1(new_n718), .A2(new_n531), .A3(new_n567), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n695), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n738), .A2(new_n638), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n603), .B1(new_n486), .B2(new_n692), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n567), .A2(new_n531), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n740), .A2(KEYINPUT51), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT51), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n631), .A2(new_n638), .A3(new_n568), .ZN(new_n745));
  OAI22_X1  g544(.A1(new_n739), .A2(new_n568), .B1(new_n744), .B2(new_n745), .ZN(G1336gat));
  NAND3_X1  g545(.A1(new_n695), .A2(new_n456), .A3(new_n737), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(G92gat), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n718), .A2(G92gat), .A3(new_n641), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n742), .B2(new_n743), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT117), .ZN(new_n751));
  INV_X1    g550(.A(new_n749), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n693), .A2(new_n668), .A3(new_n741), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n740), .A2(KEYINPUT51), .A3(new_n741), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n751), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT52), .B1(new_n748), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n747), .A2(G92gat), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT52), .B1(new_n757), .B2(KEYINPUT118), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n762), .B(new_n763), .C1(KEYINPUT118), .C2(new_n757), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(G1337gat));
  AND2_X1   g564(.A1(new_n738), .A2(new_n650), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n481), .A2(new_n631), .A3(new_n571), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n766), .A2(new_n571), .B1(new_n744), .B2(new_n767), .ZN(G1338gat));
  NAND3_X1  g567(.A1(new_n695), .A2(new_n378), .A3(new_n737), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n718), .A2(new_n377), .A3(G106gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n742), .B2(new_n743), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT53), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n770), .A2(new_n775), .A3(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(G1339gat));
  INV_X1    g576(.A(new_n567), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT121), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n627), .B1(new_n618), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n610), .A2(new_n615), .A3(new_n617), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n620), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(KEYINPUT54), .A3(new_n618), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n779), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n622), .A2(new_n627), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n787), .B2(new_n788), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n508), .A2(new_n511), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n518), .A2(new_n519), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n526), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n530), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n603), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n783), .A2(new_n786), .A3(KEYINPUT121), .A4(KEYINPUT55), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n789), .A2(new_n791), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT122), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n785), .A2(KEYINPUT54), .A3(new_n618), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n788), .B1(new_n801), .B2(new_n782), .ZN(new_n802));
  INV_X1    g601(.A(new_n790), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n802), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n804), .A2(KEYINPUT122), .A3(new_n789), .A4(new_n796), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n789), .A2(new_n791), .A3(new_n531), .A4(new_n797), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n631), .A2(new_n530), .A3(new_n794), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n668), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n778), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n607), .A2(KEYINPUT119), .A3(new_n663), .A4(new_n718), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n567), .A2(new_n603), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT104), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n814), .A2(new_n718), .A3(new_n663), .A4(new_n604), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n810), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n377), .A2(new_n315), .A3(new_n313), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n456), .A2(new_n405), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n531), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n378), .A2(new_n654), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n819), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n822), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n663), .A2(new_n212), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n826), .B1(new_n829), .B2(new_n830), .ZN(G1340gat));
  AOI21_X1  g630(.A(G120gat), .B1(new_n825), .B2(new_n631), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n718), .A2(new_n213), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n829), .B2(new_n833), .ZN(G1341gat));
  INV_X1    g633(.A(new_n829), .ZN(new_n835));
  OAI21_X1  g634(.A(G127gat), .B1(new_n835), .B2(new_n778), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n825), .A2(new_n207), .A3(new_n567), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1342gat));
  NOR3_X1   g637(.A1(new_n824), .A2(G134gat), .A3(new_n603), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT56), .ZN(new_n840));
  OAI21_X1  g639(.A(G134gat), .B1(new_n835), .B2(new_n603), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1343gat));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(KEYINPUT58), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n650), .A2(new_n822), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n377), .B1(new_n810), .B2(new_n818), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(KEYINPUT57), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  AOI211_X1 g648(.A(new_n849), .B(new_n377), .C1(new_n810), .C2(new_n818), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n531), .B(new_n846), .C1(new_n848), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(G141gat), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n847), .A2(new_n332), .A3(new_n531), .A4(new_n846), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n843), .A2(KEYINPUT58), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n845), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  AOI211_X1 g656(.A(new_n844), .B(new_n855), .C1(new_n851), .C2(G141gat), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(G1344gat));
  INV_X1    g658(.A(new_n847), .ZN(new_n860));
  INV_X1    g659(.A(new_n846), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n329), .A3(new_n631), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(G148gat), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n848), .A2(new_n850), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n861), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n867), .B2(new_n631), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n847), .A2(KEYINPUT57), .ZN(new_n869));
  INV_X1    g668(.A(new_n798), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n778), .B1(new_n809), .B2(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n815), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n849), .B1(new_n872), .B2(new_n377), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g673(.A(new_n846), .B(KEYINPUT124), .Z(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n631), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n864), .B1(new_n876), .B2(G148gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n863), .B1(new_n868), .B2(new_n877), .ZN(G1345gat));
  AOI21_X1  g677(.A(G155gat), .B1(new_n862), .B2(new_n567), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n567), .A2(G155gat), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT125), .Z(new_n881));
  AOI21_X1  g680(.A(new_n879), .B1(new_n867), .B2(new_n881), .ZN(G1346gat));
  AOI21_X1  g681(.A(G162gat), .B1(new_n862), .B2(new_n668), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n668), .A2(G162gat), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n867), .B2(new_n885), .ZN(G1347gat));
  INV_X1    g685(.A(new_n828), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n641), .A2(new_n638), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(new_n240), .A3(new_n663), .ZN(new_n890));
  INV_X1    g689(.A(new_n888), .ZN(new_n891));
  AOI211_X1 g690(.A(new_n820), .B(new_n891), .C1(new_n810), .C2(new_n818), .ZN(new_n892));
  AOI21_X1  g691(.A(G169gat), .B1(new_n892), .B2(new_n531), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n890), .A2(new_n893), .ZN(G1348gat));
  OAI21_X1  g693(.A(G176gat), .B1(new_n889), .B2(new_n718), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(new_n241), .A3(new_n631), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1349gat));
  OAI21_X1  g696(.A(G183gat), .B1(new_n889), .B2(new_n778), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n892), .A2(new_n277), .A3(new_n567), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT60), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n898), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n887), .A2(new_n668), .A3(new_n888), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G190gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT126), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n908), .A3(G190gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n909), .A3(KEYINPUT61), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n892), .A2(new_n271), .A3(new_n668), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n908), .B1(new_n905), .B2(G190gat), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n910), .A2(new_n914), .ZN(G1351gat));
  NOR2_X1   g714(.A1(new_n650), .A2(new_n891), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n860), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(G197gat), .B1(new_n918), .B2(new_n531), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n869), .B2(new_n873), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n531), .A2(G197gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  INV_X1    g721(.A(G204gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n918), .A2(new_n923), .A3(new_n631), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(KEYINPUT62), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(KEYINPUT62), .ZN(new_n926));
  AOI211_X1 g725(.A(new_n718), .B(new_n917), .C1(new_n869), .C2(new_n873), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n925), .B(new_n926), .C1(new_n923), .C2(new_n927), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n918), .A2(new_n320), .A3(new_n567), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n920), .A2(new_n567), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n931), .A2(KEYINPUT127), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n320), .B1(KEYINPUT127), .B2(new_n931), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n930), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n929), .B1(new_n934), .B2(new_n935), .ZN(G1354gat));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n321), .A3(new_n668), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n920), .A2(new_n668), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n321), .ZN(G1355gat));
endmodule


