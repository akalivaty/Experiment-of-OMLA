

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755;

  INV_X1 U383 ( .A(KEYINPUT64), .ZN(n444) );
  NOR2_X2 U384 ( .A1(n374), .A2(n630), .ZN(n643) );
  XNOR2_X2 U385 ( .A(n575), .B(n449), .ZN(n611) );
  XNOR2_X2 U386 ( .A(n448), .B(G469), .ZN(n575) );
  NOR2_X1 U387 ( .A1(n717), .A2(n726), .ZN(n718) );
  AND2_X1 U388 ( .A1(n394), .A2(n401), .ZN(n400) );
  AND2_X1 U389 ( .A1(n397), .A2(n403), .ZN(n396) );
  AND2_X1 U390 ( .A1(n574), .A2(n367), .ZN(n397) );
  XNOR2_X1 U391 ( .A(n557), .B(n556), .ZN(n561) );
  OR2_X1 U392 ( .A1(n598), .A2(n554), .ZN(n555) );
  OR2_X1 U393 ( .A1(n567), .A2(n568), .ZN(n554) );
  NAND2_X1 U394 ( .A1(n550), .A2(n627), .ZN(n606) );
  XNOR2_X1 U395 ( .A(n516), .B(n369), .ZN(n550) );
  NOR2_X1 U396 ( .A1(n713), .A2(G902), .ZN(n448) );
  XNOR2_X1 U397 ( .A(n462), .B(n452), .ZN(n739) );
  XNOR2_X1 U398 ( .A(KEYINPUT22), .B(KEYINPUT74), .ZN(n556) );
  XNOR2_X1 U399 ( .A(G128), .B(G143), .ZN(n509) );
  XNOR2_X1 U400 ( .A(n458), .B(n457), .ZN(n600) );
  NAND2_X1 U401 ( .A1(n754), .A2(n688), .ZN(n417) );
  XNOR2_X1 U402 ( .A(n409), .B(G125), .ZN(n506) );
  INV_X1 U403 ( .A(G146), .ZN(n409) );
  XNOR2_X1 U404 ( .A(G137), .B(KEYINPUT69), .ZN(n452) );
  AND2_X1 U405 ( .A1(n588), .A2(n371), .ZN(n404) );
  NAND2_X1 U406 ( .A1(n413), .A2(n410), .ZN(n403) );
  NAND2_X1 U407 ( .A1(n412), .A2(n365), .ZN(n410) );
  AND2_X1 U408 ( .A1(n416), .A2(n414), .ZN(n413) );
  NOR2_X1 U409 ( .A1(G953), .A2(G237), .ZN(n477) );
  XNOR2_X1 U410 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n589) );
  XNOR2_X1 U411 ( .A(n451), .B(n430), .ZN(n405) );
  INV_X1 U412 ( .A(KEYINPUT8), .ZN(n430) );
  XNOR2_X1 U413 ( .A(n362), .B(n428), .ZN(n427) );
  XNOR2_X1 U414 ( .A(n386), .B(n385), .ZN(n428) );
  XNOR2_X1 U415 ( .A(G119), .B(KEYINPUT92), .ZN(n385) );
  XNOR2_X1 U416 ( .A(KEYINPUT10), .B(G140), .ZN(n450) );
  XNOR2_X1 U417 ( .A(n739), .B(n447), .ZN(n713) );
  XNOR2_X1 U418 ( .A(n424), .B(KEYINPUT39), .ZN(n651) );
  INV_X1 U419 ( .A(KEYINPUT1), .ZN(n449) );
  XNOR2_X1 U420 ( .A(n620), .B(n619), .ZN(n648) );
  INV_X1 U421 ( .A(KEYINPUT106), .ZN(n619) );
  AND2_X1 U422 ( .A1(n379), .A2(n364), .ZN(n620) );
  NOR2_X1 U423 ( .A1(G902), .A2(n724), .ZN(n458) );
  XNOR2_X1 U424 ( .A(n406), .B(G478), .ZN(n567) );
  NAND2_X1 U425 ( .A1(n408), .A2(n407), .ZN(n406) );
  INV_X1 U426 ( .A(G902), .ZN(n407) );
  XNOR2_X1 U427 ( .A(n474), .B(n475), .ZN(n626) );
  NOR2_X1 U428 ( .A1(n561), .A2(n611), .ZN(n583) );
  NAND2_X1 U429 ( .A1(G234), .A2(G237), .ZN(n435) );
  XNOR2_X1 U430 ( .A(G137), .B(G146), .ZN(n463) );
  XOR2_X1 U431 ( .A(KEYINPUT76), .B(KEYINPUT5), .Z(n464) );
  XOR2_X1 U432 ( .A(KEYINPUT96), .B(G116), .Z(n466) );
  XNOR2_X1 U433 ( .A(n495), .B(n437), .ZN(n462) );
  XNOR2_X1 U434 ( .A(KEYINPUT4), .B(G131), .ZN(n437) );
  XNOR2_X1 U435 ( .A(G128), .B(G110), .ZN(n386) );
  XNOR2_X1 U436 ( .A(G101), .B(G104), .ZN(n438) );
  XOR2_X1 U437 ( .A(KEYINPUT77), .B(G140), .Z(n439) );
  XNOR2_X1 U438 ( .A(G146), .B(G107), .ZN(n441) );
  XNOR2_X1 U439 ( .A(n601), .B(KEYINPUT70), .ZN(n617) );
  AND2_X1 U440 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U441 ( .A(KEYINPUT38), .B(n631), .Z(n644) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n379) );
  INV_X1 U443 ( .A(KEYINPUT28), .ZN(n380) );
  NAND2_X1 U444 ( .A1(n617), .A2(n626), .ZN(n381) );
  NOR2_X1 U445 ( .A1(n600), .A2(n598), .ZN(n420) );
  AND2_X1 U446 ( .A1(n377), .A2(n375), .ZN(n741) );
  NOR2_X1 U447 ( .A1(n704), .A2(n376), .ZN(n375) );
  XNOR2_X1 U448 ( .A(n378), .B(n421), .ZN(n377) );
  INV_X1 U449 ( .A(n702), .ZN(n376) );
  XNOR2_X1 U450 ( .A(G119), .B(KEYINPUT3), .ZN(n469) );
  NAND2_X1 U451 ( .A1(n400), .A2(n398), .ZN(n731) );
  NAND2_X1 U452 ( .A1(n402), .A2(n589), .ZN(n401) );
  XOR2_X1 U453 ( .A(G116), .B(G107), .Z(n498) );
  XOR2_X1 U454 ( .A(KEYINPUT9), .B(G122), .Z(n493) );
  XNOR2_X1 U455 ( .A(n509), .B(G134), .ZN(n495) );
  INV_X1 U456 ( .A(n509), .ZN(n510) );
  NOR2_X1 U457 ( .A1(n434), .A2(KEYINPUT79), .ZN(n652) );
  NAND2_X1 U458 ( .A1(n618), .A2(n420), .ZN(n623) );
  XNOR2_X1 U459 ( .A(n426), .B(n425), .ZN(n724) );
  XNOR2_X1 U460 ( .A(n431), .B(n484), .ZN(n425) );
  XNOR2_X1 U461 ( .A(n429), .B(n427), .ZN(n426) );
  NOR2_X1 U462 ( .A1(n505), .A2(G952), .ZN(n726) );
  INV_X1 U463 ( .A(KEYINPUT42), .ZN(n384) );
  AND2_X1 U464 ( .A1(n651), .A2(n694), .ZN(n646) );
  XNOR2_X1 U465 ( .A(KEYINPUT78), .B(KEYINPUT35), .ZN(n419) );
  OR2_X2 U466 ( .A1(n561), .A2(n559), .ZN(n560) );
  NOR2_X1 U467 ( .A1(n519), .A2(n567), .ZN(n694) );
  NAND2_X1 U468 ( .A1(n583), .A2(n368), .ZN(n688) );
  INV_X1 U469 ( .A(KEYINPUT53), .ZN(n391) );
  XNOR2_X1 U470 ( .A(n388), .B(KEYINPUT119), .ZN(n387) );
  XNOR2_X1 U471 ( .A(n506), .B(n450), .ZN(n484) );
  XNOR2_X1 U472 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n362) );
  XNOR2_X1 U473 ( .A(KEYINPUT118), .B(n543), .ZN(n363) );
  XOR2_X1 U474 ( .A(n618), .B(KEYINPUT105), .Z(n364) );
  AND2_X1 U475 ( .A1(n753), .A2(n411), .ZN(n365) );
  XNOR2_X1 U476 ( .A(KEYINPUT102), .B(n558), .ZN(n366) );
  AND2_X1 U477 ( .A1(n404), .A2(n399), .ZN(n367) );
  AND2_X1 U478 ( .A1(n562), .A2(n600), .ZN(n368) );
  AND2_X1 U479 ( .A1(G210), .A2(n517), .ZN(n369) );
  XOR2_X1 U480 ( .A(KEYINPUT19), .B(KEYINPUT67), .Z(n370) );
  OR2_X1 U481 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n371) );
  XOR2_X1 U482 ( .A(KEYINPUT65), .B(KEYINPUT46), .Z(n372) );
  NAND2_X1 U483 ( .A1(n403), .A2(n587), .ZN(n395) );
  OR2_X2 U484 ( .A1(n659), .A2(n373), .ZN(n719) );
  NOR2_X1 U485 ( .A1(n434), .A2(n667), .ZN(n373) );
  NAND2_X1 U486 ( .A1(n626), .A2(n627), .ZN(n628) );
  XNOR2_X1 U487 ( .A(n629), .B(KEYINPUT104), .ZN(n374) );
  NAND2_X1 U488 ( .A1(n422), .A2(n423), .ZN(n378) );
  NAND2_X1 U489 ( .A1(n387), .A2(n393), .ZN(n392) );
  AND2_X1 U490 ( .A1(n383), .A2(n382), .ZN(n650) );
  INV_X1 U491 ( .A(n755), .ZN(n382) );
  XNOR2_X1 U492 ( .A(n383), .B(G137), .ZN(G39) );
  XNOR2_X1 U493 ( .A(n649), .B(n384), .ZN(n383) );
  NAND2_X1 U494 ( .A1(n389), .A2(n363), .ZN(n388) );
  XNOR2_X1 U495 ( .A(n652), .B(n390), .ZN(n389) );
  INV_X1 U496 ( .A(KEYINPUT2), .ZN(n390) );
  XNOR2_X1 U497 ( .A(n392), .B(n391), .ZN(G75) );
  INV_X1 U498 ( .A(G953), .ZN(n393) );
  NAND2_X1 U499 ( .A1(n395), .A2(n589), .ZN(n394) );
  NAND2_X1 U500 ( .A1(n574), .A2(n404), .ZN(n402) );
  NAND2_X1 U501 ( .A1(n396), .A2(n587), .ZN(n398) );
  INV_X1 U502 ( .A(n589), .ZN(n399) );
  NAND2_X1 U503 ( .A1(n405), .A2(G217), .ZN(n491) );
  NAND2_X1 U504 ( .A1(n405), .A2(G221), .ZN(n429) );
  INV_X1 U505 ( .A(n721), .ZN(n408) );
  OR2_X2 U506 ( .A1(n563), .A2(n555), .ZN(n557) );
  INV_X1 U507 ( .A(n551), .ZN(n621) );
  XNOR2_X2 U508 ( .A(n606), .B(n370), .ZN(n551) );
  NAND2_X1 U509 ( .A1(n753), .A2(n418), .ZN(n415) );
  XNOR2_X2 U510 ( .A(n570), .B(n419), .ZN(n753) );
  NOR2_X1 U511 ( .A1(n571), .A2(KEYINPUT44), .ZN(n411) );
  INV_X1 U512 ( .A(n417), .ZN(n412) );
  NAND2_X1 U513 ( .A1(n415), .A2(n571), .ZN(n414) );
  NAND2_X1 U514 ( .A1(n417), .A2(n571), .ZN(n416) );
  NAND2_X1 U515 ( .A1(n754), .A2(n688), .ZN(n585) );
  INV_X1 U516 ( .A(KEYINPUT44), .ZN(n418) );
  NAND2_X1 U517 ( .A1(n611), .A2(n420), .ZN(n532) );
  OR2_X1 U518 ( .A1(n611), .A2(n420), .ZN(n526) );
  INV_X1 U519 ( .A(KEYINPUT48), .ZN(n421) );
  NOR2_X1 U520 ( .A1(n642), .A2(n641), .ZN(n422) );
  XNOR2_X1 U521 ( .A(n650), .B(n372), .ZN(n423) );
  NAND2_X1 U522 ( .A1(n643), .A2(n644), .ZN(n424) );
  XOR2_X1 U523 ( .A(n452), .B(KEYINPUT93), .Z(n431) );
  AND2_X1 U524 ( .A1(n638), .A2(n637), .ZN(n432) );
  XOR2_X1 U525 ( .A(n715), .B(n714), .Z(n433) );
  AND2_X2 U526 ( .A1(n731), .A2(n741), .ZN(n434) );
  INV_X1 U527 ( .A(G110), .ZN(n440) );
  XNOR2_X1 U528 ( .A(n441), .B(n440), .ZN(n442) );
  INV_X1 U529 ( .A(KEYINPUT71), .ZN(n571) );
  XNOR2_X1 U530 ( .A(n443), .B(n442), .ZN(n446) );
  INV_X1 U531 ( .A(KEYINPUT18), .ZN(n511) );
  XNOR2_X1 U532 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U533 ( .A(n514), .B(n513), .ZN(n515) );
  INV_X1 U534 ( .A(KEYINPUT110), .ZN(n674) );
  INV_X1 U535 ( .A(KEYINPUT25), .ZN(n455) );
  XNOR2_X1 U536 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U537 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U538 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X1 U539 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U540 ( .A(n679), .B(KEYINPUT63), .ZN(n680) );
  XNOR2_X1 U541 ( .A(n681), .B(n680), .ZN(G57) );
  XOR2_X1 U542 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n436) );
  XNOR2_X1 U543 ( .A(n436), .B(n435), .ZN(n545) );
  NAND2_X1 U544 ( .A1(G952), .A2(n545), .ZN(n547) );
  XNOR2_X1 U545 ( .A(n439), .B(n438), .ZN(n443) );
  XNOR2_X2 U546 ( .A(n444), .B(G953), .ZN(n505) );
  NAND2_X1 U547 ( .A1(G227), .A2(n505), .ZN(n445) );
  XOR2_X1 U548 ( .A(n446), .B(n445), .Z(n447) );
  NAND2_X1 U549 ( .A1(n505), .A2(G234), .ZN(n451) );
  XOR2_X1 U550 ( .A(G902), .B(KEYINPUT15), .Z(n654) );
  INV_X1 U551 ( .A(n654), .ZN(n656) );
  NAND2_X1 U552 ( .A1(G234), .A2(n656), .ZN(n454) );
  XNOR2_X1 U553 ( .A(KEYINPUT94), .B(KEYINPUT20), .ZN(n453) );
  XNOR2_X1 U554 ( .A(n454), .B(n453), .ZN(n459) );
  NAND2_X1 U555 ( .A1(n459), .A2(G217), .ZN(n456) );
  NAND2_X1 U556 ( .A1(G221), .A2(n459), .ZN(n461) );
  XOR2_X1 U557 ( .A(KEYINPUT21), .B(KEYINPUT95), .Z(n460) );
  XNOR2_X1 U558 ( .A(n461), .B(n460), .ZN(n598) );
  XNOR2_X1 U559 ( .A(G472), .B(KEYINPUT73), .ZN(n475) );
  INV_X1 U560 ( .A(n462), .ZN(n473) );
  XNOR2_X1 U561 ( .A(n464), .B(n463), .ZN(n468) );
  NAND2_X1 U562 ( .A1(n477), .A2(G210), .ZN(n465) );
  XNOR2_X1 U563 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U564 ( .A(n467), .B(n468), .ZN(n471) );
  XOR2_X1 U565 ( .A(G113), .B(G101), .Z(n470) );
  XNOR2_X1 U566 ( .A(n470), .B(n469), .ZN(n499) );
  XNOR2_X1 U567 ( .A(n471), .B(n499), .ZN(n472) );
  XNOR2_X1 U568 ( .A(n473), .B(n472), .ZN(n673) );
  NOR2_X1 U569 ( .A1(n673), .A2(G902), .ZN(n474) );
  XNOR2_X1 U570 ( .A(n626), .B(KEYINPUT6), .ZN(n591) );
  NOR2_X1 U571 ( .A1(n532), .A2(n591), .ZN(n476) );
  XNOR2_X1 U572 ( .A(n476), .B(KEYINPUT33), .ZN(n564) );
  XNOR2_X1 U573 ( .A(KEYINPUT13), .B(G475), .ZN(n490) );
  XOR2_X1 U574 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n479) );
  NAND2_X1 U575 ( .A1(G214), .A2(n477), .ZN(n478) );
  XNOR2_X1 U576 ( .A(n479), .B(n478), .ZN(n483) );
  XOR2_X1 U577 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n481) );
  XNOR2_X1 U578 ( .A(G113), .B(KEYINPUT97), .ZN(n480) );
  XNOR2_X1 U579 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U580 ( .A(n483), .B(n482), .Z(n488) );
  XNOR2_X1 U581 ( .A(G143), .B(G131), .ZN(n485) );
  XOR2_X2 U582 ( .A(G104), .B(G122), .Z(n500) );
  XNOR2_X1 U583 ( .A(n485), .B(n500), .ZN(n486) );
  XNOR2_X1 U584 ( .A(n484), .B(n486), .ZN(n487) );
  XNOR2_X1 U585 ( .A(n488), .B(n487), .ZN(n653) );
  NOR2_X1 U586 ( .A1(G902), .A2(n653), .ZN(n489) );
  XNOR2_X1 U587 ( .A(n490), .B(n489), .ZN(n568) );
  XOR2_X1 U588 ( .A(KEYINPUT100), .B(KEYINPUT7), .Z(n492) );
  XNOR2_X1 U589 ( .A(n492), .B(n491), .ZN(n497) );
  XNOR2_X1 U590 ( .A(n493), .B(n498), .ZN(n494) );
  XNOR2_X1 U591 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U592 ( .A(n497), .B(n496), .Z(n721) );
  XNOR2_X1 U593 ( .A(n499), .B(n498), .ZN(n504) );
  XOR2_X1 U594 ( .A(n500), .B(KEYINPUT16), .Z(n502) );
  XNOR2_X1 U595 ( .A(G110), .B(KEYINPUT75), .ZN(n501) );
  XNOR2_X1 U596 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U597 ( .A(n504), .B(n503), .ZN(n735) );
  AND2_X1 U598 ( .A1(G224), .A2(n505), .ZN(n508) );
  XNOR2_X1 U599 ( .A(n506), .B(KEYINPUT17), .ZN(n507) );
  XNOR2_X1 U600 ( .A(n508), .B(n507), .ZN(n514) );
  XNOR2_X1 U601 ( .A(n510), .B(KEYINPUT4), .ZN(n512) );
  XNOR2_X1 U602 ( .A(n735), .B(n515), .ZN(n708) );
  NAND2_X1 U603 ( .A1(n708), .A2(n656), .ZN(n516) );
  OR2_X1 U604 ( .A1(G237), .A2(G902), .ZN(n517) );
  BUF_X1 U605 ( .A(n550), .Z(n631) );
  NAND2_X1 U606 ( .A1(G214), .A2(n517), .ZN(n627) );
  NOR2_X1 U607 ( .A1(n644), .A2(n627), .ZN(n518) );
  NOR2_X1 U608 ( .A1(n554), .A2(n518), .ZN(n521) );
  INV_X1 U609 ( .A(n568), .ZN(n519) );
  NAND2_X1 U610 ( .A1(n519), .A2(n567), .ZN(n700) );
  INV_X1 U611 ( .A(n700), .ZN(n689) );
  NOR2_X1 U612 ( .A1(n694), .A2(n689), .ZN(n634) );
  NAND2_X1 U613 ( .A1(n644), .A2(n627), .ZN(n524) );
  NOR2_X1 U614 ( .A1(n634), .A2(n524), .ZN(n520) );
  NOR2_X1 U615 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U616 ( .A(n522), .B(KEYINPUT116), .ZN(n523) );
  NOR2_X1 U617 ( .A1(n564), .A2(n523), .ZN(n537) );
  NOR2_X1 U618 ( .A1(n524), .A2(n554), .ZN(n525) );
  XNOR2_X1 U619 ( .A(KEYINPUT41), .B(n525), .ZN(n647) );
  XNOR2_X1 U620 ( .A(n526), .B(KEYINPUT50), .ZN(n531) );
  NAND2_X1 U621 ( .A1(n600), .A2(n598), .ZN(n527) );
  XOR2_X1 U622 ( .A(KEYINPUT49), .B(n527), .Z(n528) );
  INV_X1 U623 ( .A(n626), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n528), .A2(n562), .ZN(n529) );
  XNOR2_X1 U625 ( .A(KEYINPUT115), .B(n529), .ZN(n530) );
  NAND2_X1 U626 ( .A1(n531), .A2(n530), .ZN(n533) );
  OR2_X1 U627 ( .A1(n562), .A2(n532), .ZN(n578) );
  NAND2_X1 U628 ( .A1(n533), .A2(n578), .ZN(n534) );
  XNOR2_X1 U629 ( .A(KEYINPUT51), .B(n534), .ZN(n535) );
  NOR2_X1 U630 ( .A1(n647), .A2(n535), .ZN(n536) );
  NOR2_X1 U631 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U632 ( .A(n538), .B(KEYINPUT52), .Z(n539) );
  XNOR2_X1 U633 ( .A(KEYINPUT117), .B(n539), .ZN(n540) );
  NOR2_X1 U634 ( .A1(n547), .A2(n540), .ZN(n542) );
  NOR2_X1 U635 ( .A1(n564), .A2(n647), .ZN(n541) );
  NOR2_X1 U636 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U637 ( .A(KEYINPUT89), .B(G898), .ZN(n729) );
  NAND2_X1 U638 ( .A1(n729), .A2(G953), .ZN(n544) );
  XNOR2_X1 U639 ( .A(n544), .B(KEYINPUT90), .ZN(n736) );
  NAND2_X1 U640 ( .A1(G902), .A2(n545), .ZN(n592) );
  NOR2_X1 U641 ( .A1(n736), .A2(n592), .ZN(n546) );
  XNOR2_X1 U642 ( .A(KEYINPUT91), .B(n546), .ZN(n549) );
  NOR2_X1 U643 ( .A1(G953), .A2(n547), .ZN(n548) );
  XOR2_X1 U644 ( .A(KEYINPUT88), .B(n548), .Z(n596) );
  NAND2_X1 U645 ( .A1(n549), .A2(n596), .ZN(n552) );
  NAND2_X1 U646 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U647 ( .A(n553), .B(KEYINPUT0), .ZN(n563) );
  INV_X1 U648 ( .A(n611), .ZN(n590) );
  INV_X1 U649 ( .A(n600), .ZN(n581) );
  NOR2_X1 U650 ( .A1(n590), .A2(n581), .ZN(n558) );
  NAND2_X1 U651 ( .A1(n591), .A2(n366), .ZN(n559) );
  XNOR2_X2 U652 ( .A(n560), .B(KEYINPUT32), .ZN(n754) );
  XOR2_X1 U653 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n566) );
  INV_X1 U654 ( .A(n563), .ZN(n576) );
  NOR2_X1 U655 ( .A1(n563), .A2(n564), .ZN(n565) );
  XNOR2_X1 U656 ( .A(n566), .B(n565), .ZN(n569) );
  NAND2_X1 U657 ( .A1(n568), .A2(n567), .ZN(n633) );
  NOR2_X2 U658 ( .A1(n569), .A2(n633), .ZN(n570) );
  NAND2_X1 U659 ( .A1(n585), .A2(KEYINPUT66), .ZN(n572) );
  NAND2_X1 U660 ( .A1(n572), .A2(n753), .ZN(n573) );
  NAND2_X1 U661 ( .A1(n573), .A2(KEYINPUT44), .ZN(n574) );
  INV_X1 U662 ( .A(n575), .ZN(n618) );
  NOR2_X1 U663 ( .A1(n626), .A2(n623), .ZN(n577) );
  NAND2_X1 U664 ( .A1(n577), .A2(n576), .ZN(n683) );
  NOR2_X1 U665 ( .A1(n578), .A2(n563), .ZN(n579) );
  XNOR2_X1 U666 ( .A(n579), .B(KEYINPUT31), .ZN(n699) );
  NAND2_X1 U667 ( .A1(n683), .A2(n699), .ZN(n580) );
  INV_X1 U668 ( .A(n634), .ZN(n615) );
  NAND2_X1 U669 ( .A1(n580), .A2(n615), .ZN(n588) );
  AND2_X1 U670 ( .A1(n581), .A2(n591), .ZN(n582) );
  NAND2_X1 U671 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U672 ( .A(KEYINPUT101), .B(n584), .ZN(n752) );
  NOR2_X1 U673 ( .A1(KEYINPUT66), .A2(n585), .ZN(n586) );
  NOR2_X1 U674 ( .A1(n752), .A2(n586), .ZN(n587) );
  NAND2_X1 U675 ( .A1(n590), .A2(n627), .ZN(n603) );
  INV_X1 U676 ( .A(n694), .ZN(n697) );
  NOR2_X1 U677 ( .A1(n697), .A2(n591), .ZN(n602) );
  NOR2_X1 U678 ( .A1(G900), .A2(n592), .ZN(n594) );
  INV_X1 U679 ( .A(n505), .ZN(n593) );
  NAND2_X1 U680 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U681 ( .A1(n596), .A2(n595), .ZN(n624) );
  INV_X1 U682 ( .A(n624), .ZN(n597) );
  NOR2_X1 U683 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U684 ( .A1(n602), .A2(n617), .ZN(n607) );
  NOR2_X1 U685 ( .A1(n603), .A2(n607), .ZN(n604) );
  XNOR2_X1 U686 ( .A(n604), .B(KEYINPUT43), .ZN(n605) );
  NOR2_X1 U687 ( .A1(n631), .A2(n605), .ZN(n704) );
  NOR2_X1 U688 ( .A1(n607), .A2(n606), .ZN(n609) );
  XNOR2_X1 U689 ( .A(KEYINPUT108), .B(KEYINPUT36), .ZN(n608) );
  XNOR2_X1 U690 ( .A(n609), .B(n608), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n612), .B(KEYINPUT109), .ZN(n749) );
  NOR2_X1 U693 ( .A1(KEYINPUT47), .A2(KEYINPUT80), .ZN(n613) );
  NOR2_X1 U694 ( .A1(n749), .A2(n613), .ZN(n639) );
  XOR2_X1 U695 ( .A(KEYINPUT47), .B(KEYINPUT68), .Z(n614) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n616), .A2(KEYINPUT80), .ZN(n622) );
  NOR2_X1 U698 ( .A1(n648), .A2(n621), .ZN(n695) );
  NAND2_X1 U699 ( .A1(n622), .A2(n695), .ZN(n638) );
  XNOR2_X1 U700 ( .A(n623), .B(KEYINPUT103), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n628), .B(KEYINPUT30), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n631), .A2(n643), .ZN(n632) );
  NOR2_X1 U704 ( .A1(n633), .A2(n632), .ZN(n693) );
  NAND2_X1 U705 ( .A1(KEYINPUT47), .A2(n634), .ZN(n635) );
  XNOR2_X1 U706 ( .A(KEYINPUT81), .B(n635), .ZN(n636) );
  NOR2_X1 U707 ( .A1(n693), .A2(n636), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n639), .A2(n432), .ZN(n642) );
  NAND2_X1 U709 ( .A1(KEYINPUT47), .A2(KEYINPUT80), .ZN(n640) );
  NOR2_X1 U710 ( .A1(n695), .A2(n640), .ZN(n641) );
  XOR2_X1 U711 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n645) );
  XNOR2_X1 U712 ( .A(n646), .B(n645), .ZN(n755) );
  NAND2_X1 U713 ( .A1(n651), .A2(n689), .ZN(n702) );
  XOR2_X1 U714 ( .A(n653), .B(KEYINPUT59), .Z(n661) );
  XNOR2_X1 U715 ( .A(n654), .B(KEYINPUT82), .ZN(n655) );
  AND2_X1 U716 ( .A1(n390), .A2(n655), .ZN(n669) );
  AND2_X1 U717 ( .A1(n434), .A2(n669), .ZN(n659) );
  XNOR2_X1 U718 ( .A(KEYINPUT83), .B(n656), .ZN(n657) );
  NAND2_X1 U719 ( .A1(n657), .A2(KEYINPUT2), .ZN(n658) );
  AND2_X1 U720 ( .A1(n658), .A2(KEYINPUT82), .ZN(n667) );
  NAND2_X1 U721 ( .A1(G475), .A2(n719), .ZN(n660) );
  XNOR2_X1 U722 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X1 U723 ( .A1(n662), .A2(n726), .ZN(n665) );
  INV_X1 U724 ( .A(KEYINPUT123), .ZN(n663) );
  XNOR2_X1 U725 ( .A(n663), .B(KEYINPUT60), .ZN(n664) );
  XNOR2_X1 U726 ( .A(n665), .B(n664), .ZN(G60) );
  INV_X1 U727 ( .A(G472), .ZN(n666) );
  OR2_X1 U728 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U729 ( .A1(n434), .A2(n668), .ZN(n672) );
  AND2_X1 U730 ( .A1(G472), .A2(n669), .ZN(n670) );
  AND2_X1 U731 ( .A1(n434), .A2(n670), .ZN(n671) );
  NOR2_X1 U732 ( .A1(n672), .A2(n671), .ZN(n677) );
  XOR2_X1 U733 ( .A(n673), .B(KEYINPUT62), .Z(n675) );
  NOR2_X1 U734 ( .A1(n726), .A2(n678), .ZN(n681) );
  INV_X1 U735 ( .A(KEYINPUT86), .ZN(n679) );
  NOR2_X1 U736 ( .A1(n697), .A2(n683), .ZN(n682) );
  XOR2_X1 U737 ( .A(G104), .B(n682), .Z(G6) );
  NOR2_X1 U738 ( .A1(n683), .A2(n700), .ZN(n687) );
  XOR2_X1 U739 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n685) );
  XNOR2_X1 U740 ( .A(G107), .B(KEYINPUT111), .ZN(n684) );
  XNOR2_X1 U741 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U742 ( .A(n687), .B(n686), .ZN(G9) );
  XNOR2_X1 U743 ( .A(G110), .B(n688), .ZN(G12) );
  XOR2_X1 U744 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n691) );
  NAND2_X1 U745 ( .A1(n695), .A2(n689), .ZN(n690) );
  XNOR2_X1 U746 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U747 ( .A(G128), .B(n692), .ZN(G30) );
  XOR2_X1 U748 ( .A(G143), .B(n693), .Z(G45) );
  NAND2_X1 U749 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U750 ( .A(n696), .B(G146), .ZN(G48) );
  NOR2_X1 U751 ( .A1(n697), .A2(n699), .ZN(n698) );
  XOR2_X1 U752 ( .A(G113), .B(n698), .Z(G15) );
  NOR2_X1 U753 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U754 ( .A(G116), .B(n701), .Z(G18) );
  XNOR2_X1 U755 ( .A(G134), .B(KEYINPUT114), .ZN(n703) );
  XNOR2_X1 U756 ( .A(n703), .B(n702), .ZN(G36) );
  XOR2_X1 U757 ( .A(G140), .B(n704), .Z(G42) );
  XOR2_X1 U758 ( .A(KEYINPUT85), .B(KEYINPUT55), .Z(n706) );
  XNOR2_X1 U759 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n708), .B(n707), .ZN(n710) );
  NAND2_X1 U762 ( .A1(n719), .A2(G210), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n711), .A2(n726), .ZN(n712) );
  XNOR2_X1 U765 ( .A(n712), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U766 ( .A1(n719), .A2(G469), .ZN(n716) );
  XOR2_X1 U767 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n715) );
  XNOR2_X1 U768 ( .A(n713), .B(KEYINPUT121), .ZN(n714) );
  XNOR2_X1 U769 ( .A(n716), .B(n433), .ZN(n717) );
  XNOR2_X1 U770 ( .A(KEYINPUT122), .B(n718), .ZN(G54) );
  NAND2_X1 U771 ( .A1(G478), .A2(n719), .ZN(n720) );
  XNOR2_X1 U772 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U773 ( .A1(n726), .A2(n722), .ZN(G63) );
  NAND2_X1 U774 ( .A1(G217), .A2(n719), .ZN(n723) );
  XNOR2_X1 U775 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U776 ( .A1(n726), .A2(n725), .ZN(G66) );
  NAND2_X1 U777 ( .A1(G953), .A2(G224), .ZN(n727) );
  XOR2_X1 U778 ( .A(KEYINPUT61), .B(n727), .Z(n728) );
  NOR2_X1 U779 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U780 ( .A(KEYINPUT124), .B(n730), .Z(n733) );
  NAND2_X1 U781 ( .A1(n393), .A2(n731), .ZN(n732) );
  NAND2_X1 U782 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U783 ( .A(n734), .B(KEYINPUT125), .ZN(n738) );
  NAND2_X1 U784 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U785 ( .A(n738), .B(n737), .ZN(G69) );
  XNOR2_X1 U786 ( .A(n739), .B(n484), .ZN(n740) );
  XOR2_X1 U787 ( .A(n740), .B(KEYINPUT126), .Z(n743) );
  XOR2_X1 U788 ( .A(n743), .B(n741), .Z(n742) );
  NAND2_X1 U789 ( .A1(n742), .A2(n505), .ZN(n748) );
  XNOR2_X1 U790 ( .A(G227), .B(n743), .ZN(n744) );
  NAND2_X1 U791 ( .A1(n744), .A2(G900), .ZN(n745) );
  XOR2_X1 U792 ( .A(KEYINPUT127), .B(n745), .Z(n746) );
  NAND2_X1 U793 ( .A1(G953), .A2(n746), .ZN(n747) );
  NAND2_X1 U794 ( .A1(n748), .A2(n747), .ZN(G72) );
  XOR2_X1 U795 ( .A(KEYINPUT37), .B(KEYINPUT113), .Z(n751) );
  XNOR2_X1 U796 ( .A(G125), .B(n749), .ZN(n750) );
  XNOR2_X1 U797 ( .A(n751), .B(n750), .ZN(G27) );
  XOR2_X1 U798 ( .A(G101), .B(n752), .Z(G3) );
  XNOR2_X1 U799 ( .A(n753), .B(G122), .ZN(G24) );
  XNOR2_X1 U800 ( .A(G119), .B(n754), .ZN(G21) );
  XOR2_X1 U801 ( .A(n755), .B(G131), .Z(G33) );
endmodule

