//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(KEYINPUT65), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n207), .B1(new_n208), .B2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G13), .ZN(new_n210));
  NAND4_X1  g0010(.A1(new_n210), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT66), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n201), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT67), .Z(new_n222));
  AOI21_X1  g0022(.A(new_n214), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n208), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT68), .Z(new_n231));
  INV_X1    g0031(.A(KEYINPUT1), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n231), .A2(new_n232), .ZN(new_n234));
  AND3_X1   g0034(.A1(new_n223), .A2(new_n233), .A3(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT69), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT2), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n239), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G223), .ZN(new_n255));
  INV_X1    g0055(.A(G77), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n254), .A2(new_n255), .B1(new_n256), .B2(new_n253), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G222), .ZN(new_n260));
  OR3_X1    g0060(.A1(new_n259), .A2(KEYINPUT71), .A3(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(KEYINPUT71), .B1(new_n259), .B2(new_n260), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n216), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT70), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(KEYINPUT70), .A2(G33), .A3(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(new_n216), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(G226), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n272), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n270), .A2(G274), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n266), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT76), .B(G200), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(KEYINPUT72), .A3(new_n215), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT72), .B1(new_n281), .B2(new_n215), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n271), .A2(G13), .A3(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT74), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT74), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n288), .A2(new_n271), .A3(G13), .A4(G20), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G20), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G1), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(G50), .A3(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G33), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT73), .B1(new_n298), .B2(G20), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT73), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(new_n292), .A3(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT8), .B(G58), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n297), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n285), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n287), .A2(new_n289), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n295), .B(new_n306), .C1(G50), .C2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT9), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n277), .A2(G190), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n280), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n280), .A2(new_n309), .A3(new_n313), .A4(new_n310), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n270), .A2(G238), .A3(new_n272), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(G226), .A2(G1698), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n241), .B2(G1698), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n318), .B1(new_n320), .B2(new_n253), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n316), .B(new_n275), .C1(new_n321), .C2(new_n265), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT13), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n241), .A2(G1698), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(G226), .B2(G1698), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n317), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n265), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n332), .A2(new_n333), .A3(new_n316), .A4(new_n275), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n323), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G169), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT14), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n323), .A2(G179), .A3(new_n334), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n335), .A2(new_n339), .A3(G169), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n296), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n342), .A2(new_n202), .B1(new_n292), .B2(G68), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(G77), .B2(new_n302), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n281), .A2(new_n215), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT72), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n282), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT11), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT11), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n303), .A2(new_n256), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n350), .B(new_n285), .C1(new_n351), .C2(new_n343), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G68), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n287), .A2(new_n354), .A3(new_n289), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT77), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT12), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT12), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n293), .A2(new_n354), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n359), .A2(new_n360), .B1(new_n291), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n353), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n341), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT16), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT80), .B1(new_n327), .B2(G33), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT80), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(new_n298), .A3(KEYINPUT3), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n370), .A3(new_n328), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(G20), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n253), .B2(G20), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n354), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G58), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(new_n354), .ZN(new_n378));
  OAI21_X1  g0178(.A(G20), .B1(new_n378), .B2(new_n201), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n296), .A2(G159), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n367), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT7), .B1(new_n329), .B2(new_n292), .ZN(new_n383));
  AOI211_X1 g0183(.A(new_n372), .B(G20), .C1(new_n326), .C2(new_n328), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n381), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(KEYINPUT16), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n382), .A2(new_n285), .A3(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n304), .A2(new_n293), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n348), .A2(new_n307), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n290), .A2(new_n304), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT81), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT81), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n270), .A2(G232), .A3(new_n272), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT82), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n275), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n399), .B1(new_n275), .B2(new_n398), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n255), .A2(new_n258), .ZN(new_n404));
  INV_X1    g0204(.A(G226), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G1698), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G87), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n329), .A2(new_n407), .B1(new_n298), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n409), .A2(new_n331), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(G179), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n331), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(new_n275), .A3(new_n398), .ZN(new_n413));
  INV_X1    g0213(.A(G169), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n403), .A2(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n397), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT18), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n397), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n275), .A2(new_n398), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT82), .ZN(new_n421));
  AOI21_X1  g0221(.A(G190), .B1(new_n409), .B2(new_n331), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n400), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G200), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n410), .B2(new_n420), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(new_n388), .A3(new_n396), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n327), .A2(G33), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n431));
  OAI211_X1 g0231(.A(KEYINPUT7), .B(new_n292), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n375), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n381), .B1(new_n433), .B2(G68), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n348), .B1(new_n434), .B2(KEYINPUT16), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n435), .A2(new_n382), .B1(new_n393), .B2(new_n395), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(KEYINPUT17), .A3(new_n426), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n417), .A2(new_n419), .A3(new_n429), .A4(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n366), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G179), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n277), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n308), .C1(G169), .C2(new_n277), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n291), .A2(G77), .A3(new_n294), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT75), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n304), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n446), .A2(new_n296), .B1(G20), .B2(G77), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT15), .B(G87), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n303), .B2(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n449), .A2(new_n285), .B1(new_n256), .B2(new_n290), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n329), .A2(G107), .ZN(new_n452));
  INV_X1    g0252(.A(G238), .ZN(new_n453));
  OAI221_X1 g0253(.A(new_n452), .B1(new_n259), .B2(new_n241), .C1(new_n453), .C2(new_n254), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n331), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n270), .A2(G244), .A3(new_n272), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n275), .A3(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n457), .A2(G179), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n414), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n451), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n279), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n455), .A2(G190), .A3(new_n275), .A4(new_n456), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n461), .A2(new_n445), .A3(new_n450), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n315), .A2(new_n439), .A3(new_n442), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT78), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n323), .A2(G190), .A3(new_n334), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(new_n353), .A3(new_n362), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n424), .B1(new_n323), .B2(new_n334), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n470), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n363), .A2(new_n472), .A3(KEYINPUT78), .A4(new_n468), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT79), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n474), .B1(new_n471), .B2(new_n473), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n466), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT87), .A2(KEYINPUT21), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n271), .A2(G33), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n348), .A2(G116), .A3(new_n307), .A4(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G116), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n290), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  AND2_X1   g0285(.A1(KEYINPUT83), .A2(G97), .ZN(new_n486));
  NOR2_X1   g0286(.A1(KEYINPUT83), .A2(G97), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n292), .B(new_n485), .C1(new_n488), .C2(G33), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n281), .A2(new_n215), .B1(G20), .B2(new_n483), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT20), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g0291(.A1(KEYINPUT83), .A2(G97), .ZN(new_n492));
  NAND2_X1  g0292(.A1(KEYINPUT83), .A2(G97), .ZN(new_n493));
  AOI21_X1  g0293(.A(G33), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n485), .A2(new_n292), .ZN(new_n495));
  OAI211_X1 g0295(.A(KEYINPUT20), .B(new_n490), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n482), .B(new_n484), .C1(new_n491), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G169), .ZN(new_n499));
  INV_X1    g0299(.A(G41), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n271), .B(G45), .C1(new_n500), .C2(KEYINPUT5), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT85), .B1(new_n500), .B2(KEYINPUT5), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(KEYINPUT85), .A3(KEYINPUT5), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n503), .A2(G274), .A3(new_n270), .A4(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT85), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(G41), .ZN(new_n508));
  INV_X1    g0308(.A(G45), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G1), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(G41), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n508), .A2(new_n504), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(G270), .A3(new_n270), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n505), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n326), .A2(new_n328), .A3(G264), .A4(G1698), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n326), .A2(new_n328), .A3(G257), .A4(new_n258), .ZN(new_n516));
  INV_X1    g0316(.A(G303), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n515), .B(new_n516), .C1(new_n517), .C2(new_n253), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n331), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT86), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(KEYINPUT86), .A3(new_n331), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n514), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n480), .B1(new_n499), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(G179), .A3(new_n498), .ZN(new_n525));
  INV_X1    g0325(.A(new_n514), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n518), .A2(KEYINPUT86), .A3(new_n331), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT86), .B1(new_n518), .B2(new_n331), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n480), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n529), .A2(G169), .A3(new_n498), .A4(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n524), .A2(new_n525), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n498), .B1(new_n529), .B2(G200), .ZN(new_n533));
  OR2_X1    g0333(.A1(new_n533), .A2(KEYINPUT88), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(KEYINPUT88), .B1(G190), .B2(new_n523), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n348), .A2(new_n307), .A3(new_n481), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT84), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n448), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n348), .A2(KEYINPUT84), .A3(new_n307), .A4(new_n481), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(G107), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n492), .A2(new_n408), .A3(new_n543), .A4(new_n493), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n292), .B1(new_n317), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n253), .A2(new_n292), .A3(G68), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n299), .A2(new_n301), .B1(new_n492), .B2(new_n493), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n547), .B(new_n548), .C1(KEYINPUT19), .C2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(new_n285), .B1(new_n290), .B2(new_n448), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n542), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(G250), .B1(new_n271), .B2(G45), .ZN(new_n553));
  INV_X1    g0353(.A(G274), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(new_n510), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n555), .A2(new_n270), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n453), .A2(new_n258), .ZN(new_n557));
  INV_X1    g0357(.A(G244), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G1698), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n253), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G116), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n265), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n414), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n561), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(new_n331), .B1(new_n270), .B2(new_n555), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n440), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n552), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n539), .A2(G87), .A3(new_n541), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(G190), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n279), .B1(new_n556), .B2(new_n562), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n568), .A2(new_n551), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n539), .A2(G97), .A3(new_n541), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT6), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(G107), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n486), .B2(new_n487), .ZN(new_n577));
  AND2_X1   g0377(.A1(G97), .A2(G107), .ZN(new_n578));
  NOR2_X1   g0378(.A1(G97), .A2(G107), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G20), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n296), .A2(G77), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n543), .B1(new_n374), .B2(new_n375), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n285), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n307), .A2(G97), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n574), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n512), .A2(G257), .A3(new_n270), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n505), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n326), .A2(new_n328), .A3(G250), .A4(G1698), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n326), .A2(new_n328), .A3(G244), .A4(new_n258), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT4), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n485), .B(new_n592), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n331), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n591), .A2(new_n597), .A3(new_n440), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n591), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n414), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n589), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n539), .A2(G107), .A3(new_n541), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n307), .A2(G107), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT25), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n326), .A2(new_n328), .A3(new_n292), .A4(G87), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT22), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT22), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n253), .A2(new_n608), .A3(new_n292), .A4(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT24), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n298), .A2(new_n483), .A3(G20), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT23), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n292), .B2(G107), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n543), .A2(KEYINPUT23), .A3(G20), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n610), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n611), .B1(new_n610), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n285), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n512), .A2(new_n270), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n326), .A2(new_n328), .A3(G257), .A4(G1698), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n326), .A2(new_n328), .A3(G250), .A4(new_n258), .ZN(new_n622));
  NAND2_X1  g0422(.A1(G33), .A2(G294), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n620), .A2(G264), .B1(new_n624), .B2(new_n331), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(G190), .A3(new_n505), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n331), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n512), .A2(G264), .A3(new_n270), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n505), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G200), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n605), .A2(new_n619), .A3(new_n626), .A4(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n619), .A2(new_n602), .A3(new_n604), .ZN(new_n632));
  AOI21_X1  g0432(.A(G169), .B1(new_n625), .B2(new_n505), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n629), .A2(G179), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n329), .A2(new_n292), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n372), .B1(new_n371), .B2(new_n373), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n583), .B(new_n582), .C1(new_n638), .C2(new_n543), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n587), .B1(new_n639), .B2(new_n285), .ZN(new_n640));
  INV_X1    g0440(.A(G190), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n591), .A2(new_n597), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(G200), .B1(new_n591), .B2(new_n597), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n640), .B(new_n574), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n601), .A2(new_n631), .A3(new_n636), .A4(new_n644), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n479), .A2(new_n536), .A3(new_n573), .A4(new_n645), .ZN(G372));
  AOI21_X1  g0446(.A(KEYINPUT17), .B1(new_n436), .B2(new_n426), .ZN(new_n647));
  AND4_X1   g0447(.A1(KEYINPUT17), .A2(new_n426), .A3(new_n388), .A4(new_n396), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n460), .B1(new_n471), .B2(new_n473), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n649), .B1(new_n650), .B2(new_n366), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n421), .A2(new_n440), .A3(new_n412), .A4(new_n400), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n413), .A2(new_n414), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n436), .A2(KEYINPUT18), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n418), .B1(new_n397), .B2(new_n415), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n315), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n442), .ZN(new_n660));
  INV_X1    g0460(.A(new_n479), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n636), .A2(new_n525), .A3(new_n524), .A4(new_n531), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n566), .A2(new_n563), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n551), .B2(new_n542), .ZN(new_n664));
  INV_X1    g0464(.A(new_n569), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n568), .A2(new_n570), .A3(new_n551), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT89), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n568), .A2(new_n551), .A3(KEYINPUT89), .A4(new_n570), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n644), .A2(new_n601), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n662), .A2(new_n670), .A3(new_n671), .A4(new_n631), .ZN(new_n672));
  INV_X1    g0472(.A(new_n601), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT26), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n572), .A2(new_n675), .A3(new_n601), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n672), .B(new_n567), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n660), .B1(new_n661), .B2(new_n678), .ZN(G369));
  NAND3_X1  g0479(.A1(new_n271), .A2(new_n292), .A3(G13), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT90), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT27), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G343), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n498), .ZN(new_n688));
  MUX2_X1   g0488(.A(new_n532), .B(new_n536), .S(new_n688), .Z(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n626), .A2(new_n630), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n632), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n686), .B1(new_n605), .B2(new_n619), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n636), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n632), .A2(new_n635), .A3(new_n686), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n690), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n695), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n532), .A2(new_n686), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(new_n702), .B2(new_n694), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(G399));
  NOR2_X1   g0504(.A1(new_n544), .A2(G116), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G1), .ZN(new_n706));
  INV_X1    g0506(.A(new_n212), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  MUX2_X1   g0508(.A(new_n706), .B(new_n221), .S(new_n708), .Z(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT92), .Z(new_n710));
  XNOR2_X1  g0510(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n677), .A2(new_n686), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(KEYINPUT29), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n666), .A2(new_n667), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n569), .A3(new_n669), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n567), .A3(new_n673), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT26), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n573), .A2(new_n675), .A3(new_n673), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n672), .A2(new_n719), .A3(new_n567), .A4(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n715), .B1(new_n721), .B2(new_n686), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n714), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G330), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT93), .ZN(new_n726));
  OAI211_X1 g0526(.A(G179), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n625), .A2(new_n591), .A3(new_n597), .A4(new_n565), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n565), .A2(G179), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n730), .A2(new_n599), .A3(new_n629), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n729), .A2(KEYINPUT30), .B1(new_n731), .B2(new_n529), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n726), .B(new_n733), .C1(new_n727), .C2(new_n728), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n725), .B(new_n686), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n729), .A2(KEYINPUT30), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n731), .A2(new_n529), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT31), .B1(new_n738), .B2(new_n687), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n536), .A2(new_n645), .A3(new_n573), .A4(new_n686), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n724), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n723), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n712), .B1(new_n745), .B2(G1), .ZN(G364));
  INV_X1    g0546(.A(new_n690), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n210), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n271), .B1(new_n748), .B2(G45), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n708), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G330), .B2(new_n689), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n212), .A2(G355), .A3(new_n253), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G116), .B2(new_n212), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n248), .A2(new_n509), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n212), .A2(new_n329), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n222), .B2(new_n509), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n215), .B1(G20), .B2(new_n414), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n751), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n292), .A2(new_n440), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(G190), .A3(new_n424), .ZN(new_n768));
  INV_X1    g0568(.A(G322), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n329), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n292), .A2(G179), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n771), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n770), .B(new_n774), .C1(G329), .C2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n279), .A2(new_n641), .A3(new_n775), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G283), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n279), .A2(G190), .A3(new_n775), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G303), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n778), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n767), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n786), .A2(new_n641), .A3(new_n424), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n641), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n292), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G326), .A2(new_n787), .B1(new_n790), .B2(G294), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n767), .A2(new_n641), .A3(G200), .ZN(new_n792));
  XOR2_X1   g0592(.A(KEYINPUT33), .B(G317), .Z(new_n793));
  OAI21_X1  g0593(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n792), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n787), .A2(G50), .B1(new_n795), .B2(G68), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n776), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n796), .B1(KEYINPUT32), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n779), .A2(new_n543), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G87), .B2(new_n783), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n253), .B1(new_n772), .B2(new_n256), .ZN(new_n803));
  INV_X1    g0603(.A(new_n768), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(G58), .B2(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n799), .A2(KEYINPUT32), .B1(new_n790), .B2(G97), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n802), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n785), .A2(new_n794), .B1(new_n800), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n766), .B1(new_n808), .B2(new_n763), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n762), .B(KEYINPUT94), .Z(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n689), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n753), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(G396));
  OR2_X1    g0613(.A1(new_n460), .A2(new_n687), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n451), .A2(new_n687), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n463), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n460), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n713), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT98), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n464), .A2(new_n687), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n677), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n751), .B1(new_n824), .B2(new_n743), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n743), .B2(new_n824), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n763), .A2(new_n760), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n750), .B(new_n708), .C1(new_n256), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n763), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n779), .A2(new_n408), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G303), .A2(new_n787), .B1(new_n790), .B2(G97), .ZN(new_n831));
  INV_X1    g0631(.A(new_n772), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n804), .A2(G294), .B1(new_n832), .B2(G116), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n831), .B(new_n833), .C1(new_n773), .C2(new_n776), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n792), .A2(KEYINPUT95), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n792), .A2(KEYINPUT95), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n830), .B(new_n834), .C1(G283), .C2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n329), .B1(new_n782), .B2(new_n543), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT96), .Z(new_n841));
  AOI22_X1  g0641(.A1(new_n804), .A2(G143), .B1(new_n832), .B2(G159), .ZN(new_n842));
  INV_X1    g0642(.A(G150), .ZN(new_n843));
  INV_X1    g0643(.A(G137), .ZN(new_n844));
  INV_X1    g0644(.A(new_n787), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n842), .B1(new_n843), .B2(new_n792), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n780), .A2(G68), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n783), .A2(G50), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n790), .A2(G58), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n329), .B1(new_n777), .B2(G132), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n846), .B2(new_n847), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n839), .A2(new_n841), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n818), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n828), .B1(new_n829), .B2(new_n855), .C1(new_n856), .C2(new_n761), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n826), .A2(new_n857), .ZN(G384));
  OR2_X1    g0658(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n219), .A2(new_n859), .A3(G116), .A4(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT36), .Z(new_n862));
  OR3_X1    g0662(.A1(new_n221), .A2(new_n256), .A3(new_n378), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n202), .A2(G68), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n271), .B(G13), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n479), .B1(new_n714), .B2(new_n722), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n660), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT101), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT102), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n354), .B1(new_n375), .B2(new_n432), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n367), .B1(new_n873), .B2(new_n381), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n387), .A2(new_n874), .A3(new_n285), .ZN(new_n875));
  INV_X1    g0675(.A(new_n392), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT100), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(KEYINPUT100), .A3(new_n876), .ZN(new_n880));
  INV_X1    g0680(.A(new_n685), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n654), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n872), .B1(new_n883), .B2(new_n427), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n397), .A2(new_n685), .ZN(new_n885));
  AND4_X1   g0685(.A1(new_n872), .A2(new_n416), .A3(new_n885), .A4(new_n427), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n879), .A2(new_n685), .A3(new_n880), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n657), .B2(new_n649), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n438), .A2(new_n397), .A3(new_n685), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n416), .A2(new_n885), .A3(new_n427), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT37), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n416), .A2(new_n885), .A3(new_n872), .A4(new_n427), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n871), .B1(new_n891), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT99), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n341), .A2(new_n899), .A3(new_n364), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n899), .B1(new_n341), .B2(new_n364), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n686), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n890), .B1(new_n887), .B2(new_n889), .ZN(new_n905));
  INV_X1    g0705(.A(new_n888), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n438), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n907), .B(KEYINPUT38), .C1(new_n886), .C2(new_n884), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n905), .A2(new_n908), .A3(KEYINPUT39), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n898), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n823), .A2(new_n814), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n905), .A2(new_n908), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n365), .A2(KEYINPUT99), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n363), .A2(new_n686), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n471), .B2(new_n473), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(new_n900), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n471), .A2(new_n473), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT79), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n341), .B1(new_n918), .B2(new_n475), .ZN(new_n919));
  INV_X1    g0719(.A(new_n914), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n911), .A2(new_n912), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n881), .B1(new_n655), .B2(new_n656), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n910), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n870), .B(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT103), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n686), .B1(new_n732), .B2(new_n734), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n926), .B1(new_n927), .B2(KEYINPUT31), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT104), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n927), .A2(KEYINPUT104), .A3(KEYINPUT31), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n738), .A2(new_n687), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(KEYINPUT103), .A3(new_n725), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n741), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n341), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n476), .B2(new_n477), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n914), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n818), .B1(new_n940), .B2(new_n916), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n892), .A2(new_n896), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n908), .B1(new_n942), .B2(KEYINPUT38), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n937), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n921), .B(new_n856), .C1(new_n933), .C2(new_n936), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT40), .B1(new_n905), .B2(new_n908), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n944), .A2(KEYINPUT40), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n933), .A2(new_n936), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n948), .B1(new_n661), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n891), .A2(new_n897), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT40), .B1(new_n945), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n937), .A2(new_n941), .A3(new_n947), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n479), .A3(new_n937), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n950), .A2(G330), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n925), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n271), .B2(new_n748), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n925), .A2(new_n956), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n866), .B1(new_n958), .B2(new_n959), .ZN(G367));
  XNOR2_X1  g0760(.A(new_n697), .B(new_n701), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(new_n747), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n962), .A2(new_n723), .A3(new_n743), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT107), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n687), .A2(new_n589), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n671), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n673), .A2(new_n687), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n703), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT45), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n703), .ZN(new_n972));
  INV_X1    g0772(.A(new_n968), .ZN(new_n973));
  AOI21_X1  g0773(.A(KEYINPUT44), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n972), .A2(KEYINPUT44), .A3(new_n973), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n971), .B(new_n699), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n974), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n698), .B1(new_n977), .B2(new_n970), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n963), .A2(new_n964), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n978), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n745), .A2(new_n962), .ZN(new_n981));
  OAI21_X1  g0781(.A(KEYINPUT107), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n744), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n708), .B(KEYINPUT41), .Z(new_n984));
  OAI21_X1  g0784(.A(new_n749), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n696), .A2(new_n968), .A3(new_n702), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT105), .Z(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n601), .B1(new_n966), .B2(new_n636), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n686), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT43), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n568), .A2(new_n551), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n687), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n996), .A2(new_n567), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n670), .B2(new_n996), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n988), .A2(new_n993), .A3(new_n994), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n994), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n998), .A2(new_n994), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n987), .B(KEYINPUT105), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1000), .B(new_n1002), .C1(new_n1003), .C2(new_n992), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n999), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n699), .A2(new_n973), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT106), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1005), .B1(new_n699), .B2(new_n973), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT106), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n999), .A2(new_n1010), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n985), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n239), .A2(new_n757), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n764), .B1(new_n212), .B2(new_n448), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n751), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n768), .A2(new_n843), .B1(new_n772), .B2(new_n202), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n329), .B(new_n1018), .C1(G137), .C2(new_n777), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n838), .A2(G159), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G143), .A2(new_n787), .B1(new_n790), .B2(G68), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G58), .A2(new_n783), .B1(new_n780), .B2(G77), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n253), .B1(new_n777), .B2(G317), .ZN(new_n1024));
  INV_X1    g0824(.A(G283), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n772), .C1(new_n517), .C2(new_n768), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n845), .A2(new_n773), .B1(new_n543), .B2(new_n789), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(G294), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n837), .C1(new_n488), .C2(new_n779), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT46), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n782), .A2(new_n483), .B1(KEYINPUT108), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(KEYINPUT108), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1023), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT47), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1017), .B1(new_n1036), .B2(new_n763), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n810), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n998), .A2(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1014), .A2(new_n1041), .ZN(G387));
  OR3_X1    g0842(.A1(new_n244), .A2(new_n509), .A3(new_n253), .ZN(new_n1043));
  OAI21_X1  g0843(.A(KEYINPUT50), .B1(new_n304), .B2(G50), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1044), .B(new_n509), .C1(new_n354), .C2(new_n256), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n304), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n329), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n705), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n707), .B1(new_n1043), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n764), .B1(new_n543), .B2(new_n212), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n751), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n789), .A2(new_n448), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n253), .B1(new_n202), .B2(new_n768), .C1(new_n845), .C2(new_n797), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(G97), .C2(new_n780), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n792), .A2(new_n304), .B1(new_n772), .B2(new_n354), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT110), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n782), .A2(new_n256), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G150), .B2(new_n777), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT109), .Z(new_n1059));
  NAND3_X1  g0859(.A1(new_n1054), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n253), .B1(new_n777), .B2(G326), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n782), .A2(new_n1029), .B1(new_n789), .B2(new_n1025), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n804), .A2(G317), .B1(new_n832), .B2(G303), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n769), .B2(new_n845), .C1(new_n837), .C2(new_n773), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT48), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT49), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1061), .B1(new_n483), .B2(new_n779), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1060), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1051), .B1(new_n1071), .B2(new_n763), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n696), .B2(new_n810), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT111), .Z(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n750), .B2(new_n962), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n981), .A2(new_n708), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n745), .A2(new_n962), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(G393));
  NAND2_X1  g0878(.A1(new_n980), .A2(new_n981), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n708), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n979), .B2(new_n982), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n251), .A2(new_n757), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n764), .B1(new_n212), .B2(new_n488), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n751), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n787), .A2(G150), .B1(new_n804), .B2(G159), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT51), .Z(new_n1086));
  AOI211_X1 g0886(.A(new_n329), .B(new_n830), .C1(G143), .C2(new_n777), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(new_n354), .C2(new_n782), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n790), .A2(G77), .B1(new_n832), .B2(new_n446), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n837), .B2(new_n202), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT112), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n838), .A2(G303), .B1(G116), .B2(new_n790), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT113), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n787), .A2(G317), .B1(new_n804), .B2(G311), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT52), .Z(new_n1096));
  OAI221_X1 g0896(.A(new_n329), .B1(new_n776), .B2(new_n769), .C1(new_n1029), .C2(new_n772), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n801), .B(new_n1097), .C1(G283), .C2(new_n783), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1088), .A2(new_n1091), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1084), .B1(new_n1101), .B2(new_n763), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n762), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1102), .B1(new_n968), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n980), .B2(new_n749), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1081), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G390));
  OAI21_X1  g0907(.A(new_n903), .B1(new_n891), .B2(new_n897), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n721), .A2(new_n686), .A3(new_n817), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n814), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1108), .B1(new_n921), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n742), .A2(new_n856), .A3(new_n921), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n460), .A2(new_n687), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n677), .B2(new_n822), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n901), .A2(new_n902), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n939), .A2(new_n914), .B1(new_n1116), .B2(new_n915), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n903), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1118), .A2(KEYINPUT114), .B1(new_n898), .B2(new_n909), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT114), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1120), .B(new_n903), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1111), .B(new_n1113), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1122));
  NOR4_X1   g0922(.A1(new_n949), .A2(new_n1117), .A3(new_n724), .A4(new_n818), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1118), .A2(KEYINPUT114), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n898), .A2(new_n909), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n1126), .A3(new_n1121), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1111), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1124), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1122), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n949), .A2(new_n724), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n479), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1132), .A2(new_n867), .A3(new_n660), .ZN(new_n1133));
  OAI211_X1 g0933(.A(G330), .B(new_n856), .C1(new_n933), .C2(new_n936), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1134), .A2(new_n1117), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1109), .A2(new_n814), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1112), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT115), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n724), .B(new_n818), .C1(new_n740), .C2(new_n741), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1110), .B1(new_n1139), .B2(new_n921), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT115), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1134), .A2(new_n1117), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1139), .A2(new_n921), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n911), .B1(new_n1123), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1133), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1130), .A2(new_n1147), .ZN(new_n1148));
  AND4_X1   g0948(.A1(new_n1141), .A2(new_n1142), .A3(new_n1136), .A4(new_n1112), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1141), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1146), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1133), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1127), .A2(new_n1128), .A3(new_n1112), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1111), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1154), .B1(new_n1155), .B2(new_n1124), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1148), .A2(new_n1157), .A3(new_n708), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1126), .A2(new_n760), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n827), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n751), .B1(new_n446), .B2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT116), .Z(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n253), .B1(new_n776), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(G128), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n845), .A2(new_n1165), .B1(new_n797), .B2(new_n789), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(G132), .C2(new_n804), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n782), .A2(new_n843), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT53), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n838), .A2(G137), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT54), .B(G143), .Z(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT117), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1172), .A2(new_n832), .B1(new_n780), .B2(G50), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1167), .A2(new_n1169), .A3(new_n1170), .A4(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n837), .A2(new_n543), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n768), .A2(new_n483), .B1(new_n772), .B2(new_n488), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n253), .B(new_n1176), .C1(G294), .C2(new_n777), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n783), .A2(G87), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G283), .A2(new_n787), .B1(new_n790), .B2(G77), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n849), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1174), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1162), .B1(new_n1181), .B2(new_n763), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1130), .A2(new_n750), .B1(new_n1159), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1158), .A2(new_n1183), .ZN(G378));
  AOI22_X1  g0984(.A1(G116), .A2(new_n787), .B1(new_n790), .B2(G68), .ZN(new_n1185));
  INV_X1    g0985(.A(G97), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1185), .B1(new_n1186), .B2(new_n792), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n804), .A2(G107), .B1(new_n777), .B2(G283), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n253), .A2(G41), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n448), .C2(new_n772), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n779), .A2(new_n377), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1187), .A2(new_n1190), .A3(new_n1057), .A4(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT118), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(KEYINPUT58), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(G33), .A2(G41), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1189), .A2(G50), .A3(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT119), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1172), .A2(new_n783), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n768), .A2(new_n1165), .B1(new_n772), .B2(new_n844), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G132), .B2(new_n795), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G125), .A2(new_n787), .B1(new_n790), .B2(G150), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1199), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT59), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(KEYINPUT120), .ZN(new_n1205));
  INV_X1    g1005(.A(G124), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1195), .B1(new_n1206), .B2(new_n776), .C1(new_n779), .C2(new_n797), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1204), .B2(KEYINPUT120), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(KEYINPUT58), .A2(new_n1193), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n829), .B1(new_n1198), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n751), .B1(G50), .B2(new_n1160), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n315), .A2(new_n442), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n308), .A2(new_n685), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT55), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1212), .B(new_n1214), .ZN(new_n1215));
  XOR2_X1   g1015(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1216));
  XNOR2_X1  g1016(.A(new_n1215), .B(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1210), .B(new_n1211), .C1(new_n1218), .C2(new_n760), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n954), .A2(G330), .A3(new_n924), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n924), .B1(new_n954), .B2(G330), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1217), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n910), .A2(new_n922), .A3(new_n923), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n948), .B2(new_n724), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n954), .A2(G330), .A3(new_n924), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n1225), .A3(new_n1218), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1222), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1219), .B1(new_n1227), .B2(new_n750), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(KEYINPUT57), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1133), .B1(new_n1130), .B2(new_n1147), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n708), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1152), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT57), .B1(new_n1232), .B2(new_n1227), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1228), .B1(new_n1231), .B2(new_n1233), .ZN(G375));
  INV_X1    g1034(.A(new_n984), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1146), .B(new_n1133), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1153), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n377), .A2(new_n779), .B1(new_n782), .B2(new_n797), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G132), .A2(new_n787), .B1(new_n790), .B2(G50), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n329), .B1(new_n832), .B2(G150), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n804), .A2(G137), .B1(new_n777), .B2(G128), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1238), .B(new_n1242), .C1(new_n838), .C2(new_n1172), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n804), .A2(G283), .B1(new_n777), .B2(G303), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n329), .C1(new_n543), .C2(new_n772), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n837), .A2(new_n483), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n845), .A2(new_n1029), .B1(new_n448), .B2(new_n789), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n256), .A2(new_n779), .B1(new_n782), .B2(new_n1186), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n763), .B1(new_n1243), .B2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n751), .C1(G68), .C2(new_n1160), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1117), .B2(new_n760), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n749), .B(KEYINPUT122), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(new_n1151), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1237), .A2(new_n1254), .ZN(G381));
  OR2_X1    g1055(.A1(G393), .A2(G396), .ZN(new_n1256));
  OR4_X1    g1056(.A1(G384), .A2(G378), .A3(G381), .A4(new_n1256), .ZN(new_n1257));
  OR4_X1    g1057(.A1(G387), .A2(new_n1257), .A3(G390), .A4(G375), .ZN(G407));
  INV_X1    g1058(.A(G378), .ZN(new_n1259));
  INV_X1    g1059(.A(G343), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(G213), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT123), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G407), .B(G213), .C1(G375), .C2(new_n1263), .ZN(G409));
  INV_X1    g1064(.A(KEYINPUT124), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1220), .A2(new_n1221), .A3(new_n1217), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1218), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1235), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1265), .B1(new_n1268), .B2(new_n1230), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1232), .A2(new_n1227), .A3(KEYINPUT124), .A4(new_n1235), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1219), .B1(new_n1227), .B2(new_n1253), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1259), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G378), .B(new_n1228), .C1(new_n1231), .C2(new_n1233), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1262), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1262), .A2(G2897), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1236), .A2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1144), .A2(KEYINPUT60), .A3(new_n1146), .A4(new_n1133), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1153), .A3(new_n708), .A4(new_n1282), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1283), .A2(G384), .A3(new_n1254), .ZN(new_n1284));
  AOI21_X1  g1084(.A(G384), .B1(new_n1283), .B2(new_n1254), .ZN(new_n1285));
  OAI211_X1 g1085(.A(KEYINPUT125), .B(new_n1279), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1254), .ZN(new_n1287));
  INV_X1    g1087(.A(G384), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1283), .A2(G384), .A3(new_n1254), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1286), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1279), .B1(new_n1294), .B2(KEYINPUT125), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1277), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G387), .A2(G390), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G393), .A2(G396), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1256), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1040), .B1(new_n985), .B2(new_n1013), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1301), .B1(new_n1302), .B2(new_n1106), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1300), .A2(new_n1299), .A3(new_n1256), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1298), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1298), .B2(new_n1303), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1294), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1275), .A2(new_n1276), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT63), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1262), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(KEYINPUT63), .A3(new_n1308), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1297), .A2(new_n1307), .A3(new_n1311), .A4(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  OAI21_X1  g1115(.A(KEYINPUT125), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1278), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(new_n1286), .A3(new_n1292), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1315), .B1(new_n1318), .B2(new_n1312), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1309), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1312), .A2(KEYINPUT62), .A3(new_n1308), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1319), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1314), .B1(new_n1323), .B2(new_n1307), .ZN(G405));
  NAND2_X1  g1124(.A1(G375), .A2(new_n1259), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1274), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1308), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1326), .A2(new_n1308), .ZN(new_n1329));
  OAI22_X1  g1129(.A1(new_n1328), .A2(new_n1329), .B1(new_n1306), .B2(new_n1305), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1329), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1331), .A2(new_n1307), .A3(new_n1327), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1330), .A2(new_n1332), .ZN(G402));
endmodule


