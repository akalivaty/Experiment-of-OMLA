//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n588, new_n589,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  NAND2_X1  g034(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g037(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT67), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n469), .B1(new_n475), .B2(new_n478), .ZN(G160));
  AOI21_X1  g054(.A(new_n465), .B1(new_n462), .B2(new_n463), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(G136), .B2(new_n464), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n470), .A2(new_n486), .A3(G138), .A4(new_n465), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n465), .A2(G138), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n462), .B2(new_n463), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n489), .B2(new_n486), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT69), .A2(G114), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT69), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n480), .A2(G126), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(G62), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT72), .A2(G75), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(G651), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT73), .ZN(new_n511));
  AND3_X1   g086(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(G543), .B1(KEYINPUT70), .B2(KEYINPUT5), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT71), .B(G88), .ZN(new_n517));
  OAI21_X1  g092(.A(G543), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n522), .B(G651), .C1(new_n504), .C2(new_n509), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n511), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n520), .B1(KEYINPUT73), .B2(new_n510), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(KEYINPUT74), .A3(new_n523), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(G166));
  NAND2_X1  g104(.A1(new_n502), .A2(new_n503), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n516), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n518), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g114(.A(KEYINPUT75), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G51), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n537), .A2(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  OR2_X1    g119(.A1(KEYINPUT6), .A2(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(KEYINPUT6), .A2(G651), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n502), .A2(new_n503), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n541), .A2(G52), .B1(G90), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n549));
  INV_X1    g124(.A(G64), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n502), .B2(new_n503), .ZN(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n549), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n512), .A2(new_n513), .ZN(new_n555));
  OAI211_X1 g130(.A(KEYINPUT76), .B(new_n552), .C1(new_n555), .C2(new_n550), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n554), .A2(new_n556), .A3(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n548), .A2(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  AOI22_X1  g134(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G651), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT77), .B(G81), .Z(new_n562));
  OAI22_X1  g137(.A1(new_n560), .A2(new_n561), .B1(new_n516), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G43), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n539), .B2(new_n540), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT78), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n502), .B2(new_n503), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n573), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g153(.A(KEYINPUT79), .B(new_n576), .C1(new_n555), .C2(new_n574), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n578), .A2(new_n579), .A3(G651), .ZN(new_n580));
  INV_X1    g155(.A(G53), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT9), .B1(new_n518), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n545), .A2(new_n546), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT9), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n583), .A2(new_n584), .A3(G53), .A4(G543), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n582), .A2(new_n585), .B1(G91), .B2(new_n547), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n580), .A2(new_n586), .ZN(G299));
  AOI21_X1  g162(.A(KEYINPUT74), .B1(new_n527), .B2(new_n523), .ZN(new_n588));
  AND4_X1   g163(.A1(KEYINPUT74), .A2(new_n511), .A3(new_n521), .A4(new_n523), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n588), .A2(new_n589), .ZN(G303));
  NAND2_X1  g165(.A1(new_n547), .A2(G87), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n501), .B1(new_n545), .B2(new_n546), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G49), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n591), .A2(KEYINPUT80), .A3(new_n592), .A4(new_n594), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G288));
  AOI22_X1  g175(.A1(new_n530), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n561), .ZN(new_n602));
  INV_X1    g177(.A(G86), .ZN(new_n603));
  INV_X1    g178(.A(G48), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n516), .A2(new_n603), .B1(new_n518), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G305));
  NAND2_X1  g182(.A1(G72), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G60), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n555), .B2(new_n609), .ZN(new_n610));
  XOR2_X1   g185(.A(KEYINPUT81), .B(G85), .Z(new_n611));
  AOI22_X1  g186(.A1(new_n610), .A2(G651), .B1(new_n547), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n541), .A2(G47), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(G290));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n516), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n530), .A2(new_n583), .A3(KEYINPUT10), .A4(G92), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(KEYINPUT75), .B1(new_n583), .B2(G543), .ZN(new_n620));
  INV_X1    g195(.A(new_n540), .ZN(new_n621));
  OAI21_X1  g196(.A(G54), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(G66), .B1(new_n512), .B2(new_n513), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G651), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n619), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G171), .B2(new_n628), .ZN(G284));
  OAI21_X1  g205(.A(new_n629), .B1(G171), .B2(new_n628), .ZN(G321));
  NAND2_X1  g206(.A1(G299), .A2(new_n628), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G168), .B2(new_n628), .ZN(G297));
  OAI21_X1  g208(.A(new_n632), .B1(G168), .B2(new_n628), .ZN(G280));
  INV_X1    g209(.A(new_n627), .ZN(new_n635));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G860), .ZN(G148));
  OR2_X1    g212(.A1(new_n563), .A2(new_n565), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(new_n628), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n627), .A2(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(new_n628), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g217(.A1(new_n470), .A2(new_n467), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT12), .Z(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT13), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(new_n646));
  AOI22_X1  g221(.A1(G123), .A2(new_n480), .B1(new_n464), .B2(G135), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n649));
  INV_X1    g224(.A(G111), .ZN(new_n650));
  AOI22_X1  g225(.A1(new_n648), .A2(new_n649), .B1(new_n650), .B2(G2105), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n649), .B2(new_n648), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(G2096), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n646), .A2(new_n654), .ZN(G156));
  INV_X1    g230(.A(KEYINPUT14), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n658), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n661), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(G401));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  XOR2_X1   g246(.A(KEYINPUT84), .B(KEYINPUT17), .Z(new_n672));
  XNOR2_X1  g247(.A(G2072), .B(G2078), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT83), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n671), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(new_n673), .B2(new_n676), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT18), .Z(new_n680));
  INV_X1    g255(.A(new_n671), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n678), .B(new_n680), .C1(new_n674), .C2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2096), .B(G2100), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT85), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1961), .B(G1966), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(new_n688), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n690), .A2(new_n693), .ZN(new_n696));
  MUX2_X1   g271(.A(new_n688), .B(new_n695), .S(new_n696), .Z(new_n697));
  NOR2_X1   g272(.A1(new_n694), .A2(new_n688), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n697), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n701), .B1(new_n697), .B2(new_n700), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n686), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n704), .ZN(new_n706));
  INV_X1    g281(.A(new_n686), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n706), .A2(new_n707), .A3(new_n702), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1981), .B(G1986), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n705), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n705), .B2(new_n708), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(G229));
  NAND2_X1  g287(.A1(new_n606), .A2(G16), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G6), .B2(G16), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT32), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(KEYINPUT32), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G1981), .ZN(new_n718));
  INV_X1    g293(.A(G1981), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n715), .A2(new_n719), .A3(new_n716), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G22), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT91), .Z(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G166), .B2(new_n722), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G1971), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(G1971), .ZN(new_n727));
  NOR2_X1   g302(.A1(G16), .A2(G23), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT90), .Z(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n595), .B2(new_n722), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT33), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1976), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n721), .A2(new_n726), .A3(new_n727), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(KEYINPUT34), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT87), .B(G29), .Z(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G25), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n464), .A2(G131), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n480), .A2(G119), .ZN(new_n740));
  OR2_X1    g315(.A1(G95), .A2(G2105), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n741), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT88), .Z(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n738), .B1(new_n745), .B2(new_n737), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT35), .B(G1991), .Z(new_n747));
  XOR2_X1   g322(.A(new_n746), .B(new_n747), .Z(new_n748));
  NOR2_X1   g323(.A1(G16), .A2(G24), .ZN(new_n749));
  XOR2_X1   g324(.A(G290), .B(KEYINPUT89), .Z(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1986), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n733), .B2(KEYINPUT34), .ZN(new_n754));
  OAI21_X1  g329(.A(KEYINPUT36), .B1(new_n735), .B2(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n733), .A2(KEYINPUT34), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n756), .A2(new_n757), .A3(new_n734), .A4(new_n753), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT24), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(G34), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(G34), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n736), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G160), .ZN(new_n764));
  INV_X1    g339(.A(G29), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT94), .ZN(new_n767));
  INV_X1    g342(.A(G2084), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n722), .A2(G20), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT23), .Z(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G299), .B2(G16), .ZN(new_n773));
  INV_X1    g348(.A(G1956), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n769), .A2(new_n770), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(G162), .A2(new_n737), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n737), .A2(G35), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(KEYINPUT29), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT29), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n777), .A2(new_n781), .A3(new_n778), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G2090), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n566), .A2(G16), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G16), .B2(G19), .ZN(new_n787));
  INV_X1    g362(.A(G1341), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n765), .A2(G32), .ZN(new_n789));
  NAND3_X1  g364(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT95), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT26), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n464), .A2(G141), .B1(G105), .B2(new_n467), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n480), .A2(G129), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(G29), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT27), .B(G1996), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT96), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n787), .A2(new_n788), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n737), .A2(G27), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G164), .B2(new_n737), .ZN(new_n801));
  INV_X1    g376(.A(G2078), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n799), .B(new_n803), .C1(new_n788), .C2(new_n787), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n785), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n722), .A2(G5), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G171), .B2(new_n722), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1961), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT25), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n464), .A2(G139), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n810), .B(new_n811), .C1(new_n465), .C2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT93), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G29), .ZN(new_n815));
  NOR2_X1   g390(.A1(G29), .A2(G33), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT92), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G2072), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n808), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(G4), .A2(G16), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n635), .B2(G16), .ZN(new_n822));
  INV_X1    g397(.A(G1348), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n818), .B2(new_n819), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n722), .A2(G21), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G168), .B2(new_n722), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(G1966), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT30), .B(G28), .ZN(new_n829));
  OR2_X1    g404(.A1(KEYINPUT31), .A2(G11), .ZN(new_n830));
  NAND2_X1  g405(.A1(KEYINPUT31), .A2(G11), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n829), .A2(new_n765), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n653), .B2(new_n736), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n827), .B2(G1966), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n736), .A2(G26), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT28), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n464), .A2(G140), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n480), .A2(G128), .ZN(new_n839));
  OR2_X1    g414(.A1(G104), .A2(G2105), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n840), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n837), .B1(new_n842), .B2(G29), .ZN(new_n843));
  INV_X1    g418(.A(G2067), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n796), .A2(new_n798), .ZN(new_n846));
  NOR4_X1   g421(.A1(new_n825), .A2(new_n835), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n776), .A2(new_n805), .A3(new_n820), .A4(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT97), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n847), .A2(new_n805), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n851), .A2(KEYINPUT97), .A3(new_n776), .A4(new_n820), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n759), .A2(new_n853), .ZN(G311));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n759), .A2(new_n855), .A3(new_n853), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n759), .B2(new_n853), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(G150));
  XNOR2_X1  g433(.A(KEYINPUT99), .B(G93), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n547), .A2(new_n859), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(new_n561), .ZN(new_n862));
  INV_X1    g437(.A(G55), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n539), .B2(new_n540), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT100), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(G67), .B1(new_n512), .B2(new_n513), .ZN(new_n866));
  NAND2_X1  g441(.A1(G80), .A2(G543), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n868), .A2(G651), .B1(new_n547), .B2(new_n859), .ZN(new_n869));
  OAI21_X1  g444(.A(G55), .B1(new_n620), .B2(new_n621), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n865), .A2(new_n566), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n566), .B1(new_n865), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n635), .A2(G559), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n880));
  XNOR2_X1  g455(.A(KEYINPUT101), .B(G860), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n869), .B2(new_n870), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT37), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(G145));
  XOR2_X1   g460(.A(KEYINPUT105), .B(G37), .Z(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n464), .A2(G142), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n480), .A2(G130), .ZN(new_n889));
  OR2_X1    g464(.A1(G106), .A2(G2105), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n890), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n644), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n644), .A2(new_n892), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n894), .A2(new_n895), .A3(new_n743), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n743), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(KEYINPUT104), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n900));
  INV_X1    g475(.A(new_n743), .ZN(new_n901));
  INV_X1    g476(.A(new_n895), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(new_n893), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n900), .B1(new_n903), .B2(new_n896), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n907));
  INV_X1    g482(.A(new_n842), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n490), .A2(new_n496), .A3(KEYINPUT102), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT102), .B1(new_n490), .B2(new_n496), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n795), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n497), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n842), .A3(new_n909), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n913), .B1(new_n912), .B2(new_n916), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n907), .B(new_n813), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n912), .A2(new_n916), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n795), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n814), .A3(new_n917), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n917), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n907), .B1(new_n925), .B2(new_n813), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n906), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n813), .B1(new_n918), .B2(new_n919), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT103), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n929), .A2(new_n905), .A3(new_n923), .A4(new_n920), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(G162), .B(new_n653), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(G160), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n887), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n897), .B(new_n898), .C1(new_n924), .C2(new_n926), .ZN(new_n935));
  INV_X1    g510(.A(new_n933), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n930), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g514(.A1(G299), .A2(new_n627), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n541), .A2(G54), .B1(G651), .B2(new_n625), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n942), .A2(new_n580), .A3(new_n586), .A4(new_n619), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  XOR2_X1   g519(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n940), .B2(new_n943), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT107), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n940), .A2(new_n943), .ZN(new_n948));
  INV_X1    g523(.A(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n948), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n875), .B(new_n640), .ZN(new_n955));
  MUX2_X1   g530(.A(new_n953), .B(new_n954), .S(new_n955), .Z(new_n956));
  OR2_X1    g531(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n526), .A2(new_n528), .A3(G305), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n595), .ZN(new_n960));
  XNOR2_X1  g535(.A(G290), .B(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G305), .B1(new_n526), .B2(new_n528), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(G290), .B(new_n595), .ZN(new_n964));
  NAND2_X1  g539(.A1(G166), .A2(new_n606), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n964), .B1(new_n965), .B2(new_n958), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n957), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n957), .B2(new_n968), .ZN(new_n970));
  OAI21_X1  g545(.A(G868), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n628), .B1(new_n862), .B2(new_n864), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(G295));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n972), .ZN(G331));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n975));
  NAND2_X1  g550(.A1(G301), .A2(G286), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n548), .A2(new_n537), .A3(new_n542), .A4(new_n557), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n873), .B2(new_n874), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n862), .A2(KEYINPUT100), .A3(new_n864), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n871), .B1(new_n869), .B2(new_n870), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n638), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n865), .A2(new_n566), .A3(new_n872), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n983), .A3(new_n976), .A4(new_n977), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n984), .A3(new_n954), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n965), .A2(new_n964), .A3(new_n958), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n961), .B1(new_n959), .B2(new_n962), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n947), .A2(new_n952), .B1(new_n984), .B2(new_n979), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n975), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n979), .A2(new_n984), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n940), .A2(new_n943), .A3(new_n941), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n951), .B1(new_n950), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n946), .A2(KEYINPUT107), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n995), .A2(new_n967), .A3(KEYINPUT108), .A4(new_n985), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n990), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n985), .ZN(new_n998));
  INV_X1    g573(.A(new_n967), .ZN(new_n999));
  AOI21_X1  g574(.A(G37), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n991), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n948), .A2(new_n941), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n948), .B2(new_n945), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n985), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n887), .B1(new_n1006), .B2(new_n999), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n997), .A2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT44), .B(new_n1002), .C1(new_n1008), .C2(new_n1001), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n997), .A2(new_n1000), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT109), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1001), .B1(new_n997), .B2(new_n1000), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n997), .A2(new_n1001), .A3(new_n1007), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT110), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1016), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1020));
  AOI211_X1 g595(.A(KEYINPUT109), .B(new_n1001), .C1(new_n997), .C2(new_n1000), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT110), .B(new_n1018), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1009), .B1(new_n1019), .B2(new_n1023), .ZN(G397));
  NOR2_X1   g599(.A1(new_n476), .A2(new_n477), .ZN(new_n1025));
  AOI211_X1 g600(.A(KEYINPUT67), .B(new_n465), .C1(new_n471), .C2(new_n472), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n468), .B(G40), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1384), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT45), .B1(new_n497), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(G1384), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n915), .A2(new_n909), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1030), .A2(new_n802), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1027), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n497), .B2(new_n1028), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI211_X1 g614(.A(KEYINPUT50), .B(G1384), .C1(new_n490), .C2(new_n496), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1036), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1961), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1034), .A2(new_n1035), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n497), .A2(KEYINPUT117), .A3(new_n1032), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT117), .B1(new_n497), .B2(new_n1032), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1030), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1044), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(G301), .B(KEYINPUT54), .ZN(new_n1051));
  INV_X1    g626(.A(G40), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n476), .A2(new_n1052), .A3(new_n1049), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1033), .A2(new_n468), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n915), .A2(new_n1028), .A3(new_n909), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1031), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1051), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1050), .A2(new_n1051), .B1(new_n1057), .B2(new_n1044), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1042), .A2(G2084), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1966), .B1(new_n1047), .B2(new_n1030), .ZN(new_n1060));
  OAI211_X1 g635(.A(G8), .B(G286), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1060), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1027), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n768), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1062), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G168), .A2(new_n1062), .ZN(new_n1067));
  XOR2_X1   g642(.A(new_n1067), .B(KEYINPUT124), .Z(new_n1068));
  OAI211_X1 g643(.A(new_n1061), .B(KEYINPUT51), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(G8), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1067), .A2(KEYINPUT51), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1058), .A2(new_n1069), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n960), .A2(G1976), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n497), .A2(new_n1028), .ZN(new_n1075));
  OAI211_X1 g650(.A(G8), .B(new_n1074), .C1(new_n1027), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1976), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n597), .A2(new_n1078), .A3(new_n598), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1079), .A2(KEYINPUT114), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT114), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1077), .B(KEYINPUT115), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n1076), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n1087));
  OAI21_X1  g662(.A(G1981), .B1(new_n602), .B2(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1088), .A2(new_n606), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n606), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT49), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n1027), .B2(new_n1075), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(KEYINPUT49), .A3(new_n1090), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1076), .A2(KEYINPUT52), .ZN(new_n1096));
  AND4_X1   g671(.A1(new_n1083), .A2(new_n1086), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1098));
  INV_X1    g673(.A(G1971), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1064), .A2(new_n784), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1062), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(G303), .B(G8), .C1(KEYINPUT112), .C2(KEYINPUT55), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(G166), .B2(new_n1062), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT113), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1103), .A2(new_n1109), .A3(new_n1105), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1102), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1097), .A2(new_n1108), .A3(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1073), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G1996), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1030), .A2(new_n1116), .A3(new_n1033), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(G1341), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1027), .B2(new_n1075), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n638), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1121), .B(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(G299), .B(KEYINPUT57), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT119), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1042), .A2(new_n774), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT56), .B(G2072), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1030), .A2(new_n1033), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1125), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1124), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1126), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1130), .A2(KEYINPUT61), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(KEYINPUT121), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1131), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1129), .A2(new_n1137), .A3(new_n1124), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1123), .B(new_n1133), .C1(new_n1136), .C2(new_n1140), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1027), .A2(G2067), .A3(new_n1075), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1042), .B2(new_n823), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT60), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(new_n627), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n627), .B(KEYINPUT122), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1143), .A2(KEYINPUT60), .A3(new_n1147), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1143), .A2(KEYINPUT60), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT123), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1146), .A2(new_n1149), .A3(new_n1152), .A4(new_n1148), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1141), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1143), .A2(new_n627), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1132), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1130), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1115), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1069), .A2(new_n1159), .A3(new_n1072), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1112), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n1110), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1107), .B1(new_n1164), .B2(new_n1102), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1165), .A2(G171), .A3(new_n1097), .A4(new_n1050), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT125), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1070), .A2(G286), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1097), .A2(new_n1108), .A3(new_n1113), .A4(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT63), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1165), .A2(new_n1172), .A3(new_n1097), .A4(new_n1168), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1095), .A2(new_n1078), .A3(new_n599), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n606), .A2(new_n719), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1092), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1113), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1176), .B1(new_n1177), .B2(new_n1097), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1171), .A2(new_n1173), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1050), .A2(G171), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1114), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1181), .B(new_n1182), .C1(new_n1161), .C2(new_n1160), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1158), .A2(new_n1167), .A3(new_n1179), .A4(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1056), .A2(new_n1027), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1185), .A2(G1996), .A3(new_n795), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT111), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n842), .B(new_n844), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(G1996), .B2(new_n795), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1187), .B1(new_n1185), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1185), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n743), .B(new_n747), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g768(.A(G290), .B(G1986), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1193), .B1(new_n1185), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1184), .A2(new_n1195), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1191), .A2(G1986), .A3(G290), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT48), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1185), .A2(new_n1116), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT46), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT126), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT47), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n913), .A2(new_n1188), .ZN(new_n1204));
  AOI22_X1  g779(.A1(new_n1199), .A2(new_n1200), .B1(new_n1185), .B2(new_n1204), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1203), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1207));
  OAI22_X1  g782(.A1(new_n1193), .A2(new_n1198), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1190), .A2(new_n747), .A3(new_n745), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n908), .A2(new_n844), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1191), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1196), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g788(.A(G319), .ZN(new_n1215));
  NOR3_X1   g789(.A1(G401), .A2(new_n1215), .A3(G227), .ZN(new_n1216));
  OAI21_X1  g790(.A(new_n1216), .B1(new_n710), .B2(new_n711), .ZN(new_n1217));
  AOI21_X1  g791(.A(new_n1217), .B1(new_n934), .B2(new_n937), .ZN(new_n1218));
  OAI21_X1  g792(.A(new_n1218), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n1219), .A2(KEYINPUT127), .ZN(new_n1220));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n1221));
  NAND3_X1  g795(.A1(new_n1017), .A2(new_n1221), .A3(new_n1218), .ZN(new_n1222));
  AND2_X1   g796(.A1(new_n1220), .A2(new_n1222), .ZN(G308));
  NAND2_X1  g797(.A1(new_n1220), .A2(new_n1222), .ZN(G225));
endmodule


