//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(G127gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(G127gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n206), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G155gat), .ZN(new_n214));
  INV_X1    g013(.A(G162gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT78), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n218), .B1(G155gat), .B2(G162gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G155gat), .B(G162gat), .Z(new_n221));
  AND2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n220), .B(new_n221), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n208), .A2(new_n212), .A3(new_n226), .ZN(new_n231));
  XOR2_X1   g030(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(KEYINPUT4), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n231), .A2(KEYINPUT4), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT81), .B1(new_n238), .B2(new_n233), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n230), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT5), .ZN(new_n241));
  NAND2_X1  g040(.A1(G225gat), .A2(G233gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n213), .A2(new_n224), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n231), .ZN(new_n245));
  INV_X1    g044(.A(new_n242), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n208), .A2(new_n212), .A3(new_n226), .A4(KEYINPUT4), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n229), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n232), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n246), .B1(new_n231), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT80), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  AND4_X1   g051(.A1(KEYINPUT80), .A2(new_n251), .A3(new_n248), .A4(new_n229), .ZN(new_n253));
  OAI211_X1 g052(.A(KEYINPUT5), .B(new_n247), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n243), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G1gat), .B(G29gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT0), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(G57gat), .ZN(new_n259));
  INV_X1    g058(.A(G85gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT6), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n261), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n255), .A2(KEYINPUT6), .A3(new_n263), .ZN(new_n266));
  XNOR2_X1  g065(.A(G211gat), .B(G218gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT75), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n269));
  INV_X1    g068(.A(G197gat), .ZN(new_n270));
  INV_X1    g069(.A(G204gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G197gat), .A2(G204gat), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n268), .B(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT25), .ZN(new_n278));
  XOR2_X1   g077(.A(G183gat), .B(G190gat), .Z(new_n279));
  INV_X1    g078(.A(KEYINPUT24), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT66), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI22_X1  g087(.A1(KEYINPUT65), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n281), .A2(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n282), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n291), .B(KEYINPUT24), .ZN(new_n294));
  INV_X1    g093(.A(G183gat), .ZN(new_n295));
  INV_X1    g094(.A(G190gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT64), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT64), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n294), .A2(new_n300), .A3(new_n297), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n290), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n293), .B1(new_n302), .B2(new_n278), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n305));
  NAND2_X1  g104(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT27), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(KEYINPUT67), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n295), .A2(KEYINPUT27), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n306), .A2(new_n308), .B1(new_n309), .B2(KEYINPUT67), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n311), .A2(new_n296), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n305), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT27), .B(G183gat), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n296), .A2(KEYINPUT28), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT70), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT67), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n306), .A2(new_n320), .A3(KEYINPUT27), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT67), .B1(new_n307), .B2(G183gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n311), .A2(new_n296), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n319), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT70), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n316), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n318), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT26), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n283), .B1(new_n286), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT71), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n286), .A2(new_n329), .ZN(new_n333));
  OAI211_X1 g132(.A(KEYINPUT71), .B(new_n283), .C1(new_n286), .C2(new_n329), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n335), .A2(new_n291), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT72), .B1(new_n328), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n291), .ZN(new_n339));
  AOI211_X1 g138(.A(new_n338), .B(new_n339), .C1(new_n318), .C2(new_n327), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n304), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT76), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n321), .A2(new_n322), .A3(new_n296), .A4(new_n311), .ZN(new_n343));
  AOI221_X4 g142(.A(KEYINPUT70), .B1(new_n314), .B2(new_n315), .C1(new_n343), .C2(new_n319), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n326), .B1(new_n325), .B2(new_n316), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n336), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n338), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n336), .B(KEYINPUT72), .C1(new_n344), .C2(new_n345), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n304), .ZN(new_n351));
  AOI211_X1 g150(.A(KEYINPUT29), .B(new_n277), .C1(new_n342), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n304), .A2(new_n346), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(new_n276), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n275), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n277), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n350), .B1(new_n349), .B2(new_n304), .ZN(new_n358));
  AOI211_X1 g157(.A(KEYINPUT76), .B(new_n303), .C1(new_n347), .C2(new_n348), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n277), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(KEYINPUT77), .B(new_n277), .C1(new_n358), .C2(new_n359), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n357), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n355), .B1(new_n364), .B2(new_n275), .ZN(new_n365));
  XOR2_X1   g164(.A(G8gat), .B(G36gat), .Z(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(G64gat), .ZN(new_n367));
  INV_X1    g166(.A(G92gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n265), .A2(new_n266), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n357), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n342), .A2(new_n351), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT77), .B1(new_n374), .B2(new_n277), .ZN(new_n375));
  INV_X1    g174(.A(new_n363), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(KEYINPUT86), .A3(new_n275), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT86), .ZN(new_n379));
  INV_X1    g178(.A(new_n275), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n379), .B1(new_n364), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n380), .B1(new_n352), .B2(new_n354), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT37), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT37), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n370), .B1(new_n365), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT38), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n277), .A2(KEYINPUT29), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n354), .B1(new_n374), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(new_n380), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n377), .B2(new_n380), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT37), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(KEYINPUT38), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n372), .B1(new_n387), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n369), .B(new_n355), .C1(new_n364), .C2(new_n275), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n371), .A2(KEYINPUT30), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n244), .A2(new_n242), .A3(new_n231), .ZN(new_n398));
  OAI211_X1 g197(.A(KEYINPUT39), .B(new_n398), .C1(new_n240), .C2(new_n242), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n235), .B1(new_n234), .B2(new_n236), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n238), .A2(new_n233), .A3(KEYINPUT81), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n229), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT39), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(new_n403), .A3(new_n246), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n399), .A2(new_n261), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n264), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n405), .A2(new_n406), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n365), .A2(new_n411), .A3(new_n370), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n227), .B1(new_n275), .B2(KEYINPUT29), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n224), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n228), .A2(new_n356), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n275), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT83), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G228gat), .A2(G233gat), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  OR3_X1    g221(.A1(new_n421), .A2(new_n422), .A3(G22gat), .ZN(new_n423));
  OAI21_X1  g222(.A(G22gat), .B1(new_n421), .B2(new_n422), .ZN(new_n424));
  XOR2_X1   g223(.A(G78gat), .B(G106gat), .Z(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT31), .ZN(new_n426));
  INV_X1    g225(.A(G50gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AND4_X1   g228(.A1(new_n414), .A2(new_n423), .A3(new_n424), .A4(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n423), .B2(new_n424), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n424), .A2(new_n414), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n413), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n395), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n341), .A2(new_n213), .ZN(new_n436));
  NAND2_X1  g235(.A1(G227gat), .A2(G233gat), .ZN(new_n437));
  INV_X1    g236(.A(new_n213), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n349), .A2(new_n438), .A3(new_n304), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT73), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT34), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n440), .B2(KEYINPUT34), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n437), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n438), .B1(new_n349), .B2(new_n304), .ZN(new_n447));
  AOI211_X1 g246(.A(new_n213), .B(new_n303), .C1(new_n347), .C2(new_n348), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450));
  XNOR2_X1  g249(.A(G15gat), .B(G43gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(G71gat), .ZN(new_n452));
  INV_X1    g251(.A(G99gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n449), .B(KEYINPUT32), .C1(new_n450), .C2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n449), .B2(new_n450), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n449), .A2(KEYINPUT32), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n447), .A2(new_n448), .A3(new_n446), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT34), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n445), .A2(new_n456), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n456), .ZN(new_n464));
  INV_X1    g263(.A(new_n444), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(new_n462), .A3(new_n442), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT36), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n466), .A2(KEYINPUT74), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n468), .B2(KEYINPUT74), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n473), .B2(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n397), .A2(new_n412), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n264), .A2(KEYINPUT82), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n255), .A2(new_n477), .A3(new_n263), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n262), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n266), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n433), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n377), .A2(new_n380), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n369), .B1(new_n483), .B2(new_n355), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n396), .A2(KEYINPUT30), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n412), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n480), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n464), .A2(new_n466), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n445), .A2(new_n462), .B1(new_n456), .B2(new_n459), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT74), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n472), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n433), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT35), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT35), .B1(new_n265), .B2(new_n266), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n475), .A2(new_n495), .A3(new_n433), .A4(new_n469), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n435), .A2(new_n482), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G8gat), .ZN(new_n498));
  XOR2_X1   g297(.A(G15gat), .B(G22gat), .Z(new_n499));
  INV_X1    g298(.A(G1gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT16), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(G1gat), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n501), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n503), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT87), .B(G36gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(G29gat), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR3_X1   g311(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(G43gat), .B(G50gat), .Z(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(KEYINPUT15), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT88), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n519), .B(KEYINPUT15), .Z(new_n520));
  NAND2_X1  g319(.A1(new_n511), .A2(KEYINPUT89), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT90), .ZN(new_n522));
  INV_X1    g321(.A(new_n513), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n523), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n510), .B(KEYINPUT91), .Z(new_n526));
  NAND4_X1  g325(.A1(new_n520), .A2(new_n524), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n508), .B1(new_n517), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n527), .A2(KEYINPUT17), .A3(new_n517), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT17), .B1(new_n527), .B2(new_n517), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n528), .B1(new_n531), .B2(new_n508), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT18), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n527), .A2(new_n517), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT93), .B1(new_n537), .B2(new_n507), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n538), .A2(new_n528), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n533), .B(KEYINPUT13), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n528), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n532), .A2(KEYINPUT18), .A3(new_n533), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n536), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(G197gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT11), .ZN(new_n547));
  INV_X1    g346(.A(G169gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT12), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n536), .A2(new_n542), .A3(new_n550), .A4(new_n543), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(KEYINPUT94), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n544), .A2(new_n555), .A3(new_n551), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n497), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(KEYINPUT41), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G134gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G190gat), .B(G218gat), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT102), .ZN(new_n565));
  NAND2_X1  g364(.A1(G85gat), .A2(G92gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n566), .B(new_n567), .Z(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n569), .B1(new_n260), .B2(new_n368), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT100), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT100), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n568), .A2(new_n575), .A3(new_n572), .A4(new_n570), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(KEYINPUT101), .A3(new_n576), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n529), .A2(new_n530), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n576), .ZN(new_n579));
  NOR2_X1   g378(.A1(KEYINPUT101), .A2(KEYINPUT17), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(new_n537), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n560), .A2(KEYINPUT41), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n565), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(G162gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n584), .A2(G162gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n564), .A2(KEYINPUT102), .ZN(new_n588));
  NOR3_X1   g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n584), .A2(G162gat), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n590), .B1(new_n591), .B2(new_n585), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n563), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n588), .B1(new_n586), .B2(new_n587), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n590), .A3(new_n585), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n562), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G57gat), .B(G64gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(KEYINPUT95), .Z(new_n599));
  NAND2_X1  g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  OR2_X1    g399(.A1(G71gat), .A2(G78gat), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT9), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n600), .B(new_n601), .C1(new_n598), .C2(new_n602), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n507), .B1(new_n607), .B2(KEYINPUT21), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT97), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G127gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n609), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT98), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT96), .B(G155gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n618), .B(new_n619), .Z(new_n620));
  NAND2_X1  g419(.A1(new_n612), .A2(new_n616), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n620), .B1(new_n617), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT103), .Z(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n607), .B1(new_n574), .B2(new_n576), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n573), .A2(new_n606), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n579), .A2(KEYINPUT10), .A3(new_n607), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n626), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n628), .A2(new_n633), .A3(new_n629), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT105), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT104), .ZN(new_n639));
  INV_X1    g438(.A(G176gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(new_n271), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n637), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n597), .A2(new_n624), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT106), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n558), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n266), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n477), .B1(new_n255), .B2(new_n263), .ZN(new_n650));
  AOI211_X1 g449(.A(KEYINPUT82), .B(new_n261), .C1(new_n243), .C2(new_n254), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n652), .B2(new_n262), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  INV_X1    g454(.A(new_n475), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n504), .A2(new_n498), .ZN(new_n657));
  NAND2_X1  g456(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n648), .A2(new_n656), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n648), .ZN(new_n664));
  OAI21_X1  g463(.A(G8gat), .B1(new_n664), .B2(new_n475), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT42), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT107), .B1(new_n666), .B2(new_n659), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n663), .B1(new_n667), .B2(new_n661), .ZN(G1325gat));
  AND3_X1   g467(.A1(new_n648), .A2(G15gat), .A3(new_n474), .ZN(new_n669));
  AOI21_X1  g468(.A(G15gat), .B1(new_n648), .B2(new_n469), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(G1326gat));
  INV_X1    g470(.A(new_n433), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n648), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  NAND2_X1  g474(.A1(new_n494), .A2(new_n496), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n413), .A2(new_n433), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n369), .B1(new_n391), .B2(KEYINPUT37), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(KEYINPUT37), .B2(new_n383), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n393), .B1(new_n679), .B2(KEYINPUT38), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n677), .B1(new_n680), .B2(new_n372), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n491), .A2(new_n492), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT36), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n653), .B1(new_n412), .B2(new_n397), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n683), .B(new_n471), .C1(new_n684), .C2(new_n433), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n676), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n597), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n624), .A2(new_n557), .A3(new_n644), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n691), .A2(G29gat), .A3(new_n480), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT45), .Z(new_n693));
  OAI21_X1  g492(.A(KEYINPUT44), .B1(new_n497), .B2(new_n597), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n686), .A2(new_n695), .A3(new_n687), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n690), .ZN(new_n698));
  OAI21_X1  g497(.A(G29gat), .B1(new_n698), .B2(new_n480), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n693), .A2(new_n699), .ZN(G1328gat));
  OR2_X1    g499(.A1(new_n691), .A2(new_n509), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n702));
  OAI22_X1  g501(.A1(new_n701), .A2(new_n475), .B1(new_n702), .B2(KEYINPUT46), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(KEYINPUT108), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n509), .B1(new_n698), .B2(new_n475), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n702), .B(KEYINPUT46), .C1(new_n701), .C2(new_n475), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(G1329gat));
  INV_X1    g507(.A(new_n474), .ZN(new_n709));
  OAI21_X1  g508(.A(G43gat), .B1(new_n698), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(G43gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n469), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n691), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1330gat));
  NOR3_X1   g514(.A1(new_n691), .A2(G50gat), .A3(new_n433), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n697), .A2(new_n672), .A3(new_n690), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(G50gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT48), .ZN(G1331gat));
  OR2_X1    g518(.A1(new_n622), .A2(new_n623), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n687), .A2(new_n720), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n686), .A2(new_n721), .A3(new_n557), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n480), .A2(new_n645), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT109), .B(G57gat), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1332gat));
  NOR2_X1   g525(.A1(new_n475), .A2(new_n645), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT49), .B(G64gat), .Z(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(G1333gat));
  NAND2_X1  g530(.A1(new_n722), .A2(new_n644), .ZN(new_n732));
  OAI21_X1  g531(.A(G71gat), .B1(new_n732), .B2(new_n709), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n732), .A2(G71gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(new_n468), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1334gat));
  NOR2_X1   g536(.A1(new_n433), .A2(new_n645), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G78gat), .ZN(G1335gat));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  INV_X1    g540(.A(new_n557), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n624), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n741), .B1(new_n688), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n686), .A2(KEYINPUT51), .A3(new_n687), .A4(new_n743), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(G85gat), .B1(new_n747), .B2(new_n723), .ZN(new_n748));
  AOI211_X1 g547(.A(new_n645), .B(new_n744), .C1(new_n694), .C2(new_n696), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n480), .A2(new_n260), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(G1336gat));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n697), .A2(new_n644), .A3(new_n656), .A4(new_n743), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G92gat), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n747), .A2(new_n368), .A3(new_n727), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n756), .B(new_n758), .ZN(G1337gat));
  NAND3_X1  g558(.A1(new_n469), .A2(new_n453), .A3(new_n644), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT111), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n747), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n749), .A2(new_n474), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(new_n453), .ZN(G1338gat));
  AOI21_X1  g563(.A(G106gat), .B1(new_n745), .B2(new_n746), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n765), .A2(new_n738), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n497), .A2(KEYINPUT44), .A3(new_n597), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n695), .B1(new_n686), .B2(new_n687), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n738), .B(new_n743), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT53), .B1(new_n766), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n697), .A2(KEYINPUT112), .A3(new_n738), .A4(new_n743), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(G106gat), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT53), .B1(new_n765), .B2(new_n738), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n771), .B1(new_n778), .B2(new_n779), .ZN(G1339gat));
  NOR2_X1   g579(.A1(new_n532), .A2(new_n533), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n549), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n553), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n630), .A2(new_n631), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n633), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n630), .A2(new_n626), .A3(new_n631), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(KEYINPUT54), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n643), .B1(new_n632), .B2(new_n789), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n788), .A2(KEYINPUT55), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT55), .B1(new_n788), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n635), .A2(new_n642), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n593), .A2(new_n784), .A3(new_n596), .A4(new_n794), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n795), .A2(KEYINPUT114), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n554), .A2(new_n556), .A3(new_n794), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n644), .A2(new_n784), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n597), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n795), .A2(KEYINPUT114), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n796), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n720), .ZN(new_n803));
  NOR4_X1   g602(.A1(new_n742), .A2(new_n687), .A3(new_n720), .A4(new_n644), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(new_n433), .A3(new_n469), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n656), .A2(new_n480), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G113gat), .B1(new_n810), .B2(new_n557), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n804), .B1(new_n802), .B2(new_n720), .ZN(new_n812));
  NOR4_X1   g611(.A1(new_n812), .A2(new_n480), .A3(new_n656), .A4(new_n493), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(new_n204), .A3(new_n742), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(G1340gat));
  OAI21_X1  g614(.A(G120gat), .B1(new_n810), .B2(new_n645), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n813), .A2(new_n202), .A3(new_n644), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1341gat));
  NOR3_X1   g617(.A1(new_n810), .A2(new_n209), .A3(new_n720), .ZN(new_n819));
  AOI21_X1  g618(.A(G127gat), .B1(new_n813), .B2(new_n624), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(G1342gat));
  NAND3_X1  g620(.A1(new_n813), .A2(new_n211), .A3(new_n687), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n822), .A2(KEYINPUT56), .ZN(new_n823));
  OAI21_X1  g622(.A(G134gat), .B1(new_n810), .B2(new_n597), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(KEYINPUT56), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT115), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n823), .A2(new_n828), .A3(new_n824), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(G1343gat));
  NAND2_X1  g629(.A1(new_n709), .A2(new_n809), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n812), .B2(new_n433), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n795), .B(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n624), .B1(new_n835), .B2(new_n800), .ZN(new_n836));
  OAI211_X1 g635(.A(KEYINPUT57), .B(new_n672), .C1(new_n836), .C2(new_n804), .ZN(new_n837));
  AOI211_X1 g636(.A(new_n557), .B(new_n831), .C1(new_n833), .C2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(G141gat), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT116), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT58), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n806), .A2(KEYINPUT117), .A3(new_n653), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n812), .B2(new_n480), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n709), .A2(new_n672), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n656), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n843), .A2(new_n845), .A3(new_n742), .A4(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n842), .B1(new_n848), .B2(G141gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n837), .ZN(new_n850));
  INV_X1    g649(.A(new_n831), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n742), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n853), .A3(G141gat), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n843), .A2(new_n845), .A3(new_n847), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n855), .A2(new_n841), .A3(new_n839), .A4(new_n742), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n849), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT58), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n838), .A2(new_n839), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n859), .A2(new_n849), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1344gat));
  INV_X1    g660(.A(G148gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n855), .A2(new_n862), .A3(new_n644), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n593), .A2(new_n596), .A3(new_n794), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(KEYINPUT121), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(KEYINPUT121), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n784), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n800), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n869), .A2(new_n720), .B1(new_n647), .B2(new_n557), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n832), .B1(new_n870), .B2(new_n433), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n837), .A2(KEYINPUT120), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n806), .A2(new_n873), .A3(KEYINPUT57), .A4(new_n672), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n831), .B(KEYINPUT119), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n644), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n864), .B1(new_n877), .B2(G148gat), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n831), .B1(new_n833), .B2(new_n837), .ZN(new_n879));
  AOI211_X1 g678(.A(KEYINPUT59), .B(new_n862), .C1(new_n879), .C2(new_n644), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n863), .B1(new_n878), .B2(new_n880), .ZN(G1345gat));
  AOI21_X1  g680(.A(G155gat), .B1(new_n855), .B2(new_n624), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n720), .A2(new_n214), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n879), .B2(new_n883), .ZN(G1346gat));
  AOI21_X1  g683(.A(G162gat), .B1(new_n855), .B2(new_n687), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n597), .A2(new_n215), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n879), .B2(new_n886), .ZN(G1347gat));
  NAND2_X1  g686(.A1(new_n656), .A2(new_n480), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT122), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n808), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G169gat), .B1(new_n890), .B2(new_n557), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n812), .A2(new_n653), .A3(new_n493), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n656), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n742), .A2(new_n548), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(G1348gat));
  OAI21_X1  g694(.A(G176gat), .B1(new_n890), .B2(new_n645), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n640), .A3(new_n727), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1349gat));
  NAND4_X1  g697(.A1(new_n892), .A2(new_n624), .A3(new_n314), .A4(new_n656), .ZN(new_n899));
  INV_X1    g698(.A(new_n889), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n807), .A2(new_n720), .A3(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n899), .B(KEYINPUT124), .C1(new_n901), .C2(new_n295), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT60), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n899), .B1(new_n901), .B2(new_n295), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n906), .B(new_n907), .C1(new_n903), .C2(new_n908), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n890), .B2(new_n597), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(KEYINPUT61), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(KEYINPUT61), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n687), .A2(new_n296), .ZN(new_n913));
  OAI22_X1  g712(.A1(new_n911), .A2(new_n912), .B1(new_n893), .B2(new_n913), .ZN(G1351gat));
  NOR2_X1   g713(.A1(new_n900), .A2(new_n474), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n875), .A2(new_n742), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G197gat), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n846), .A2(new_n475), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT125), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n812), .A2(new_n653), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n270), .A3(new_n742), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT126), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n917), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1352gat));
  XNOR2_X1  g727(.A(KEYINPUT127), .B(G204gat), .ZN(new_n929));
  OR3_X1    g728(.A1(new_n921), .A2(new_n645), .A3(new_n929), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n875), .A2(new_n644), .A3(new_n915), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(G1353gat));
  OR3_X1    g734(.A1(new_n921), .A2(G211gat), .A3(new_n720), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n875), .A2(new_n624), .A3(new_n915), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n937), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT63), .B1(new_n937), .B2(G211gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1354gat));
  AOI21_X1  g739(.A(G218gat), .B1(new_n922), .B2(new_n687), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n875), .A2(new_n915), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n687), .A2(G218gat), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(G1355gat));
endmodule


