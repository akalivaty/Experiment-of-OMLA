

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U550 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U551 ( .A1(n525), .A2(n524), .ZN(G160) );
  XNOR2_X2 U552 ( .A(n628), .B(n627), .ZN(n763) );
  NOR2_X1 U553 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U554 ( .A(n594), .B(n593), .ZN(n595) );
  NOR2_X1 U555 ( .A1(n720), .A2(n604), .ZN(n638) );
  NAND2_X1 U556 ( .A1(G160), .A2(G40), .ZN(n720) );
  NOR2_X2 U557 ( .A1(G2104), .A2(n521), .ZN(n873) );
  XNOR2_X1 U558 ( .A(KEYINPUT30), .B(KEYINPUT96), .ZN(n593) );
  XNOR2_X1 U559 ( .A(KEYINPUT32), .B(KEYINPUT102), .ZN(n666) );
  XNOR2_X1 U560 ( .A(n667), .B(n666), .ZN(n687) );
  NAND2_X1 U561 ( .A1(G8), .A2(n629), .ZN(n695) );
  AND2_X2 U562 ( .A1(n521), .A2(G2104), .ZN(n878) );
  NOR2_X1 U563 ( .A1(G651), .A2(n565), .ZN(n780) );
  NOR2_X1 U564 ( .A1(G651), .A2(G543), .ZN(n784) );
  INV_X1 U565 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U566 ( .A1(G101), .A2(n878), .ZN(n516) );
  XNOR2_X1 U567 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n514) );
  XNOR2_X1 U568 ( .A(n514), .B(KEYINPUT64), .ZN(n515) );
  XNOR2_X1 U569 ( .A(n516), .B(n515), .ZN(n519) );
  AND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n872) );
  NAND2_X1 U571 ( .A1(G113), .A2(n872), .ZN(n517) );
  XNOR2_X1 U572 ( .A(n517), .B(KEYINPUT66), .ZN(n518) );
  NAND2_X1 U573 ( .A1(n519), .A2(n518), .ZN(n525) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n520), .Z(n880) );
  NAND2_X1 U576 ( .A1(G137), .A2(n880), .ZN(n523) );
  NAND2_X1 U577 ( .A1(G125), .A2(n873), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U579 ( .A1(n784), .A2(G89), .ZN(n526) );
  XNOR2_X1 U580 ( .A(n526), .B(KEYINPUT4), .ZN(n528) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n565) );
  INV_X1 U582 ( .A(G651), .ZN(n530) );
  NOR2_X1 U583 ( .A1(n565), .A2(n530), .ZN(n785) );
  NAND2_X1 U584 ( .A1(G76), .A2(n785), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U586 ( .A(n529), .B(KEYINPUT5), .ZN(n536) );
  NAND2_X1 U587 ( .A1(G51), .A2(n780), .ZN(n533) );
  NOR2_X1 U588 ( .A1(G543), .A2(n530), .ZN(n531) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n531), .Z(n781) );
  NAND2_X1 U590 ( .A1(G63), .A2(n781), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U592 ( .A(KEYINPUT6), .B(n534), .Z(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U594 ( .A(n537), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U595 ( .A1(G90), .A2(n784), .ZN(n539) );
  NAND2_X1 U596 ( .A1(G77), .A2(n785), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U598 ( .A(KEYINPUT9), .B(n540), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n780), .A2(G52), .ZN(n542) );
  NAND2_X1 U600 ( .A1(G64), .A2(n781), .ZN(n541) );
  AND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(G301) );
  NAND2_X1 U603 ( .A1(G78), .A2(n785), .ZN(n545) );
  XOR2_X1 U604 ( .A(KEYINPUT68), .B(n545), .Z(n550) );
  NAND2_X1 U605 ( .A1(G53), .A2(n780), .ZN(n547) );
  NAND2_X1 U606 ( .A1(G65), .A2(n781), .ZN(n546) );
  NAND2_X1 U607 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U608 ( .A(KEYINPUT69), .B(n548), .Z(n549) );
  NOR2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n784), .A2(G91), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(G299) );
  XOR2_X1 U612 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U613 ( .A1(n780), .A2(G50), .ZN(n553) );
  XNOR2_X1 U614 ( .A(KEYINPUT78), .B(n553), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n781), .A2(G62), .ZN(n554) );
  XOR2_X1 U616 ( .A(KEYINPUT77), .B(n554), .Z(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U618 ( .A(KEYINPUT79), .B(n557), .ZN(n561) );
  NAND2_X1 U619 ( .A1(G88), .A2(n784), .ZN(n559) );
  NAND2_X1 U620 ( .A1(G75), .A2(n785), .ZN(n558) );
  AND2_X1 U621 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U622 ( .A1(n561), .A2(n560), .ZN(G303) );
  NAND2_X1 U623 ( .A1(G49), .A2(n780), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G74), .A2(G651), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U626 ( .A1(n781), .A2(n564), .ZN(n567) );
  NAND2_X1 U627 ( .A1(n565), .A2(G87), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(G288) );
  NAND2_X1 U629 ( .A1(n781), .A2(G61), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT75), .B(n568), .Z(n570) );
  NAND2_X1 U631 ( .A1(n784), .A2(G86), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U633 ( .A(KEYINPUT76), .B(n571), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n785), .A2(G73), .ZN(n572) );
  XOR2_X1 U635 ( .A(KEYINPUT2), .B(n572), .Z(n573) );
  NOR2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n780), .A2(G48), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(G305) );
  NAND2_X1 U639 ( .A1(G60), .A2(n781), .ZN(n578) );
  NAND2_X1 U640 ( .A1(G72), .A2(n785), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G85), .A2(n784), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT67), .B(n579), .ZN(n580) );
  NOR2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n780), .A2(G47), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(G290) );
  INV_X1 U647 ( .A(G1384), .ZN(n589) );
  AND2_X1 U648 ( .A1(G138), .A2(n589), .ZN(n584) );
  AND2_X1 U649 ( .A1(n880), .A2(n584), .ZN(n591) );
  NAND2_X1 U650 ( .A1(G114), .A2(n872), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G126), .A2(n873), .ZN(n585) );
  AND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G102), .A2(n878), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n753) );
  AND2_X1 U655 ( .A1(n589), .A2(n753), .ZN(n590) );
  OR2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n719) );
  INV_X1 U657 ( .A(n719), .ZN(n604) );
  OR2_X1 U658 ( .A1(n720), .A2(n604), .ZN(n629) );
  NOR2_X1 U659 ( .A1(G1966), .A2(n695), .ZN(n671) );
  NOR2_X1 U660 ( .A1(G2084), .A2(n629), .ZN(n668) );
  NOR2_X1 U661 ( .A1(n671), .A2(n668), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G8), .A2(n592), .ZN(n594) );
  NOR2_X1 U663 ( .A1(G168), .A2(n595), .ZN(n596) );
  XNOR2_X1 U664 ( .A(n596), .B(KEYINPUT97), .ZN(n600) );
  XOR2_X1 U665 ( .A(G2078), .B(KEYINPUT25), .Z(n969) );
  NOR2_X1 U666 ( .A1(n969), .A2(n629), .ZN(n598) );
  NOR2_X1 U667 ( .A1(n638), .A2(G1961), .ZN(n597) );
  NOR2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n651) );
  NAND2_X1 U669 ( .A1(n651), .A2(G301), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n600), .A2(n599), .ZN(n602) );
  XNOR2_X1 U671 ( .A(KEYINPUT31), .B(KEYINPUT98), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n602), .B(n601), .ZN(n655) );
  AND2_X1 U673 ( .A1(G40), .A2(G1996), .ZN(n603) );
  NAND2_X1 U674 ( .A1(G160), .A2(n603), .ZN(n605) );
  NOR2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U676 ( .A(n606), .B(KEYINPUT26), .Z(n608) );
  NAND2_X1 U677 ( .A1(n629), .A2(G1341), .ZN(n607) );
  NAND2_X1 U678 ( .A1(n608), .A2(n607), .ZN(n619) );
  NAND2_X1 U679 ( .A1(n784), .A2(G81), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n609), .B(KEYINPUT12), .ZN(n611) );
  NAND2_X1 U681 ( .A1(G68), .A2(n785), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U683 ( .A(KEYINPUT13), .B(n612), .ZN(n618) );
  NAND2_X1 U684 ( .A1(G43), .A2(n780), .ZN(n613) );
  XOR2_X1 U685 ( .A(KEYINPUT70), .B(n613), .Z(n616) );
  NAND2_X1 U686 ( .A1(n781), .A2(G56), .ZN(n614) );
  XOR2_X1 U687 ( .A(KEYINPUT14), .B(n614), .Z(n615) );
  NOR2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n955) );
  NOR2_X1 U690 ( .A1(n619), .A2(n955), .ZN(n633) );
  NAND2_X1 U691 ( .A1(G92), .A2(n784), .ZN(n626) );
  NAND2_X1 U692 ( .A1(G54), .A2(n780), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G66), .A2(n781), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U695 ( .A1(G79), .A2(n785), .ZN(n622) );
  XNOR2_X1 U696 ( .A(KEYINPUT71), .B(n622), .ZN(n623) );
  NOR2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n628) );
  INV_X1 U699 ( .A(KEYINPUT15), .ZN(n627) );
  NOR2_X1 U700 ( .A1(G2067), .A2(n629), .ZN(n631) );
  NOR2_X1 U701 ( .A1(n638), .A2(G1348), .ZN(n630) );
  NOR2_X1 U702 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n763), .A2(n634), .ZN(n632) );
  NAND2_X1 U704 ( .A1(n633), .A2(n632), .ZN(n636) );
  OR2_X1 U705 ( .A1(n634), .A2(n763), .ZN(n635) );
  NAND2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n637), .B(KEYINPUT94), .ZN(n643) );
  NAND2_X1 U708 ( .A1(n638), .A2(G2072), .ZN(n639) );
  XOR2_X1 U709 ( .A(KEYINPUT27), .B(n639), .Z(n641) );
  NAND2_X1 U710 ( .A1(G1956), .A2(n629), .ZN(n640) );
  NAND2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n645) );
  NOR2_X1 U712 ( .A1(G299), .A2(n645), .ZN(n642) );
  XNOR2_X1 U713 ( .A(n644), .B(KEYINPUT95), .ZN(n649) );
  XOR2_X1 U714 ( .A(KEYINPUT93), .B(KEYINPUT28), .Z(n647) );
  NAND2_X1 U715 ( .A1(n645), .A2(G299), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U718 ( .A(n650), .B(KEYINPUT29), .ZN(n653) );
  NOR2_X1 U719 ( .A1(G301), .A2(n651), .ZN(n652) );
  NAND2_X1 U720 ( .A1(n655), .A2(n654), .ZN(n669) );
  AND2_X1 U721 ( .A1(G286), .A2(G8), .ZN(n656) );
  NAND2_X1 U722 ( .A1(n669), .A2(n656), .ZN(n665) );
  INV_X1 U723 ( .A(G8), .ZN(n663) );
  NOR2_X1 U724 ( .A1(G1971), .A2(n695), .ZN(n657) );
  XNOR2_X1 U725 ( .A(n657), .B(KEYINPUT100), .ZN(n659) );
  NOR2_X1 U726 ( .A1(n629), .A2(G2090), .ZN(n658) );
  NOR2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U728 ( .A(KEYINPUT101), .B(n660), .Z(n661) );
  NAND2_X1 U729 ( .A1(n661), .A2(G303), .ZN(n662) );
  OR2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  AND2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n667) );
  NAND2_X1 U732 ( .A1(n668), .A2(G8), .ZN(n673) );
  XNOR2_X1 U733 ( .A(n669), .B(KEYINPUT99), .ZN(n670) );
  NOR2_X1 U734 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U735 ( .A1(n673), .A2(n672), .ZN(n688) );
  NAND2_X1 U736 ( .A1(G1976), .A2(G288), .ZN(n940) );
  AND2_X1 U737 ( .A1(n688), .A2(n940), .ZN(n674) );
  NAND2_X1 U738 ( .A1(n687), .A2(n674), .ZN(n679) );
  INV_X1 U739 ( .A(n940), .ZN(n677) );
  NOR2_X1 U740 ( .A1(G1976), .A2(G288), .ZN(n939) );
  NOR2_X1 U741 ( .A1(G1971), .A2(G303), .ZN(n675) );
  NOR2_X1 U742 ( .A1(n939), .A2(n675), .ZN(n676) );
  OR2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n678) );
  AND2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n695), .A2(n680), .ZN(n681) );
  NOR2_X1 U746 ( .A1(KEYINPUT33), .A2(n681), .ZN(n682) );
  XNOR2_X1 U747 ( .A(n682), .B(KEYINPUT103), .ZN(n686) );
  XOR2_X1 U748 ( .A(G1981), .B(G305), .Z(n948) );
  NAND2_X1 U749 ( .A1(n939), .A2(KEYINPUT33), .ZN(n683) );
  OR2_X1 U750 ( .A1(n683), .A2(n695), .ZN(n684) );
  AND2_X1 U751 ( .A1(n948), .A2(n684), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n699) );
  NAND2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n691) );
  NOR2_X1 U754 ( .A1(G2090), .A2(G303), .ZN(n689) );
  NAND2_X1 U755 ( .A1(G8), .A2(n689), .ZN(n690) );
  NAND2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U757 ( .A1(n695), .A2(n692), .ZN(n697) );
  NOR2_X1 U758 ( .A1(G1981), .A2(G305), .ZN(n693) );
  XOR2_X1 U759 ( .A(n693), .B(KEYINPUT24), .Z(n694) );
  OR2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n696) );
  AND2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U763 ( .A(n700), .B(KEYINPUT104), .ZN(n737) );
  NAND2_X1 U764 ( .A1(G95), .A2(n878), .ZN(n702) );
  NAND2_X1 U765 ( .A1(G131), .A2(n880), .ZN(n701) );
  NAND2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U767 ( .A(KEYINPUT90), .B(n703), .ZN(n707) );
  NAND2_X1 U768 ( .A1(G107), .A2(n872), .ZN(n705) );
  NAND2_X1 U769 ( .A1(G119), .A2(n873), .ZN(n704) );
  NAND2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n706) );
  OR2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n885) );
  AND2_X1 U772 ( .A1(n885), .A2(G1991), .ZN(n718) );
  NAND2_X1 U773 ( .A1(n873), .A2(G129), .ZN(n708) );
  XOR2_X1 U774 ( .A(KEYINPUT91), .B(n708), .Z(n710) );
  NAND2_X1 U775 ( .A1(n872), .A2(G117), .ZN(n709) );
  NAND2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U777 ( .A(KEYINPUT92), .B(n711), .ZN(n714) );
  NAND2_X1 U778 ( .A1(n878), .A2(G105), .ZN(n712) );
  XOR2_X1 U779 ( .A(KEYINPUT38), .B(n712), .Z(n713) );
  NOR2_X1 U780 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n880), .A2(G141), .ZN(n715) );
  NAND2_X1 U782 ( .A1(n716), .A2(n715), .ZN(n867) );
  AND2_X1 U783 ( .A1(n867), .A2(G1996), .ZN(n717) );
  NOR2_X1 U784 ( .A1(n718), .A2(n717), .ZN(n994) );
  NOR2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n749) );
  INV_X1 U786 ( .A(n749), .ZN(n721) );
  NOR2_X1 U787 ( .A1(n994), .A2(n721), .ZN(n741) );
  INV_X1 U788 ( .A(n741), .ZN(n732) );
  NAND2_X1 U789 ( .A1(G104), .A2(n878), .ZN(n723) );
  NAND2_X1 U790 ( .A1(G140), .A2(n880), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U792 ( .A(KEYINPUT34), .B(n724), .ZN(n729) );
  NAND2_X1 U793 ( .A1(G116), .A2(n872), .ZN(n726) );
  NAND2_X1 U794 ( .A1(G128), .A2(n873), .ZN(n725) );
  NAND2_X1 U795 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U796 ( .A(n727), .B(KEYINPUT35), .Z(n728) );
  NOR2_X1 U797 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U798 ( .A(KEYINPUT36), .B(n730), .Z(n731) );
  XNOR2_X1 U799 ( .A(KEYINPUT89), .B(n731), .ZN(n890) );
  XNOR2_X1 U800 ( .A(G2067), .B(KEYINPUT37), .ZN(n746) );
  NOR2_X1 U801 ( .A1(n890), .A2(n746), .ZN(n1010) );
  NAND2_X1 U802 ( .A1(n749), .A2(n1010), .ZN(n744) );
  NAND2_X1 U803 ( .A1(n732), .A2(n744), .ZN(n735) );
  XNOR2_X1 U804 ( .A(G1986), .B(G290), .ZN(n945) );
  NAND2_X1 U805 ( .A1(n945), .A2(n749), .ZN(n733) );
  XOR2_X1 U806 ( .A(KEYINPUT88), .B(n733), .Z(n734) );
  NOR2_X1 U807 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U808 ( .A1(n737), .A2(n736), .ZN(n751) );
  NOR2_X1 U809 ( .A1(G1996), .A2(n867), .ZN(n738) );
  XOR2_X1 U810 ( .A(KEYINPUT105), .B(n738), .Z(n1000) );
  NOR2_X1 U811 ( .A1(G1986), .A2(G290), .ZN(n739) );
  NOR2_X1 U812 ( .A1(G1991), .A2(n885), .ZN(n1007) );
  NOR2_X1 U813 ( .A1(n739), .A2(n1007), .ZN(n740) );
  NOR2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U815 ( .A1(n1000), .A2(n742), .ZN(n743) );
  XNOR2_X1 U816 ( .A(n743), .B(KEYINPUT39), .ZN(n745) );
  NAND2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n747) );
  NAND2_X1 U818 ( .A1(n890), .A2(n746), .ZN(n993) );
  NAND2_X1 U819 ( .A1(n747), .A2(n993), .ZN(n748) );
  NAND2_X1 U820 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U821 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U822 ( .A(n752), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U823 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U824 ( .A(G57), .ZN(G237) );
  AND2_X1 U825 ( .A1(G138), .A2(n880), .ZN(n754) );
  NOR2_X1 U826 ( .A1(n754), .A2(n753), .ZN(G164) );
  NAND2_X1 U827 ( .A1(G7), .A2(G661), .ZN(n755) );
  XNOR2_X1 U828 ( .A(n755), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U829 ( .A(G223), .ZN(n825) );
  NAND2_X1 U830 ( .A1(n825), .A2(G567), .ZN(n756) );
  XOR2_X1 U831 ( .A(KEYINPUT11), .B(n756), .Z(G234) );
  INV_X1 U832 ( .A(G860), .ZN(n762) );
  OR2_X1 U833 ( .A1(n955), .A2(n762), .ZN(G153) );
  NOR2_X1 U834 ( .A1(G868), .A2(n763), .ZN(n758) );
  INV_X1 U835 ( .A(G868), .ZN(n792) );
  NOR2_X1 U836 ( .A1(n792), .A2(G301), .ZN(n757) );
  NOR2_X1 U837 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U838 ( .A(KEYINPUT72), .B(n759), .ZN(G284) );
  NOR2_X1 U839 ( .A1(G868), .A2(G299), .ZN(n761) );
  NOR2_X1 U840 ( .A1(G286), .A2(n792), .ZN(n760) );
  NOR2_X1 U841 ( .A1(n761), .A2(n760), .ZN(G297) );
  NAND2_X1 U842 ( .A1(n762), .A2(G559), .ZN(n764) );
  INV_X1 U843 ( .A(n763), .ZN(n943) );
  NAND2_X1 U844 ( .A1(n764), .A2(n943), .ZN(n765) );
  XNOR2_X1 U845 ( .A(n765), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U846 ( .A1(G868), .A2(n955), .ZN(n768) );
  NAND2_X1 U847 ( .A1(G868), .A2(n943), .ZN(n766) );
  NOR2_X1 U848 ( .A1(G559), .A2(n766), .ZN(n767) );
  NOR2_X1 U849 ( .A1(n768), .A2(n767), .ZN(G282) );
  NAND2_X1 U850 ( .A1(G111), .A2(n872), .ZN(n770) );
  NAND2_X1 U851 ( .A1(G135), .A2(n880), .ZN(n769) );
  NAND2_X1 U852 ( .A1(n770), .A2(n769), .ZN(n773) );
  NAND2_X1 U853 ( .A1(n873), .A2(G123), .ZN(n771) );
  XOR2_X1 U854 ( .A(KEYINPUT18), .B(n771), .Z(n772) );
  NOR2_X1 U855 ( .A1(n773), .A2(n772), .ZN(n775) );
  NAND2_X1 U856 ( .A1(n878), .A2(G99), .ZN(n774) );
  NAND2_X1 U857 ( .A1(n775), .A2(n774), .ZN(n1008) );
  XNOR2_X1 U858 ( .A(n1008), .B(G2096), .ZN(n776) );
  XNOR2_X1 U859 ( .A(n776), .B(KEYINPUT73), .ZN(n778) );
  INV_X1 U860 ( .A(G2100), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n778), .A2(n777), .ZN(G156) );
  NAND2_X1 U862 ( .A1(n943), .A2(G559), .ZN(n801) );
  XNOR2_X1 U863 ( .A(n955), .B(n801), .ZN(n779) );
  NOR2_X1 U864 ( .A1(G860), .A2(n779), .ZN(n791) );
  NAND2_X1 U865 ( .A1(G55), .A2(n780), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G67), .A2(n781), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n789) );
  NAND2_X1 U868 ( .A1(G93), .A2(n784), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G80), .A2(n785), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U871 ( .A1(n789), .A2(n788), .ZN(n793) );
  XNOR2_X1 U872 ( .A(n793), .B(KEYINPUT74), .ZN(n790) );
  XNOR2_X1 U873 ( .A(n791), .B(n790), .ZN(G145) );
  INV_X1 U874 ( .A(G303), .ZN(G166) );
  NAND2_X1 U875 ( .A1(n792), .A2(n793), .ZN(n804) );
  XNOR2_X1 U876 ( .A(n793), .B(G288), .ZN(n794) );
  XNOR2_X1 U877 ( .A(n794), .B(G290), .ZN(n795) );
  XNOR2_X1 U878 ( .A(KEYINPUT19), .B(n795), .ZN(n797) );
  XNOR2_X1 U879 ( .A(G305), .B(KEYINPUT80), .ZN(n796) );
  XNOR2_X1 U880 ( .A(n797), .B(n796), .ZN(n798) );
  XOR2_X1 U881 ( .A(n798), .B(G299), .Z(n799) );
  XNOR2_X1 U882 ( .A(n955), .B(n799), .ZN(n800) );
  XNOR2_X1 U883 ( .A(G166), .B(n800), .ZN(n894) );
  XOR2_X1 U884 ( .A(n894), .B(n801), .Z(n802) );
  NAND2_X1 U885 ( .A1(G868), .A2(n802), .ZN(n803) );
  NAND2_X1 U886 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U887 ( .A(n805), .B(KEYINPUT81), .ZN(G295) );
  NAND2_X1 U888 ( .A1(G2078), .A2(G2084), .ZN(n806) );
  XOR2_X1 U889 ( .A(KEYINPUT20), .B(n806), .Z(n807) );
  NAND2_X1 U890 ( .A1(G2090), .A2(n807), .ZN(n809) );
  XNOR2_X1 U891 ( .A(KEYINPUT21), .B(KEYINPUT82), .ZN(n808) );
  XNOR2_X1 U892 ( .A(n809), .B(n808), .ZN(n810) );
  NAND2_X1 U893 ( .A1(n810), .A2(G2072), .ZN(n811) );
  XOR2_X1 U894 ( .A(KEYINPUT83), .B(n811), .Z(G158) );
  XNOR2_X1 U895 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U896 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n813) );
  NAND2_X1 U897 ( .A1(G132), .A2(G82), .ZN(n812) );
  XNOR2_X1 U898 ( .A(n813), .B(n812), .ZN(n814) );
  XNOR2_X1 U899 ( .A(n814), .B(KEYINPUT84), .ZN(n815) );
  NOR2_X1 U900 ( .A1(G218), .A2(n815), .ZN(n816) );
  NAND2_X1 U901 ( .A1(G96), .A2(n816), .ZN(n913) );
  NAND2_X1 U902 ( .A1(G2106), .A2(n913), .ZN(n820) );
  NAND2_X1 U903 ( .A1(G108), .A2(G120), .ZN(n817) );
  NOR2_X1 U904 ( .A1(G237), .A2(n817), .ZN(n818) );
  NAND2_X1 U905 ( .A1(G69), .A2(n818), .ZN(n914) );
  NAND2_X1 U906 ( .A1(G567), .A2(n914), .ZN(n819) );
  NAND2_X1 U907 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U908 ( .A(KEYINPUT86), .B(n821), .Z(G319) );
  INV_X1 U909 ( .A(G319), .ZN(n823) );
  NAND2_X1 U910 ( .A1(G661), .A2(G483), .ZN(n822) );
  NOR2_X1 U911 ( .A1(n823), .A2(n822), .ZN(n828) );
  NAND2_X1 U912 ( .A1(n828), .A2(G36), .ZN(n824) );
  XOR2_X1 U913 ( .A(KEYINPUT87), .B(n824), .Z(G176) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n825), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U916 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n828), .A2(n827), .ZN(G188) );
  XNOR2_X1 U919 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  XOR2_X1 U920 ( .A(G2100), .B(G2096), .Z(n830) );
  XNOR2_X1 U921 ( .A(KEYINPUT42), .B(G2678), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U923 ( .A(KEYINPUT43), .B(G2067), .Z(n832) );
  XNOR2_X1 U924 ( .A(G2090), .B(G2072), .ZN(n831) );
  XNOR2_X1 U925 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U926 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U927 ( .A(G2078), .B(G2084), .ZN(n835) );
  XNOR2_X1 U928 ( .A(n836), .B(n835), .ZN(G227) );
  XNOR2_X1 U929 ( .A(G1956), .B(KEYINPUT108), .ZN(n846) );
  XOR2_X1 U930 ( .A(G1986), .B(G1981), .Z(n838) );
  XNOR2_X1 U931 ( .A(G1961), .B(G1966), .ZN(n837) );
  XNOR2_X1 U932 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U933 ( .A(G1991), .B(G1976), .Z(n840) );
  XNOR2_X1 U934 ( .A(G1971), .B(G1996), .ZN(n839) );
  XNOR2_X1 U935 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U936 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U937 ( .A(G2474), .B(KEYINPUT41), .ZN(n843) );
  XNOR2_X1 U938 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U939 ( .A(n846), .B(n845), .ZN(G229) );
  NAND2_X1 U940 ( .A1(G112), .A2(n872), .ZN(n848) );
  NAND2_X1 U941 ( .A1(G100), .A2(n878), .ZN(n847) );
  NAND2_X1 U942 ( .A1(n848), .A2(n847), .ZN(n855) );
  NAND2_X1 U943 ( .A1(n880), .A2(G136), .ZN(n849) );
  XNOR2_X1 U944 ( .A(KEYINPUT109), .B(n849), .ZN(n852) );
  NAND2_X1 U945 ( .A1(n873), .A2(G124), .ZN(n850) );
  XOR2_X1 U946 ( .A(KEYINPUT44), .B(n850), .Z(n851) );
  NOR2_X1 U947 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U948 ( .A(KEYINPUT110), .B(n853), .Z(n854) );
  NOR2_X1 U949 ( .A1(n855), .A2(n854), .ZN(G162) );
  NAND2_X1 U950 ( .A1(G118), .A2(n872), .ZN(n857) );
  NAND2_X1 U951 ( .A1(G130), .A2(n873), .ZN(n856) );
  NAND2_X1 U952 ( .A1(n857), .A2(n856), .ZN(n864) );
  XNOR2_X1 U953 ( .A(KEYINPUT112), .B(KEYINPUT45), .ZN(n862) );
  NAND2_X1 U954 ( .A1(n878), .A2(G106), .ZN(n860) );
  NAND2_X1 U955 ( .A1(n880), .A2(G142), .ZN(n858) );
  XOR2_X1 U956 ( .A(KEYINPUT111), .B(n858), .Z(n859) );
  NAND2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U958 ( .A(n862), .B(n861), .Z(n863) );
  NOR2_X1 U959 ( .A1(n864), .A2(n863), .ZN(n889) );
  XOR2_X1 U960 ( .A(KEYINPUT48), .B(KEYINPUT116), .Z(n866) );
  XNOR2_X1 U961 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n866), .B(n865), .ZN(n868) );
  XNOR2_X1 U963 ( .A(n868), .B(n867), .ZN(n870) );
  XNOR2_X1 U964 ( .A(G160), .B(G164), .ZN(n869) );
  XNOR2_X1 U965 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U966 ( .A(n1008), .B(n871), .ZN(n887) );
  XNOR2_X1 U967 ( .A(KEYINPUT115), .B(KEYINPUT47), .ZN(n877) );
  NAND2_X1 U968 ( .A1(G115), .A2(n872), .ZN(n875) );
  NAND2_X1 U969 ( .A1(G127), .A2(n873), .ZN(n874) );
  NAND2_X1 U970 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U971 ( .A(n877), .B(n876), .ZN(n884) );
  NAND2_X1 U972 ( .A1(n878), .A2(G103), .ZN(n879) );
  XNOR2_X1 U973 ( .A(n879), .B(KEYINPUT114), .ZN(n882) );
  NAND2_X1 U974 ( .A1(G139), .A2(n880), .ZN(n881) );
  NAND2_X1 U975 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U976 ( .A1(n884), .A2(n883), .ZN(n995) );
  XOR2_X1 U977 ( .A(n885), .B(n995), .Z(n886) );
  XNOR2_X1 U978 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U979 ( .A(n889), .B(n888), .ZN(n892) );
  XNOR2_X1 U980 ( .A(n890), .B(G162), .ZN(n891) );
  XNOR2_X1 U981 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U982 ( .A1(G37), .A2(n893), .ZN(G395) );
  INV_X1 U983 ( .A(G301), .ZN(G171) );
  XOR2_X1 U984 ( .A(n894), .B(n943), .Z(n896) );
  XNOR2_X1 U985 ( .A(G286), .B(G171), .ZN(n895) );
  XNOR2_X1 U986 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U987 ( .A1(G37), .A2(n897), .ZN(G397) );
  XOR2_X1 U988 ( .A(G2438), .B(G2435), .Z(n899) );
  XNOR2_X1 U989 ( .A(G2443), .B(KEYINPUT106), .ZN(n898) );
  XNOR2_X1 U990 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U991 ( .A(n900), .B(G2454), .Z(n902) );
  XNOR2_X1 U992 ( .A(G1348), .B(G1341), .ZN(n901) );
  XNOR2_X1 U993 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U994 ( .A(G2451), .B(G2427), .Z(n904) );
  XNOR2_X1 U995 ( .A(G2430), .B(G2446), .ZN(n903) );
  XNOR2_X1 U996 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U997 ( .A(n906), .B(n905), .Z(n907) );
  NAND2_X1 U998 ( .A1(G14), .A2(n907), .ZN(n915) );
  NAND2_X1 U999 ( .A1(n915), .A2(G319), .ZN(n910) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1002 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1004 ( .A1(n912), .A2(n911), .ZN(G225) );
  XNOR2_X1 U1005 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G132), .ZN(G219) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  INV_X1 U1009 ( .A(G96), .ZN(G221) );
  INV_X1 U1010 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(G325) );
  INV_X1 U1012 ( .A(G325), .ZN(G261) );
  INV_X1 U1013 ( .A(G69), .ZN(G235) );
  INV_X1 U1014 ( .A(n915), .ZN(G401) );
  XOR2_X1 U1015 ( .A(KEYINPUT125), .B(G16), .Z(n938) );
  XNOR2_X1 U1016 ( .A(G1961), .B(G5), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(G1966), .B(G21), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(G1956), .B(G20), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(G6), .B(G1981), .ZN(n918) );
  NOR2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n925) );
  XOR2_X1 U1022 ( .A(G4), .B(KEYINPUT126), .Z(n921) );
  XNOR2_X1 U1023 ( .A(G1348), .B(KEYINPUT59), .ZN(n920) );
  XNOR2_X1 U1024 ( .A(n921), .B(n920), .ZN(n923) );
  XNOR2_X1 U1025 ( .A(G1341), .B(G19), .ZN(n922) );
  NOR2_X1 U1026 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1028 ( .A(KEYINPUT60), .B(n926), .Z(n927) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(G1971), .B(G22), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(G24), .B(G1986), .ZN(n929) );
  NOR2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n932) );
  XOR2_X1 U1033 ( .A(G1976), .B(G23), .Z(n931) );
  NAND2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(KEYINPUT58), .B(n933), .ZN(n934) );
  NOR2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1037 ( .A(KEYINPUT61), .B(n936), .Z(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n991) );
  XOR2_X1 U1039 ( .A(G16), .B(KEYINPUT56), .Z(n963) );
  XNOR2_X1 U1040 ( .A(n939), .B(KEYINPUT123), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(n942), .B(KEYINPUT124), .ZN(n961) );
  XNOR2_X1 U1043 ( .A(G1348), .B(n943), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(G1956), .B(G299), .ZN(n944) );
  NOR2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G166), .B(G1971), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(G168), .B(G1966), .ZN(n949) );
  NAND2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(n950), .B(KEYINPUT57), .ZN(n951) );
  NAND2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(G301), .B(G1961), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(n955), .B(G1341), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n988) );
  XOR2_X1 U1059 ( .A(G29), .B(KEYINPUT121), .Z(n985) );
  XOR2_X1 U1060 ( .A(G2067), .B(G26), .Z(n965) );
  XOR2_X1 U1061 ( .A(G1991), .B(G25), .Z(n964) );
  NAND2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n976) );
  XNOR2_X1 U1063 ( .A(KEYINPUT119), .B(G2072), .ZN(n966) );
  XNOR2_X1 U1064 ( .A(n966), .B(G33), .ZN(n974) );
  INV_X1 U1065 ( .A(G1996), .ZN(n967) );
  XNOR2_X1 U1066 ( .A(G32), .B(n967), .ZN(n968) );
  NAND2_X1 U1067 ( .A1(n968), .A2(G28), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(G27), .B(n969), .ZN(n970) );
  XNOR2_X1 U1069 ( .A(KEYINPUT120), .B(n970), .ZN(n971) );
  NOR2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1073 ( .A(KEYINPUT53), .B(n977), .Z(n980) );
  XOR2_X1 U1074 ( .A(KEYINPUT54), .B(G34), .Z(n978) );
  XNOR2_X1 U1075 ( .A(G2084), .B(n978), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(G35), .B(G2090), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1079 ( .A(KEYINPUT55), .B(n983), .Z(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(KEYINPUT122), .B(n986), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(G11), .A2(n989), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(n992), .B(KEYINPUT127), .ZN(n1020) );
  INV_X1 U1086 ( .A(G29), .ZN(n1018) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n1005) );
  XOR2_X1 U1088 ( .A(G2072), .B(n995), .Z(n997) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT50), .B(n998), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(G2090), .B(G162), .Z(n999) );
  NOR2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1094 ( .A(KEYINPUT51), .B(n1001), .Z(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1013) );
  XOR2_X1 U1097 ( .A(G2084), .B(G160), .Z(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT52), .B(n1014), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(n1015), .B(KEYINPUT118), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(KEYINPUT55), .A2(n1016), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1021), .ZN(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

