//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT83), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207));
  AND2_X1   g006(.A1(G211gat), .A2(G218gat), .ZN(new_n208));
  OAI22_X1  g007(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(KEYINPUT22), .ZN(new_n209));
  NOR2_X1   g008(.A1(G211gat), .A2(G218gat), .ZN(new_n210));
  NOR3_X1   g009(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT74), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(G197gat), .A2(G204gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT22), .ZN(new_n214));
  NAND2_X1  g013(.A1(G211gat), .A2(G218gat), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n213), .A2(new_n205), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G211gat), .ZN(new_n217));
  INV_X1    g016(.A(G218gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT74), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(new_n215), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n212), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(G155gat), .ZN(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G141gat), .B(G148gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n224), .B(new_n227), .C1(new_n228), .C2(KEYINPUT2), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230));
  INV_X1    g029(.A(G141gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G148gat), .ZN(new_n232));
  INV_X1    g031(.A(G148gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G141gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n227), .A2(new_n224), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n224), .A2(KEYINPUT2), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n229), .A2(new_n230), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n223), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT84), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n219), .A2(new_n242), .A3(new_n215), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT84), .B1(new_n208), .B2(new_n210), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n216), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n240), .B1(new_n216), .B2(new_n244), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n230), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n238), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT85), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n241), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n247), .A2(KEYINPUT85), .A3(new_n248), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n204), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT29), .B1(new_n212), .B2(new_n222), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n248), .B1(new_n254), .B2(KEYINPUT3), .ZN(new_n255));
  INV_X1    g054(.A(new_n202), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n240), .ZN(new_n258));
  INV_X1    g057(.A(new_n223), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT86), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n241), .A2(KEYINPUT86), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(KEYINPUT89), .B(G22gat), .C1(new_n253), .C2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G78gat), .B(G106gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT31), .B(G50gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n242), .B1(new_n219), .B2(new_n215), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT29), .B1(new_n209), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n216), .A2(new_n243), .A3(new_n244), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT3), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n248), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n250), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n259), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n252), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n203), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT86), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n255), .B(new_n256), .C1(new_n277), .C2(new_n260), .ZN(new_n278));
  NAND2_X1  g077(.A1(KEYINPUT89), .A2(G22gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n267), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT87), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(new_n253), .B2(new_n263), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n276), .A2(new_n278), .A3(KEYINPUT87), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(G22gat), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT87), .B1(new_n276), .B2(new_n278), .ZN(new_n286));
  INV_X1    g085(.A(G22gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n267), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT88), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n285), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n285), .B2(new_n288), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n281), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT90), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT90), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n294), .B(new_n281), .C1(new_n290), .C2(new_n291), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G183gat), .ZN(new_n301));
  INV_X1    g100(.A(G190gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT66), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(G183gat), .A3(G190gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT24), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G169gat), .ZN(new_n313));
  INV_X1    g112(.A(G176gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT65), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT65), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(G169gat), .B2(G176gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT23), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT25), .ZN(new_n319));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n313), .A2(new_n314), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n312), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n310), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(new_n303), .A3(new_n304), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(G169gat), .ZN(new_n328));
  OR2_X1    g127(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n321), .A2(new_n322), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n326), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n319), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n324), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n301), .A2(KEYINPUT27), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT27), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G183gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n338), .A3(new_n302), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT27), .B(G183gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(KEYINPUT28), .A3(new_n302), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT67), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT67), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n347), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT26), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n315), .A2(new_n317), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n320), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n344), .A2(new_n352), .A3(new_n306), .ZN(new_n353));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n335), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(new_n335), .B2(new_n353), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n259), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n335), .A2(new_n353), .A3(new_n354), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n344), .A2(new_n306), .A3(new_n352), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n323), .A2(new_n318), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n361), .A2(new_n312), .B1(new_n333), .B2(new_n319), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n223), .B(new_n359), .C1(new_n363), .C2(new_n356), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n358), .A2(new_n364), .A3(KEYINPUT75), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n366), .B(new_n259), .C1(new_n355), .C2(new_n357), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n300), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n367), .A3(new_n300), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(KEYINPUT30), .A3(new_n370), .ZN(new_n371));
  AOI211_X1 g170(.A(KEYINPUT30), .B(new_n300), .C1(new_n365), .C2(new_n367), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT81), .ZN(new_n376));
  XOR2_X1   g175(.A(G1gat), .B(G29gat), .Z(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n230), .B1(new_n229), .B2(new_n238), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT70), .ZN(new_n383));
  AND2_X1   g182(.A1(G113gat), .A2(G120gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(G113gat), .A2(G120gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G113gat), .ZN(new_n387));
  INV_X1    g186(.A(G120gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G113gat), .A2(G120gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(KEYINPUT70), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G134gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G127gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT68), .ZN(new_n396));
  INV_X1    g195(.A(G127gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G134gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT69), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT68), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n394), .A3(G127gat), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT69), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n397), .A3(G134gat), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n396), .A2(new_n399), .A3(new_n401), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n393), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n395), .A2(new_n398), .A3(new_n392), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n390), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n382), .A2(new_n239), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n408), .B1(new_n393), .B2(new_n404), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n412), .B1(new_n272), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n405), .A2(new_n229), .A3(new_n238), .A4(new_n409), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n415), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n420));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n416), .A2(new_n418), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n272), .A2(new_n413), .A3(new_n412), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(KEYINPUT77), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n421), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n229), .A2(new_n230), .A3(new_n238), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n381), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n429), .B2(new_n410), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT77), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n431), .A3(new_n418), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n248), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n416), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n420), .B1(new_n435), .B2(new_n427), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n433), .A2(KEYINPUT79), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT79), .B1(new_n433), .B2(new_n436), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n380), .B(new_n423), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n424), .A2(KEYINPUT77), .A3(new_n425), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n432), .A2(new_n421), .A3(new_n411), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n436), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n433), .A2(KEYINPUT79), .A3(new_n436), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n380), .B1(new_n448), .B2(new_n423), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n441), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n446), .A2(new_n447), .B1(new_n419), .B2(new_n422), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n451), .A2(new_n440), .A3(new_n380), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n374), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT82), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT6), .B1(new_n451), .B2(new_n380), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n448), .A2(new_n423), .ZN(new_n456));
  INV_X1    g255(.A(new_n380), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n449), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n374), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT71), .B1(new_n360), .B2(new_n362), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT71), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n335), .A2(new_n465), .A3(new_n353), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n410), .A3(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(KEYINPUT71), .B(new_n413), .C1(new_n360), .C2(new_n362), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(G227gat), .ZN(new_n470));
  INV_X1    g269(.A(G233gat), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT34), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n470), .A2(new_n471), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n467), .A2(new_n474), .A3(new_n468), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT32), .ZN(new_n476));
  XNOR2_X1  g275(.A(G15gat), .B(G43gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(G71gat), .B(G99gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT33), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n475), .A2(new_n480), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT72), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT72), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n475), .A2(new_n485), .A3(new_n480), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n479), .B1(new_n475), .B2(KEYINPUT32), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n482), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT73), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n473), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT34), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n472), .B(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n479), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n484), .B2(new_n486), .ZN(new_n496));
  OAI211_X1 g295(.A(KEYINPUT73), .B(new_n493), .C1(new_n496), .C2(new_n482), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n296), .A2(new_n454), .A3(new_n463), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n370), .A2(KEYINPUT30), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(new_n368), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n503), .B2(new_n372), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n371), .A2(KEYINPUT91), .A3(new_n373), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n450), .A2(new_n452), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n473), .B1(new_n496), .B2(new_n482), .ZN(new_n509));
  INV_X1    g308(.A(new_n486), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n485), .B1(new_n475), .B2(new_n480), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n488), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n482), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n493), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  NOR4_X1   g314(.A1(new_n507), .A2(new_n508), .A3(new_n515), .A4(KEYINPUT35), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n296), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT36), .B1(new_n509), .B2(new_n514), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n498), .B2(KEYINPUT36), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n434), .A2(new_n416), .A3(new_n421), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT39), .ZN(new_n521));
  INV_X1    g320(.A(new_n416), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n411), .A2(new_n414), .B1(new_n522), .B2(new_n417), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n521), .B1(new_n427), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT92), .B(KEYINPUT39), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n427), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n525), .A2(KEYINPUT40), .A3(new_n380), .A4(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT40), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n380), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(new_n524), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n449), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n504), .A2(new_n533), .A3(new_n505), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT93), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT93), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n504), .A2(new_n533), .A3(new_n505), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n300), .A2(KEYINPUT37), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n370), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n358), .A2(new_n364), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT38), .B1(new_n541), .B2(KEYINPUT37), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT38), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n365), .A2(KEYINPUT37), .A3(new_n367), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n543), .A2(new_n546), .A3(new_n368), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n293), .A2(new_n295), .B1(new_n508), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n519), .B1(new_n538), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n454), .A2(new_n463), .ZN(new_n550));
  INV_X1    g349(.A(new_n296), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n500), .A2(new_n517), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g356(.A1(KEYINPUT94), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(G71gat), .B2(G78gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n557), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT21), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G127gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G15gat), .B(G22gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT16), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n568), .B2(G1gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(G1gat), .B2(new_n567), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G8gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n562), .B2(new_n561), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n566), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(new_n225), .ZN(new_n576));
  XOR2_X1   g375(.A(G183gat), .B(G211gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n574), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT95), .Z(new_n581));
  INV_X1    g380(.A(KEYINPUT41), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT96), .ZN(new_n584));
  XOR2_X1   g383(.A(G190gat), .B(G218gat), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT100), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT101), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n584), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590));
  INV_X1    g389(.A(G36gat), .ZN(new_n591));
  AND2_X1   g390(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G29gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n597), .A2(KEYINPUT15), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(KEYINPUT15), .ZN(new_n599));
  XNOR2_X1  g398(.A(G43gat), .B(G50gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G99gat), .A2(G106gat), .ZN(new_n605));
  INV_X1    g404(.A(G85gat), .ZN(new_n606));
  INV_X1    g405(.A(G92gat), .ZN(new_n607));
  AOI22_X1  g406(.A1(KEYINPUT8), .A2(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT7), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G99gat), .B(G106gat), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n614), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n610), .A2(new_n616), .A3(new_n612), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OAI22_X1  g417(.A1(new_n604), .A2(new_n618), .B1(new_n582), .B2(new_n581), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n603), .A2(KEYINPUT17), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n621), .B1(new_n601), .B2(new_n602), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n618), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT99), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n625), .B(new_n618), .C1(new_n620), .C2(new_n622), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n619), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n586), .A2(KEYINPUT101), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n590), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n627), .A2(new_n628), .A3(new_n590), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n589), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(new_n588), .A3(new_n629), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n572), .B1(new_n620), .B2(new_n622), .ZN(new_n637));
  NAND2_X1  g436(.A1(G229gat), .A2(G233gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n603), .A2(new_n571), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT18), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n603), .B(new_n571), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n638), .B(KEYINPUT13), .Z(new_n644));
  AOI22_X1  g443(.A1(new_n640), .A2(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G113gat), .B(G141gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G197gat), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT11), .B(G169gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT12), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n642), .A2(new_n645), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n642), .B2(new_n645), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(G230gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(new_n471), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n615), .A2(new_n560), .A3(new_n617), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n560), .B1(new_n615), .B2(new_n617), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n618), .A2(new_n561), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT10), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n662), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n663), .A2(KEYINPUT10), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n661), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n659), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n665), .B(KEYINPUT102), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  INV_X1    g474(.A(new_n661), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n658), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n673), .A2(KEYINPUT103), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR4_X1   g482(.A1(new_n579), .A2(new_n636), .A3(new_n655), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n554), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n508), .A2(KEYINPUT104), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n461), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g492(.A1(new_n554), .A2(new_n507), .A3(new_n684), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n694), .B2(G8gat), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n698), .B(KEYINPUT105), .C1(new_n701), .C2(new_n697), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n699), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n699), .B2(new_n702), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(G1325gat));
  OR3_X1    g505(.A1(new_n685), .A2(G15gat), .A3(new_n515), .ZN(new_n707));
  INV_X1    g506(.A(new_n519), .ZN(new_n708));
  OAI21_X1  g507(.A(G15gat), .B1(new_n685), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(G1326gat));
  NOR2_X1   g509(.A1(new_n685), .A2(new_n296), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT43), .B(G22gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  NOR2_X1   g512(.A1(new_n553), .A2(new_n635), .ZN(new_n714));
  INV_X1    g513(.A(new_n579), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(new_n655), .A3(new_n683), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n595), .A3(new_n691), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT45), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n553), .B2(new_n635), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n538), .A2(new_n548), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n552), .A2(new_n723), .A3(new_n708), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n499), .A2(KEYINPUT35), .B1(new_n516), .B2(new_n296), .ZN(new_n725));
  OAI211_X1 g524(.A(KEYINPUT44), .B(new_n636), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n716), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n728), .B2(new_n690), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n720), .A2(new_n729), .ZN(G1328gat));
  NOR3_X1   g529(.A1(new_n717), .A2(G36gat), .A3(new_n506), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT46), .ZN(new_n732));
  OAI21_X1  g531(.A(G36gat), .B1(new_n728), .B2(new_n506), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1329gat));
  NAND4_X1  g533(.A1(new_n722), .A2(new_n519), .A3(new_n726), .A4(new_n716), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G43gat), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n515), .A2(G43gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n718), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(new_n738), .A3(KEYINPUT47), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n736), .A2(KEYINPUT107), .B1(new_n718), .B2(new_n737), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n735), .A2(new_n742), .A3(G43gat), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n740), .B(KEYINPUT47), .C1(new_n741), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n736), .A2(KEYINPUT107), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(new_n743), .A3(new_n738), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT108), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n739), .B1(new_n744), .B2(new_n748), .ZN(G1330gat));
  NOR3_X1   g548(.A1(new_n717), .A2(G50gat), .A3(new_n296), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT48), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(KEYINPUT109), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G50gat), .B1(new_n728), .B2(new_n296), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n751), .A2(KEYINPUT109), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1331gat));
  INV_X1    g555(.A(new_n683), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n653), .A2(new_n654), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n579), .A2(new_n636), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n690), .B(KEYINPUT110), .Z(new_n760));
  NAND3_X1  g559(.A1(new_n554), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g561(.A1(new_n554), .A2(new_n759), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n507), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT49), .B(G64gat), .Z(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(G1333gat));
  NAND3_X1  g568(.A1(new_n765), .A2(G71gat), .A3(new_n519), .ZN(new_n770));
  INV_X1    g569(.A(G71gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n763), .B2(new_n515), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n765), .A2(new_n551), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g575(.A1(new_n715), .A2(new_n758), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n714), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n780), .A2(new_n606), .A3(new_n683), .A4(new_n691), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n715), .A2(new_n758), .A3(new_n757), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n727), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783), .B2(new_n690), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT112), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n781), .A2(new_n787), .A3(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(G1336gat));
  NAND3_X1  g588(.A1(new_n727), .A2(new_n507), .A3(new_n782), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(G92gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n779), .A2(KEYINPUT113), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n778), .B(new_n792), .Z(new_n793));
  NOR3_X1   g592(.A1(new_n757), .A2(G92gat), .A3(new_n506), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n794), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n796), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n795), .A2(new_n796), .B1(new_n798), .B2(new_n791), .ZN(G1337gat));
  INV_X1    g598(.A(new_n515), .ZN(new_n800));
  XNOR2_X1  g599(.A(KEYINPUT114), .B(G99gat), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n780), .A2(new_n800), .A3(new_n683), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n783), .A2(new_n708), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n803), .B2(new_n801), .ZN(G1338gat));
  NAND3_X1  g603(.A1(new_n727), .A2(new_n551), .A3(new_n782), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n805), .A2(G106gat), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n296), .A2(new_n757), .A3(G106gat), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n793), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n780), .A2(new_n807), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n809), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n808), .A2(new_n809), .B1(new_n811), .B2(new_n806), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n670), .A2(new_n671), .A3(new_n661), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n677), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n658), .B1(new_n672), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n678), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n820), .A2(KEYINPUT115), .A3(new_n678), .A4(new_n821), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n638), .B1(new_n637), .B2(new_n639), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n643), .A2(new_n644), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n649), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n652), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n632), .A2(new_n634), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n813), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n832), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n834), .A2(KEYINPUT116), .A3(new_n824), .A4(new_n825), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n683), .A2(new_n831), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n826), .B2(new_n655), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n635), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n715), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NOR4_X1   g639(.A1(new_n579), .A2(new_n636), .A3(new_n758), .A4(new_n683), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(new_n760), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n296), .A2(new_n498), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n843), .A2(new_n506), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n758), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n842), .A2(new_n296), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n690), .A2(new_n507), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n800), .A3(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n850), .A2(new_n387), .A3(new_n655), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n847), .A2(new_n851), .ZN(G1340gat));
  AOI21_X1  g651(.A(G120gat), .B1(new_n846), .B2(new_n683), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n850), .A2(new_n388), .A3(new_n757), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(G1341gat));
  NAND3_X1  g654(.A1(new_n846), .A2(new_n397), .A3(new_n715), .ZN(new_n856));
  OAI21_X1  g655(.A(G127gat), .B1(new_n850), .B2(new_n579), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1342gat));
  NOR2_X1   g657(.A1(new_n635), .A2(new_n507), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n394), .A3(new_n845), .A4(new_n859), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n850), .B2(new_n635), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G1343gat));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n842), .A2(new_n865), .A3(new_n551), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n708), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT117), .Z(new_n868));
  NAND4_X1  g667(.A1(new_n715), .A2(new_n655), .A3(new_n635), .A4(new_n757), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n821), .A2(new_n678), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT55), .B1(new_n815), .B2(new_n817), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT118), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n820), .A2(new_n873), .A3(new_n678), .A4(new_n821), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n758), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n636), .B1(new_n837), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n876), .B1(new_n833), .B2(new_n835), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n869), .B1(new_n877), .B2(new_n715), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(new_n551), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n866), .B(new_n868), .C1(new_n865), .C2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G141gat), .B1(new_n880), .B2(new_n655), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n519), .A2(new_n296), .ZN(new_n882));
  AND4_X1   g681(.A1(new_n506), .A2(new_n842), .A3(new_n760), .A4(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n655), .A2(G141gat), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n883), .A2(new_n884), .B1(new_n885), .B2(KEYINPUT58), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n885), .A2(KEYINPUT58), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n881), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n881), .B2(new_n886), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n233), .A2(KEYINPUT59), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n891), .B1(new_n880), .B2(new_n757), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n655), .B1(new_n822), .B2(KEYINPUT118), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n895), .A2(new_n874), .B1(new_n683), .B2(new_n831), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n896), .A2(new_n636), .B1(new_n832), .B2(new_n822), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n841), .B1(new_n897), .B2(new_n579), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n894), .B(new_n865), .C1(new_n898), .C2(new_n296), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n832), .A2(new_n822), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n579), .B1(new_n876), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n296), .B1(new_n901), .B2(new_n869), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT121), .B1(new_n902), .B2(KEYINPUT57), .ZN(new_n903));
  OAI211_X1 g702(.A(KEYINPUT57), .B(new_n551), .C1(new_n840), .C2(new_n841), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n899), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n868), .A2(new_n683), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G148gat), .ZN(new_n908));
  XOR2_X1   g707(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n893), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  AOI211_X1 g710(.A(KEYINPUT122), .B(new_n909), .C1(new_n907), .C2(G148gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n892), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n883), .A2(new_n233), .A3(new_n683), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1345gat));
  OAI21_X1  g714(.A(G155gat), .B1(new_n880), .B2(new_n579), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n883), .A2(new_n225), .A3(new_n715), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1346gat));
  NAND4_X1  g717(.A1(new_n843), .A2(new_n226), .A3(new_n859), .A4(new_n882), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n880), .B2(new_n635), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G162gat), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n880), .A2(new_n920), .A3(new_n635), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(G1347gat));
  NOR3_X1   g723(.A1(new_n760), .A2(new_n506), .A3(new_n515), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n848), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n926), .A2(new_n313), .A3(new_n655), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n842), .A2(new_n507), .A3(new_n845), .A4(new_n690), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n758), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n927), .A2(new_n930), .ZN(G1348gat));
  AOI21_X1  g730(.A(G176gat), .B1(new_n929), .B2(new_n683), .ZN(new_n932));
  INV_X1    g731(.A(new_n926), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n757), .B1(new_n329), .B2(new_n330), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(G1349gat));
  OAI21_X1  g734(.A(G183gat), .B1(new_n926), .B2(new_n579), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n929), .A2(new_n342), .A3(new_n715), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT60), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n929), .A2(new_n302), .A3(new_n636), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n933), .A2(new_n636), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(G190gat), .ZN(new_n946));
  AOI211_X1 g745(.A(KEYINPUT61), .B(new_n302), .C1(new_n933), .C2(new_n636), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1351gat));
  AND2_X1   g747(.A1(new_n842), .A2(new_n690), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n882), .A2(new_n507), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT124), .Z(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  XNOR2_X1  g752(.A(KEYINPUT125), .B(G197gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n758), .A3(new_n954), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n760), .A2(new_n506), .A3(new_n519), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n905), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n957), .A2(new_n655), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n958), .B2(new_n954), .ZN(G1352gat));
  INV_X1    g758(.A(new_n957), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(KEYINPUT126), .A3(new_n683), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n962), .B1(new_n957), .B2(new_n757), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n961), .A2(G204gat), .A3(new_n963), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n757), .A2(G204gat), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT62), .B1(new_n952), .B2(new_n965), .ZN(new_n966));
  OR3_X1    g765(.A1(new_n952), .A2(KEYINPUT62), .A3(new_n965), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n217), .A3(new_n715), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n960), .A2(new_n715), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n970), .B2(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  NAND3_X1  g772(.A1(new_n953), .A2(new_n218), .A3(new_n636), .ZN(new_n974));
  OAI21_X1  g773(.A(G218gat), .B1(new_n957), .B2(new_n635), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT127), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n974), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1355gat));
endmodule


