//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1383,
    new_n1384, new_n1385;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  AND2_X1   g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n225), .A2(G20), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n212), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0029(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G226), .B(G232), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n214), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G58), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G169), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(new_n226), .A3(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT67), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n206), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n251), .A2(new_n254), .A3(G274), .A4(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n251), .A2(G238), .A3(new_n252), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n216), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G226), .A2(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(G232), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n258), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n259), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n226), .A2(new_n247), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n256), .B(new_n257), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT13), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n261), .A2(G1698), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G226), .B2(G1698), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI22_X1  g0075(.A1(new_n272), .A2(new_n275), .B1(new_n258), .B2(new_n216), .ZN(new_n276));
  INV_X1    g0076(.A(new_n268), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT13), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n278), .A2(new_n279), .A3(new_n256), .A4(new_n257), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n246), .B1(new_n270), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT14), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n270), .A2(new_n280), .ZN(new_n283));
  INV_X1    g0083(.A(G179), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n281), .A2(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n281), .A2(KEYINPUT72), .A3(new_n282), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT72), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n283), .A2(G169), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n288), .B1(new_n289), .B2(KEYINPUT14), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n286), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G1), .A2(G13), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT69), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(new_n207), .A3(new_n258), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT69), .B1(G20), .B2(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G50), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n207), .A2(G33), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G68), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n302), .A2(G77), .B1(G20), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n295), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT11), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(G68), .ZN(new_n308));
  XOR2_X1   g0108(.A(new_n308), .B(KEYINPUT12), .Z(new_n309));
  AOI21_X1  g0109(.A(new_n294), .B1(new_n206), .B2(G20), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n306), .B(new_n309), .C1(new_n303), .C2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n305), .A2(KEYINPUT11), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n291), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n283), .A2(G200), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n314), .B(new_n317), .C1(new_n318), .C2(new_n283), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n320), .A2(KEYINPUT73), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(KEYINPUT73), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n251), .A2(G226), .A3(new_n252), .ZN(new_n323));
  INV_X1    g0123(.A(G1698), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G222), .ZN(new_n325));
  NAND2_X1  g0125(.A1(G223), .A2(G1698), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n266), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n327), .B(new_n277), .C1(G77), .C2(new_n266), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n323), .A2(new_n328), .A3(new_n256), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(new_n318), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(G200), .B2(new_n329), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT8), .B(G58), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n333), .A2(new_n302), .B1(new_n299), .B2(G150), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT70), .B1(new_n203), .B2(G20), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT70), .ZN(new_n336));
  AOI211_X1 g0136(.A(new_n336), .B(new_n207), .C1(new_n201), .C2(new_n202), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n334), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n294), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT9), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n307), .A2(G50), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(new_n310), .B2(G50), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n340), .B1(new_n339), .B2(new_n342), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n331), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT10), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT17), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n333), .A2(new_n307), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n310), .B2(new_n333), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n299), .A2(G159), .ZN(new_n351));
  INV_X1    g0151(.A(G58), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n303), .ZN(new_n353));
  OAI21_X1  g0153(.A(G20), .B1(new_n353), .B2(new_n202), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  NOR4_X1   g0156(.A1(new_n273), .A2(new_n274), .A3(new_n356), .A4(G20), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT74), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n303), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n264), .A2(new_n207), .A3(new_n265), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n356), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n265), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(KEYINPUT74), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n355), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n295), .B1(new_n364), .B2(KEYINPUT16), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n303), .B1(new_n361), .B2(new_n362), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(new_n355), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n350), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(G223), .A2(G1698), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n215), .B2(G1698), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n266), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT75), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT75), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(G33), .A3(G87), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n277), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n251), .A2(G232), .A3(new_n252), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n380), .A2(new_n318), .A3(new_n256), .A4(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n377), .B1(new_n266), .B2(new_n371), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n256), .B(new_n381), .C1(new_n383), .C2(new_n268), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n347), .B1(new_n369), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n355), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n361), .A2(KEYINPUT74), .A3(new_n362), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n362), .B2(KEYINPUT74), .ZN(new_n391));
  OAI211_X1 g0191(.A(KEYINPUT16), .B(new_n389), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(new_n294), .A3(new_n368), .ZN(new_n393));
  AND4_X1   g0193(.A1(new_n347), .A2(new_n393), .A3(new_n349), .A4(new_n387), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n380), .A2(G179), .A3(new_n256), .A4(new_n381), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n384), .A2(G169), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT18), .B1(new_n369), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n393), .A2(new_n349), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n396), .A2(new_n397), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n339), .A2(new_n342), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n329), .A2(new_n246), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n406), .B(new_n407), .C1(G179), .C2(new_n329), .ZN(new_n408));
  INV_X1    g0208(.A(new_n307), .ZN(new_n409));
  INV_X1    g0209(.A(G77), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n311), .B2(new_n410), .ZN(new_n412));
  XOR2_X1   g0212(.A(KEYINPUT15), .B(G87), .Z(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n302), .B1(G20), .B2(G77), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n333), .A2(new_n299), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n295), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G107), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n268), .B1(new_n275), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G238), .A2(G1698), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n261), .B2(G1698), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n275), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n251), .A2(G244), .A3(new_n252), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n256), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT71), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT71), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n422), .A2(new_n426), .A3(new_n256), .A4(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n417), .B1(new_n428), .B2(new_n385), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n318), .B1(new_n425), .B2(new_n427), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n425), .A2(new_n427), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n417), .B1(new_n432), .B2(new_n246), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n428), .A2(new_n284), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n346), .A2(new_n405), .A3(new_n408), .A4(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n321), .A2(new_n322), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT4), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(G1698), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(G244), .C1(new_n274), .C2(new_n273), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G283), .ZN(new_n443));
  INV_X1    g0243(.A(G244), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n264), .B2(new_n265), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n442), .B(new_n443), .C1(new_n445), .C2(KEYINPUT4), .ZN(new_n446));
  OAI21_X1  g0246(.A(G250), .B1(new_n273), .B2(new_n274), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n324), .B1(new_n447), .B2(KEYINPUT4), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n277), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n206), .A2(G45), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT5), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(G41), .ZN(new_n452));
  INV_X1    g0252(.A(G41), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT5), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n452), .A2(new_n251), .A3(G274), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(G41), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n454), .A2(new_n456), .A3(new_n206), .A4(G45), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(new_n251), .A3(G257), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n449), .A2(new_n459), .A3(G190), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n449), .A2(new_n459), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n460), .A2(KEYINPUT79), .B1(new_n461), .B2(G200), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT78), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n361), .A2(new_n362), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G107), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT6), .ZN(new_n466));
  AND2_X1   g0266(.A1(G97), .A2(G107), .ZN(new_n467));
  NOR2_X1   g0267(.A1(G97), .A2(G107), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT76), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT6), .A2(G97), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(G107), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n418), .A2(KEYINPUT76), .A3(KEYINPUT6), .A4(G97), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n474), .A2(G20), .B1(G77), .B2(new_n299), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n295), .B1(new_n465), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n206), .A2(G33), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n307), .A2(new_n477), .A3(new_n293), .A4(new_n292), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n307), .A2(new_n216), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n479), .A2(KEYINPUT77), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT77), .B1(new_n479), .B2(new_n480), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n463), .B1(new_n476), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n474), .A2(G20), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n299), .A2(G77), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n418), .B1(new_n361), .B2(new_n362), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n294), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n479), .A2(new_n480), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT77), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n479), .A2(KEYINPUT77), .A3(new_n480), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n489), .A2(KEYINPUT78), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT79), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n449), .A2(new_n459), .A3(new_n496), .A4(G190), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n462), .A2(new_n484), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n266), .A2(new_n207), .A3(G68), .ZN(new_n499));
  INV_X1    g0299(.A(G87), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(new_n216), .A3(new_n418), .ZN(new_n501));
  OAI211_X1 g0301(.A(KEYINPUT19), .B(new_n501), .C1(new_n259), .C2(G20), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n301), .A2(new_n216), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n499), .B(new_n502), .C1(KEYINPUT19), .C2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n413), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n504), .A2(new_n294), .B1(new_n409), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n478), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G87), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G45), .ZN(new_n510));
  OAI211_X1 g0310(.A(KEYINPUT80), .B(G250), .C1(new_n510), .C2(G1), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT80), .ZN(new_n512));
  AOI21_X1  g0312(.A(G274), .B1(new_n512), .B2(G250), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n511), .B1(new_n513), .B2(new_n450), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n251), .ZN(new_n515));
  INV_X1    g0315(.A(G116), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n258), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G238), .A2(G1698), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(new_n444), .B2(G1698), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n517), .B1(new_n519), .B2(new_n266), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n515), .B1(new_n520), .B2(new_n268), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G200), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n515), .B(G190), .C1(new_n520), .C2(new_n268), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(G169), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n284), .B2(new_n521), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n507), .A2(new_n413), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n506), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n509), .A2(new_n524), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n449), .A2(new_n459), .A3(G179), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n246), .B1(new_n449), .B2(new_n459), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n531), .A2(new_n532), .B1(new_n476), .B2(new_n483), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n207), .B2(G107), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n418), .A2(KEYINPUT23), .A3(G20), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n535), .A2(new_n536), .B1(new_n517), .B2(new_n207), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n207), .B(G87), .C1(new_n273), .C2(new_n274), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n538), .A2(KEYINPUT22), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n538), .A2(KEYINPUT22), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(KEYINPUT24), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT24), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n538), .B(KEYINPUT22), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(new_n537), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n294), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n409), .A2(new_n418), .ZN(new_n547));
  OR2_X1    g0347(.A1(new_n547), .A2(KEYINPUT25), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(KEYINPUT25), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n548), .B(new_n549), .C1(new_n418), .C2(new_n478), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n266), .A2(G257), .A3(G1698), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n266), .A2(G250), .A3(new_n324), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G294), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n277), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n457), .A2(new_n251), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G264), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n455), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G200), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n556), .A2(G190), .A3(new_n455), .A4(new_n558), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n546), .A2(new_n551), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n498), .A2(new_n529), .A3(new_n533), .A4(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n443), .B(new_n207), .C1(G33), .C2(new_n216), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n516), .A2(G20), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n294), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n566), .B(KEYINPUT20), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n409), .A2(new_n516), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n478), .B2(new_n516), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n557), .A2(G270), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n455), .ZN(new_n572));
  AND2_X1   g0372(.A1(G264), .A2(G1698), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n273), .B2(new_n274), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n264), .A2(G303), .A3(new_n265), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT81), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n217), .B1(new_n264), .B2(new_n265), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(new_n324), .ZN(new_n580));
  OAI211_X1 g0380(.A(G257), .B(new_n324), .C1(new_n273), .C2(new_n274), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n581), .A2(KEYINPUT81), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n577), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(KEYINPUT82), .A3(new_n277), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT82), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(KEYINPUT81), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n266), .A2(new_n578), .A3(G257), .A4(new_n324), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n576), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n585), .B1(new_n588), .B2(new_n268), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n572), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n570), .B1(new_n590), .B2(new_n385), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT83), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(KEYINPUT83), .B(new_n570), .C1(new_n590), .C2(new_n385), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n590), .A2(G190), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n572), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT82), .B1(new_n583), .B2(new_n277), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n588), .A2(new_n585), .A3(new_n268), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  OAI21_X1  g0401(.A(G169), .B1(new_n567), .B2(new_n569), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT21), .B1(new_n590), .B2(new_n602), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n570), .A2(new_n284), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n604), .A2(new_n605), .B1(new_n590), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n596), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n559), .A2(new_n246), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n556), .A2(new_n284), .A3(new_n455), .A4(new_n558), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n541), .A2(KEYINPUT24), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n544), .A2(new_n543), .A3(new_n537), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n295), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n609), .B(new_n610), .C1(new_n613), .C2(new_n550), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NOR4_X1   g0415(.A1(new_n439), .A2(new_n563), .A3(new_n608), .A4(new_n615), .ZN(G372));
  AOI21_X1  g0416(.A(new_n563), .B1(new_n607), .B2(new_n614), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n526), .A2(new_n528), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n506), .A2(new_n522), .A3(new_n508), .A4(new_n523), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT26), .B1(new_n620), .B2(new_n533), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n484), .A2(new_n495), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  INV_X1    g0423(.A(new_n532), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n530), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n529), .A2(new_n622), .A3(new_n623), .A4(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n621), .A2(new_n626), .A3(new_n618), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n438), .B1(new_n617), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n408), .ZN(new_n629));
  AOI221_X4 g0429(.A(KEYINPUT18), .B1(new_n397), .B2(new_n396), .C1(new_n393), .C2(new_n349), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n401), .B1(new_n400), .B2(new_n402), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n316), .ZN(new_n633));
  INV_X1    g0433(.A(new_n435), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n633), .B1(new_n319), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n632), .B1(new_n635), .B2(new_n395), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n629), .B1(new_n636), .B2(new_n346), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n628), .A2(new_n637), .ZN(G369));
  NAND3_X1  g0438(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G213), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n596), .B(new_n607), .C1(new_n570), .C2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n590), .A2(new_n606), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n601), .B1(new_n600), .B2(new_n603), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n590), .A2(KEYINPUT21), .A3(new_n602), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n570), .A2(new_n645), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n644), .B1(new_n613), .B2(new_n550), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n614), .A2(new_n562), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n546), .A2(new_n551), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n656), .A2(new_n609), .A3(new_n610), .A4(new_n644), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n653), .A2(G330), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n655), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT84), .B1(new_n607), .B2(new_n644), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT84), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n650), .A2(new_n662), .A3(new_n645), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n660), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g0464(.A(new_n644), .B(KEYINPUT85), .Z(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n614), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n659), .A2(new_n668), .ZN(G399));
  INV_X1    g0469(.A(new_n210), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G41), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n501), .A2(G116), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G1), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n225), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n672), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT89), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n498), .A2(new_n533), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n647), .B(new_n614), .C1(new_n648), .C2(new_n649), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n562), .A2(new_n619), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n678), .B1(new_n683), .B2(new_n618), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n618), .A2(new_n678), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n624), .A2(new_n530), .B1(new_n489), .B2(new_n494), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT26), .B1(new_n686), .B2(new_n529), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n687), .A2(KEYINPUT90), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n529), .A2(new_n622), .A3(KEYINPUT26), .A4(new_n625), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n687), .B2(KEYINPUT90), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n685), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OAI211_X1 g0491(.A(KEYINPUT29), .B(new_n645), .C1(new_n684), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n460), .A2(KEYINPUT79), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n461), .A2(G200), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n497), .A3(new_n694), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n529), .B(new_n533), .C1(new_n695), .C2(new_n622), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(new_n681), .A3(new_n562), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n621), .A2(new_n626), .A3(new_n618), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n666), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n692), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n614), .A2(new_n562), .A3(new_n665), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n697), .A2(new_n596), .A3(new_n607), .A4(new_n703), .ZN(new_n704));
  XOR2_X1   g0504(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n461), .A2(new_n559), .A3(KEYINPUT88), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT88), .B1(new_n461), .B2(new_n559), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n444), .A2(G1698), .ZN(new_n710));
  OAI221_X1 g0510(.A(new_n710), .B1(G238), .B2(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n711));
  INV_X1    g0511(.A(new_n517), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n713), .A2(new_n277), .B1(new_n251), .B2(new_n514), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G179), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n600), .A2(KEYINPUT87), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT87), .ZN(new_n717));
  INV_X1    g0517(.A(new_n715), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n590), .B2(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n709), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n714), .A2(new_n556), .A3(G179), .A4(new_n558), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n461), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n590), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(KEYINPUT30), .A3(new_n590), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n666), .B(new_n706), .C1(new_n720), .C2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n726), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT30), .B1(new_n722), .B2(new_n590), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n709), .A2(new_n716), .A3(new_n719), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n645), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n704), .B(new_n728), .C1(KEYINPUT31), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n702), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n677), .B1(new_n737), .B2(G1), .ZN(G364));
  NOR2_X1   g0538(.A1(new_n653), .A2(G330), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT91), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n653), .A2(G330), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n207), .A2(G13), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G45), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n672), .A2(G1), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n293), .B1(G20), .B2(new_n246), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT92), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n670), .A2(new_n266), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n225), .A2(new_n510), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n752), .B(new_n753), .C1(new_n241), .C2(new_n510), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n670), .A2(new_n275), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n755), .A2(G355), .B1(new_n516), .B2(new_n670), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n751), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n749), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n284), .A2(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n207), .A2(G190), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n385), .A2(G179), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n762), .A2(new_n410), .B1(new_n418), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n207), .A2(new_n318), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n766), .A2(new_n759), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(G58), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n760), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT32), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n207), .A2(new_n284), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G190), .A3(G200), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n774), .A2(new_n318), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G50), .A2(new_n776), .B1(new_n778), .B2(G68), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n766), .A2(new_n763), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n500), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n207), .B1(new_n769), .B2(G190), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n275), .B(new_n781), .C1(G97), .C2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n768), .A2(new_n773), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G326), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n775), .A2(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n266), .B(new_n787), .C1(G322), .C2(new_n767), .ZN(new_n788));
  INV_X1    g0588(.A(new_n764), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G283), .A2(new_n789), .B1(new_n761), .B2(G311), .ZN(new_n790));
  INV_X1    g0590(.A(new_n780), .ZN(new_n791));
  INV_X1    g0591(.A(new_n770), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G303), .A2(new_n791), .B1(new_n792), .B2(G329), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT33), .B(G317), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n778), .A2(new_n794), .B1(new_n783), .B2(G294), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n788), .A2(new_n790), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n758), .B1(new_n785), .B2(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n757), .A2(new_n797), .A3(new_n744), .ZN(new_n798));
  INV_X1    g0598(.A(new_n748), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n653), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n745), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  INV_X1    g0602(.A(new_n744), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n429), .A2(new_n430), .B1(new_n417), .B2(new_n645), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n435), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n433), .A2(new_n434), .A3(new_n645), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n747), .ZN(new_n808));
  INV_X1    g0608(.A(new_n767), .ZN(new_n809));
  INV_X1    g0609(.A(G294), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n809), .A2(new_n810), .B1(new_n762), .B2(new_n516), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n275), .B1(new_n782), .B2(new_n216), .C1(new_n418), .C2(new_n780), .ZN(new_n812));
  INV_X1    g0612(.A(G283), .ZN(new_n813));
  INV_X1    g0613(.A(G303), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n777), .A2(new_n813), .B1(new_n775), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n764), .A2(new_n500), .B1(new_n770), .B2(new_n816), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n811), .A2(new_n812), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G150), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n777), .A2(new_n819), .B1(new_n775), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT93), .ZN(new_n822));
  INV_X1    g0622(.A(G143), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n809), .A2(new_n823), .B1(new_n762), .B2(new_n771), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(KEYINPUT34), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G50), .A2(new_n791), .B1(new_n792), .B2(G132), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n783), .A2(G58), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n789), .A2(G68), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n827), .A2(new_n266), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n825), .B2(KEYINPUT34), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n818), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n749), .A2(new_n746), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n832), .A2(new_n758), .B1(G77), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n803), .B1(new_n808), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT95), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n665), .B1(new_n617), .B2(new_n627), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n805), .A2(new_n806), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n839), .A2(KEYINPUT94), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(KEYINPUT94), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n807), .B(new_n665), .C1(new_n617), .C2(new_n627), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n837), .B1(new_n844), .B2(new_n735), .ZN(new_n845));
  INV_X1    g0645(.A(new_n735), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n846), .A2(KEYINPUT95), .A3(new_n842), .A4(new_n843), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n845), .A2(new_n847), .B1(new_n735), .B2(new_n844), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n836), .B1(new_n848), .B2(new_n803), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT96), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT96), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n851), .B(new_n836), .C1(new_n848), .C2(new_n803), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n852), .ZN(G384));
  NOR2_X1   g0653(.A1(new_n742), .A2(new_n206), .ZN(new_n854));
  INV_X1    g0654(.A(G330), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n392), .A2(new_n294), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n364), .A2(KEYINPUT16), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n349), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n642), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n395), .B2(new_n404), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n400), .B1(new_n402), .B2(new_n859), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n393), .A2(new_n387), .A3(new_n349), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  INV_X1    g0666(.A(new_n864), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(new_n866), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n858), .B1(new_n402), .B2(new_n859), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n865), .A2(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n862), .A2(new_n870), .A3(KEYINPUT38), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n398), .A2(new_n642), .B1(new_n393), .B2(new_n349), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n872), .B2(KEYINPUT98), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n865), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n863), .A2(KEYINPUT98), .A3(KEYINPUT37), .A4(new_n864), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n369), .A2(new_n642), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT99), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n388), .B2(new_n394), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n369), .A2(new_n347), .A3(new_n387), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n864), .A2(KEYINPUT17), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT99), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n879), .A2(new_n632), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n876), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n871), .B1(new_n884), .B2(KEYINPUT38), .ZN(new_n885));
  OAI211_X1 g0685(.A(KEYINPUT31), .B(new_n644), .C1(new_n720), .C2(new_n727), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n704), .B(new_n886), .C1(new_n733), .C2(new_n706), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n314), .A2(new_n645), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n287), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT72), .B1(new_n281), .B2(new_n282), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n890), .A2(new_n285), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n319), .B(new_n889), .C1(new_n892), .C2(new_n314), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n291), .A2(new_n888), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n839), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n887), .A2(KEYINPUT40), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n880), .A2(new_n881), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n860), .B1(new_n632), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n869), .A2(KEYINPUT37), .A3(new_n864), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n866), .B1(new_n872), .B2(new_n867), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n862), .B2(new_n870), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n887), .B(new_n895), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n885), .A2(new_n896), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n438), .A2(new_n887), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n855), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT100), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n912), .B(new_n913), .C1(new_n908), .C2(new_n909), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n893), .A2(new_n894), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n843), .B2(new_n806), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n899), .B1(new_n898), .B2(new_n902), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n871), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n404), .A2(new_n642), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n316), .A2(new_n644), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n917), .B2(new_n871), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n924), .B(new_n871), .C1(new_n884), .C2(KEYINPUT38), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n438), .A2(new_n701), .A3(new_n692), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n637), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n854), .B1(new_n914), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n914), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n675), .A2(new_n410), .A3(new_n353), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(G68), .B2(new_n201), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n936), .A2(new_n206), .A3(G13), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT97), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT36), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n226), .A2(G20), .A3(G116), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n474), .B2(KEYINPUT35), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(KEYINPUT35), .B2(new_n474), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n938), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n939), .B2(new_n942), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n934), .A2(new_n944), .ZN(G367));
  AND2_X1   g0745(.A1(new_n622), .A2(new_n625), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n666), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n666), .A2(new_n622), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n947), .B1(new_n679), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n615), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n666), .B1(new_n951), .B2(new_n533), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n607), .A2(KEYINPUT84), .A3(new_n644), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n662), .B1(new_n650), .B2(new_n645), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n658), .B(new_n950), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT42), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(KEYINPUT42), .B1(new_n664), .B2(new_n950), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT102), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT43), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n956), .A2(new_n957), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n664), .A2(KEYINPUT42), .A3(new_n950), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n952), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT43), .B1(new_n966), .B2(KEYINPUT102), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n529), .B(KEYINPUT101), .C1(new_n509), .C2(new_n645), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT101), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n509), .A2(new_n645), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n620), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n528), .A3(new_n526), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n968), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n963), .A2(new_n967), .A3(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n963), .A2(new_n967), .B1(new_n973), .B2(new_n960), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT103), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT103), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n963), .A2(new_n967), .A3(new_n973), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n963), .A2(new_n967), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n960), .A2(new_n973), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n977), .B(new_n978), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n950), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n659), .A2(new_n982), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n976), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n983), .B1(new_n976), .B2(new_n981), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n743), .A2(G1), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n855), .B(new_n660), .C1(new_n646), .C2(new_n652), .ZN(new_n987));
  AOI21_X1  g0787(.A(KEYINPUT45), .B1(new_n668), .B2(new_n950), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT45), .ZN(new_n989));
  NOR4_X1   g0789(.A1(new_n664), .A2(new_n982), .A3(new_n989), .A4(new_n667), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT44), .B1(new_n668), .B2(new_n950), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT44), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n993), .B(new_n982), .C1(new_n664), .C2(new_n667), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n987), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n661), .A2(new_n663), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n658), .ZN(new_n998));
  INV_X1    g0798(.A(new_n667), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n998), .A2(new_n999), .A3(new_n950), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n989), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n668), .A2(KEYINPUT45), .A3(new_n950), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1003), .A2(new_n659), .A3(new_n992), .A4(new_n994), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n658), .B1(new_n653), .B2(G330), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n663), .B(new_n661), .C1(new_n1005), .C2(new_n987), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n741), .A2(new_n660), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1007), .A2(new_n659), .A3(new_n997), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n996), .A2(new_n1004), .A3(new_n737), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n737), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n671), .B(KEYINPUT41), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n986), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n984), .A2(new_n985), .A3(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n780), .A2(new_n516), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1015), .A2(KEYINPUT46), .B1(G107), .B2(new_n783), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(KEYINPUT46), .B2(new_n1015), .C1(new_n816), .C2(new_n775), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G97), .A2(new_n789), .B1(new_n761), .B2(G283), .ZN(new_n1018));
  INV_X1    g0818(.A(G317), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n770), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n275), .B1(new_n810), .B2(new_n777), .C1(new_n809), .C2(new_n814), .ZN(new_n1021));
  NOR3_X1   g0821(.A1(new_n1017), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT104), .Z(new_n1023));
  NOR2_X1   g0823(.A1(new_n782), .A2(new_n303), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n275), .B(new_n1024), .C1(G150), .C2(new_n767), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n201), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n761), .A2(new_n1026), .B1(new_n791), .B2(G58), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n764), .A2(new_n410), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G137), .B2(new_n792), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G143), .A2(new_n776), .B1(new_n778), .B2(G159), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1025), .A2(new_n1027), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1023), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT47), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n749), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n973), .A2(new_n799), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n751), .B1(new_n670), .B2(new_n413), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n752), .A2(new_n237), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n744), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1034), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT105), .B1(new_n1014), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n985), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1013), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n976), .A2(new_n981), .A3(new_n983), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT105), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n1046), .A3(new_n1039), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1041), .A2(new_n1047), .ZN(G387));
  OAI21_X1  g0848(.A(new_n275), .B1(new_n770), .B2(new_n786), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n780), .A2(new_n810), .B1(new_n782), .B2(new_n813), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G317), .A2(new_n767), .B1(new_n761), .B2(G303), .ZN(new_n1051));
  XOR2_X1   g0851(.A(KEYINPUT107), .B(G322), .Z(new_n1052));
  OAI221_X1 g0852(.A(new_n1051), .B1(new_n816), .B2(new_n777), .C1(new_n775), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT48), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n1054), .B2(new_n1053), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT49), .Z(new_n1057));
  AOI211_X1 g0857(.A(new_n1049), .B(new_n1057), .C1(G116), .C2(new_n789), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n809), .A2(new_n214), .B1(new_n762), .B2(new_n303), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n791), .A2(G77), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n819), .B2(new_n770), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n266), .B1(new_n764), .B2(new_n216), .C1(new_n777), .C2(new_n332), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n505), .A2(new_n782), .B1(new_n771), .B2(new_n775), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n749), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT106), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n333), .A2(new_n214), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT50), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n673), .B(new_n510), .C1(new_n303), .C2(new_n410), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n752), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1066), .A2(new_n1070), .B1(new_n234), .B2(G45), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n755), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1072), .B1(G107), .B2(new_n210), .C1(new_n673), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n751), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n744), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1065), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(KEYINPUT108), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n660), .B2(new_n748), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(KEYINPUT108), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1079), .A2(new_n1080), .B1(new_n986), .B2(new_n1009), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT109), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n1009), .B2(new_n737), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1009), .A2(new_n737), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n736), .A3(KEYINPUT109), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1083), .A2(new_n671), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1081), .A2(new_n1087), .ZN(G393));
  NAND2_X1  g0888(.A1(new_n996), .A2(new_n1004), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n986), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n982), .A2(new_n748), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1075), .B1(new_n216), .B2(new_n210), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n244), .A2(new_n670), .A3(new_n266), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n803), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n809), .A2(new_n771), .B1(new_n819), .B2(new_n775), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT51), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n782), .A2(new_n410), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n266), .B1(new_n764), .B2(new_n500), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(new_n1026), .C2(new_n778), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n762), .A2(new_n332), .B1(new_n770), .B2(new_n823), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G68), .B2(new_n791), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1097), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT110), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n776), .A2(G317), .B1(new_n767), .B2(G311), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT52), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1052), .A2(new_n770), .B1(new_n780), .B2(new_n813), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT111), .Z(new_n1109));
  OAI221_X1 g0909(.A(new_n275), .B1(new_n418), .B2(new_n764), .C1(new_n762), .C2(new_n810), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n777), .A2(new_n814), .B1(new_n782), .B2(new_n516), .ZN(new_n1111));
  OR4_X1    g0911(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1105), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1095), .B1(new_n1114), .B2(new_n749), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1091), .B1(new_n1092), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1089), .A2(new_n1084), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n671), .A3(new_n1010), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(G390));
  OAI21_X1  g0919(.A(KEYINPUT112), .B1(new_n916), .B2(new_n922), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n883), .A2(new_n877), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n874), .A2(new_n875), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n903), .B1(new_n1123), .B2(new_n899), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n925), .B1(new_n1124), .B2(new_n924), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT112), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n700), .A2(new_n807), .B1(new_n634), .B2(new_n645), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1126), .B(new_n923), .C1(new_n1127), .C2(new_n915), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1120), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n645), .B(new_n805), .C1(new_n684), .C2(new_n691), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n806), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n915), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1124), .A2(new_n922), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n704), .A2(new_n728), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n733), .A2(KEYINPUT31), .ZN(new_n1137));
  OAI211_X1 g0937(.A(G330), .B(new_n807), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1138), .A2(new_n915), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1129), .A2(new_n1135), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n887), .A2(G330), .A3(new_n895), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT113), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n887), .A2(new_n895), .A3(KEYINPUT113), .A4(G330), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1129), .A2(new_n1135), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n438), .A2(G330), .A3(new_n887), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n930), .A2(new_n1147), .A3(new_n637), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1138), .A2(new_n915), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1143), .A2(new_n1149), .A3(new_n1144), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1127), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n840), .A2(new_n841), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n887), .A2(G330), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n915), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1139), .A2(new_n1155), .A3(new_n806), .A4(new_n1130), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1148), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n672), .B1(new_n1146), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1148), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1161), .B(KEYINPUT114), .C1(new_n1140), .C2(new_n1145), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1129), .A2(new_n1135), .A3(new_n1139), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT114), .B1(new_n1168), .B2(new_n1161), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1158), .B1(new_n1163), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT115), .B1(new_n1168), .B2(new_n1090), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT115), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1146), .A2(new_n1172), .A3(new_n986), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1125), .A2(new_n746), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n762), .A2(new_n216), .B1(new_n813), .B2(new_n775), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G107), .B2(new_n778), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT117), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n829), .B1(new_n810), .B2(new_n770), .C1(new_n809), .C2(new_n516), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n1178), .A2(new_n266), .A3(new_n781), .A4(new_n1098), .ZN(new_n1179));
  INV_X1    g0979(.A(G125), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n266), .B1(new_n770), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(G128), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n777), .A2(new_n820), .B1(new_n775), .B2(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1181), .B(new_n1183), .C1(G159), .C2(new_n783), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT54), .B(G143), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1026), .A2(new_n789), .B1(new_n761), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(G132), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n809), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT53), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n780), .B2(new_n819), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n791), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1189), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1177), .A2(new_n1179), .B1(new_n1184), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(new_n758), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n744), .B1(new_n332), .B2(new_n833), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(KEYINPUT116), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1196), .A2(KEYINPUT116), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1171), .A2(new_n1173), .B1(new_n1174), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1170), .A2(new_n1200), .ZN(G378));
  AOI21_X1  g1001(.A(new_n744), .B1(new_n201), .B2(new_n833), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n775), .A2(new_n1180), .B1(new_n782), .B2(new_n819), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n791), .A2(new_n1186), .B1(new_n767), .B2(G128), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n820), .B2(new_n762), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(G132), .C2(new_n778), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n789), .A2(G159), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n792), .C2(G124), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT59), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(new_n1213), .B2(new_n1207), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1024), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n266), .A2(G41), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1060), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n809), .A2(new_n418), .B1(new_n764), .B2(new_n352), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n762), .A2(new_n505), .B1(new_n770), .B2(new_n813), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n777), .A2(new_n216), .B1(new_n775), .B2(new_n516), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(KEYINPUT58), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(KEYINPUT58), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1222), .B(new_n1223), .C1(new_n1216), .C2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n749), .B1(new_n1214), .B2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT118), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n642), .B1(new_n339), .B2(new_n342), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT119), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n346), .A2(new_n408), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1232), .B1(new_n346), .B2(new_n408), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1230), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1235), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(new_n1229), .A3(new_n1233), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1203), .B(new_n1227), .C1(new_n746), .C2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n921), .A2(new_n928), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(KEYINPUT120), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n896), .A2(new_n885), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n905), .A2(new_n906), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(G330), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1239), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n907), .A2(G330), .A3(new_n1239), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT121), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1243), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1239), .B1(new_n907), .B2(G330), .ZN(new_n1254));
  AND4_X1   g1054(.A1(G330), .A2(new_n1244), .A3(new_n1245), .A4(new_n1239), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT121), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n1242), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1253), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1240), .B1(new_n1259), .B2(new_n986), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1166), .A2(new_n1167), .A3(new_n1157), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1160), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT57), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n929), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1248), .A2(new_n1249), .A3(new_n1241), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1264), .A2(KEYINPUT57), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n671), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1260), .B1(new_n1263), .B2(new_n1268), .ZN(G375));
  OAI22_X1  g1069(.A1(new_n809), .A2(new_n820), .B1(new_n762), .B2(new_n819), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n780), .A2(new_n771), .B1(new_n770), .B2(new_n1182), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n266), .B1(new_n764), .B2(new_n352), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n775), .A2(new_n1188), .B1(new_n782), .B2(new_n214), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1273), .B(new_n1274), .C1(new_n778), .C2(new_n1186), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n777), .A2(new_n516), .B1(new_n775), .B2(new_n810), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n505), .A2(new_n782), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(new_n1276), .A2(new_n1277), .A3(new_n266), .A4(new_n1028), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n809), .A2(new_n813), .B1(new_n762), .B2(new_n418), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n780), .A2(new_n216), .B1(new_n770), .B2(new_n814), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1272), .A2(new_n1275), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1282));
  OAI221_X1 g1082(.A(new_n803), .B1(G68), .B2(new_n834), .C1(new_n1282), .C2(new_n758), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(new_n915), .B2(new_n746), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(new_n1159), .B2(new_n986), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(KEYINPUT122), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1152), .A2(new_n1156), .A3(new_n1148), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1161), .A2(new_n1012), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(G381));
  NAND3_X1  g1089(.A1(new_n1081), .A2(new_n801), .A3(new_n1087), .ZN(new_n1290));
  OR4_X1    g1090(.A1(G384), .A2(G381), .A3(G390), .A4(new_n1290), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(G387), .A2(new_n1291), .A3(G378), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G375), .A2(KEYINPUT123), .ZN(new_n1293));
  OR2_X1    g1093(.A1(G375), .A2(KEYINPUT123), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .ZN(G407));
  NAND2_X1  g1095(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1174), .A2(new_n1199), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1261), .A2(new_n671), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT114), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1146), .B2(new_n1157), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1299), .B1(new_n1301), .B2(new_n1162), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1298), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n643), .A2(G213), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1294), .A2(new_n1303), .A3(new_n1293), .A4(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(G407), .A2(G213), .A3(new_n1306), .ZN(G409));
  AND3_X1   g1107(.A1(new_n1256), .A2(new_n1242), .A3(new_n1257), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1242), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1262), .B(new_n1012), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1240), .B1(new_n1311), .B2(new_n986), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(new_n1170), .A3(new_n1200), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(G375), .B2(new_n1303), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT124), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G384), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n850), .A2(KEYINPUT124), .A3(new_n852), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT60), .ZN(new_n1319));
  OR2_X1    g1119(.A1(new_n1287), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1287), .A2(new_n1319), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1320), .A2(new_n671), .A3(new_n1161), .A4(new_n1321), .ZN(new_n1322));
  AOI22_X1  g1122(.A1(new_n1317), .A2(new_n1318), .B1(new_n1286), .B2(new_n1322), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1286), .A2(new_n1322), .A3(new_n1318), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1315), .A2(new_n1304), .A3(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1290), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n801), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1045), .A2(new_n1039), .ZN(new_n1331));
  INV_X1    g1131(.A(G390), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n985), .A2(new_n1013), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1040), .B1(new_n1334), .B2(new_n1044), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1335), .A2(G390), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1330), .B1(new_n1333), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT125), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(G390), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT125), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1041), .A2(new_n1047), .A3(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1330), .B1(new_n1335), .B2(G390), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  AOI22_X1  g1144(.A1(new_n1326), .A2(new_n1327), .B1(new_n1337), .B2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1315), .A2(new_n1304), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1286), .A2(new_n1322), .A3(new_n1318), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1305), .A2(G2897), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1349));
  AND2_X1   g1149(.A1(new_n1286), .A2(new_n1322), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n1347), .B(new_n1348), .C1(new_n1349), .C2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1348), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1352), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1353));
  AND2_X1   g1153(.A1(new_n1351), .A2(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(KEYINPUT61), .B1(new_n1346), .B2(new_n1354), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1315), .A2(KEYINPUT63), .A3(new_n1304), .A4(new_n1325), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(KEYINPUT126), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n672), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1358));
  AOI22_X1  g1158(.A1(new_n1253), .A2(new_n1258), .B1(new_n1160), .B2(new_n1261), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1358), .B1(new_n1359), .B2(KEYINPUT57), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(G378), .A2(new_n1360), .A3(new_n1260), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1305), .B1(new_n1361), .B2(new_n1314), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT126), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1362), .A2(new_n1363), .A3(KEYINPUT63), .A4(new_n1325), .ZN(new_n1364));
  NAND4_X1  g1164(.A1(new_n1345), .A2(new_n1355), .A3(new_n1357), .A4(new_n1364), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(new_n1326), .A2(KEYINPUT62), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT61), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1351), .A2(new_n1353), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1367), .B1(new_n1362), .B2(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT62), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1370), .B1(new_n1362), .B2(new_n1325), .ZN(new_n1371));
  NOR3_X1   g1171(.A1(new_n1366), .A2(new_n1369), .A3(new_n1371), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1344), .A2(new_n1337), .ZN(new_n1373));
  INV_X1    g1173(.A(KEYINPUT127), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1373), .A2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1335), .A2(G390), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1376), .A2(new_n1377), .ZN(new_n1378));
  AOI22_X1  g1178(.A1(new_n1378), .A2(new_n1330), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1379), .A2(KEYINPUT127), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1375), .A2(new_n1380), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1365), .B1(new_n1372), .B2(new_n1381), .ZN(G405));
  NAND2_X1  g1182(.A1(G375), .A2(new_n1303), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1383), .A2(new_n1361), .ZN(new_n1384));
  XNOR2_X1  g1184(.A(new_n1384), .B(new_n1325), .ZN(new_n1385));
  XNOR2_X1  g1185(.A(new_n1385), .B(new_n1379), .ZN(G402));
endmodule


