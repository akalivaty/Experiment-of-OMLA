//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n456), .A2(new_n457), .B1(new_n458), .B2(new_n452), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n457), .B2(new_n456), .ZN(G319));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  INV_X1    g045(.A(new_n465), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI211_X1 g047(.A(G137), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n463), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  AOI21_X1  g050(.A(KEYINPUT68), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n473), .A2(KEYINPUT68), .A3(new_n475), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n469), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT69), .ZN(G160));
  AOI21_X1  g055(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n470), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n464), .A2(new_n465), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI221_X1 g062(.A(new_n482), .B1(new_n483), .B2(new_n484), .C1(new_n485), .C2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT70), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT72), .A2(G138), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n481), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n470), .B(new_n491), .C1(new_n471), .C2(new_n472), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G126), .B(G2105), .C1(new_n471), .C2(new_n472), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT71), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n496), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n495), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n512), .B(G62), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(G651), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n509), .A2(new_n510), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(G88), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n521), .A2(G50), .A3(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n525), .B1(new_n523), .B2(new_n524), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n518), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n518), .B(KEYINPUT75), .C1(new_n526), .C2(new_n527), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(G166));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT76), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT7), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n508), .B1(new_n519), .B2(new_n520), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G51), .ZN(new_n538));
  AND2_X1   g113(.A1(G63), .A2(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n522), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n521), .A2(new_n522), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n538), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n536), .A2(new_n543), .ZN(G168));
  NAND2_X1  g119(.A1(new_n537), .A2(G52), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n546), .B2(new_n542), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G651), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(G171));
  NAND2_X1  g126(.A1(new_n537), .A2(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n542), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT77), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n549), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(new_n537), .A2(G53), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n521), .A2(new_n522), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n514), .A2(new_n515), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(G91), .A2(new_n566), .B1(new_n570), .B2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n565), .A2(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  XNOR2_X1  g148(.A(new_n534), .B(KEYINPUT7), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n566), .A2(G89), .B1(new_n522), .B2(new_n539), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n574), .A2(new_n538), .A3(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G168), .A2(KEYINPUT78), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(G286));
  INV_X1    g155(.A(G166), .ZN(G303));
  NAND2_X1  g156(.A1(new_n537), .A2(G49), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n521), .A2(new_n522), .A3(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT79), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n566), .A2(G87), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n587), .A2(new_n588), .A3(new_n583), .A4(new_n582), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(new_n522), .A2(G61), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n549), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n521), .A2(new_n522), .A3(G86), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n521), .A2(G48), .A3(G543), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G60), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n568), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(KEYINPUT82), .B(G85), .Z(new_n608));
  AOI22_X1  g183(.A1(new_n566), .A2(new_n608), .B1(G47), .B2(new_n537), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n605), .A2(new_n606), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(G290));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NOR2_X1   g188(.A1(G301), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n616));
  OR3_X1    g191(.A1(new_n542), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n568), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n620), .A2(G651), .B1(G54), .B2(new_n537), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n616), .B1(new_n542), .B2(new_n615), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT84), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n614), .B1(new_n625), .B2(new_n613), .ZN(G284));
  AOI21_X1  g201(.A(new_n614), .B1(new_n625), .B2(new_n613), .ZN(G321));
  NOR2_X1   g202(.A1(G299), .A2(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n578), .A2(new_n579), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G297));
  AOI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G280));
  NOR2_X1   g206(.A1(new_n624), .A2(G559), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(G860), .B2(new_n625), .ZN(G148));
  OAI21_X1  g208(.A(new_n613), .B1(new_n555), .B2(new_n557), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n632), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n486), .A2(new_n474), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT85), .B(KEYINPUT12), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n640), .A2(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT86), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n481), .A2(G135), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n470), .A2(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  INV_X1    g220(.A(G123), .ZN(new_n646));
  OAI221_X1 g221(.A(new_n643), .B1(new_n644), .B2(new_n645), .C1(new_n646), .C2(new_n487), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2096), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n640), .B2(G2100), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n642), .A2(new_n649), .ZN(G156));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n654), .B2(new_n653), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(G401));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n666), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT87), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2096), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT18), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n667), .A2(new_n668), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT88), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n673), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n685), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n687), .B(new_n689), .C1(new_n682), .C2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(KEYINPUT34), .ZN(new_n698));
  NOR2_X1   g273(.A1(G16), .A2(G22), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G166), .B2(G16), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1971), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n600), .A2(G16), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G6), .B2(G16), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT32), .B(G1981), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT91), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n702), .B(new_n705), .C1(G6), .C2(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n701), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT92), .B1(new_n584), .B2(new_n585), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT92), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n587), .A2(new_n713), .A3(new_n583), .A4(new_n582), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n711), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n711), .A2(G23), .ZN(new_n716));
  OR3_X1    g291(.A1(new_n715), .A2(KEYINPUT93), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(KEYINPUT93), .B1(new_n715), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT33), .B(G1976), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n710), .A2(KEYINPUT94), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(KEYINPUT94), .B1(new_n710), .B2(new_n721), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n698), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G1971), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n700), .B(new_n726), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n721), .A2(new_n727), .A3(new_n708), .A4(new_n707), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT94), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n730), .A2(KEYINPUT34), .A3(new_n722), .ZN(new_n731));
  MUX2_X1   g306(.A(G24), .B(G290), .S(G16), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1986), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n481), .A2(G131), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n470), .A2(G107), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n736));
  INV_X1    g311(.A(G119), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n734), .B1(new_n735), .B2(new_n736), .C1(new_n737), .C2(new_n487), .ZN(new_n738));
  MUX2_X1   g313(.A(G25), .B(new_n738), .S(G29), .Z(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT90), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n739), .B(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n733), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n725), .A2(new_n731), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(KEYINPUT95), .A2(KEYINPUT36), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n725), .A2(new_n745), .A3(new_n731), .A4(new_n743), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G29), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G32), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n470), .A2(G105), .A3(G2104), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT98), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G141), .ZN(new_n755));
  INV_X1    g330(.A(new_n481), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(KEYINPUT26), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(KEYINPUT26), .ZN(new_n760));
  INV_X1    g335(.A(G129), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n759), .B(new_n760), .C1(new_n487), .C2(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n751), .B1(new_n764), .B2(new_n750), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT27), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1996), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n750), .A2(G27), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n750), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(G2078), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n750), .A2(G33), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n486), .A2(G127), .ZN(new_n772));
  INV_X1    g347(.A(G115), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n463), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT97), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n470), .B1(new_n774), .B2(KEYINPUT97), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT25), .Z(new_n779));
  INV_X1    g354(.A(G139), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n756), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n771), .B1(new_n782), .B2(new_n750), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(G2072), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G2078), .B2(new_n769), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n711), .A2(G5), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G171), .B2(new_n711), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(G1961), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n783), .B2(G2072), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n767), .A2(new_n770), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n711), .A2(G21), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G168), .B2(new_n711), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G1966), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(G1966), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT30), .B(G28), .ZN(new_n795));
  OR2_X1    g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  NAND2_X1  g371(.A1(KEYINPUT31), .A2(G11), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n795), .A2(new_n750), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n647), .B2(new_n750), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n787), .B2(G1961), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n793), .A2(new_n794), .A3(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  INV_X1    g377(.A(G34), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n803), .A2(KEYINPUT24), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(KEYINPUT24), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n750), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G160), .B2(new_n750), .ZN(new_n807));
  INV_X1    g382(.A(G2084), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n802), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n790), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT100), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT100), .B1(new_n790), .B2(new_n810), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n750), .A2(G35), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G162), .B2(new_n750), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT29), .B(G2090), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT101), .B(KEYINPUT23), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n711), .A2(G20), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G299), .B2(G16), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1956), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n481), .A2(G140), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n470), .A2(G116), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n826));
  INV_X1    g401(.A(G128), .ZN(new_n827));
  OAI221_X1 g402(.A(new_n824), .B1(new_n825), .B2(new_n826), .C1(new_n827), .C2(new_n487), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G29), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n750), .A2(G26), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT28), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G2067), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n818), .A2(new_n823), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(G4), .A2(G16), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n625), .B2(G16), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT96), .B(G1348), .Z(new_n838));
  AND2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n711), .A2(G19), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n558), .B2(new_n711), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G1341), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n837), .A2(new_n838), .ZN(new_n843));
  NOR4_X1   g418(.A1(new_n835), .A2(new_n839), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n813), .A2(new_n814), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT102), .B1(new_n749), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n848));
  AOI211_X1 g423(.A(new_n848), .B(new_n845), .C1(new_n747), .C2(new_n748), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n847), .A2(new_n849), .ZN(G311));
  NAND2_X1  g425(.A1(new_n749), .A2(new_n846), .ZN(G150));
  NAND2_X1  g426(.A1(new_n625), .A2(G559), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT38), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n537), .A2(G55), .ZN(new_n854));
  INV_X1    g429(.A(G93), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(new_n542), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(new_n549), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n558), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n853), .B(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  INV_X1    g437(.A(G860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n859), .A2(new_n863), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(G145));
  XNOR2_X1  g443(.A(G160), .B(new_n647), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G162), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n763), .B(new_n828), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n639), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n481), .A2(G142), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n470), .A2(G118), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  INV_X1    g450(.A(G130), .ZN(new_n876));
  OAI221_X1 g451(.A(new_n873), .B1(new_n874), .B2(new_n875), .C1(new_n876), .C2(new_n487), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n738), .B(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n872), .B(new_n878), .Z(new_n879));
  INV_X1    g454(.A(new_n499), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n495), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n872), .B(new_n878), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n499), .B1(new_n494), .B2(new_n492), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n782), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n782), .B1(new_n882), .B2(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n870), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  INV_X1    g465(.A(new_n870), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n891), .A3(new_n886), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(KEYINPUT103), .B(KEYINPUT40), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(G395));
  NAND2_X1  g471(.A1(new_n712), .A2(new_n714), .ZN(new_n897));
  XNOR2_X1  g472(.A(G166), .B(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n600), .B(G290), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n901), .A2(KEYINPUT42), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(KEYINPUT42), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n860), .B(new_n632), .ZN(new_n906));
  XOR2_X1   g481(.A(G299), .B(new_n623), .Z(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT41), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n907), .B2(new_n906), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n905), .A2(new_n910), .ZN(new_n912));
  OAI21_X1  g487(.A(G868), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n859), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n613), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(G295));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n913), .A2(new_n917), .A3(new_n915), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n913), .B2(new_n915), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(G331));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n921));
  NAND3_X1  g496(.A1(G286), .A2(new_n921), .A3(G171), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n576), .B2(G171), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n629), .B2(G301), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n558), .B(new_n914), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n860), .A2(new_n922), .A3(new_n924), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n928), .A3(new_n907), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n908), .B1(new_n927), .B2(new_n928), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n932), .B2(new_n900), .ZN(new_n933));
  INV_X1    g508(.A(new_n900), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n930), .B2(new_n931), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n933), .A2(KEYINPUT43), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT107), .B1(new_n930), .B2(new_n931), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n927), .A2(new_n928), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n938), .B(new_n929), .C1(new_n939), .C2(new_n908), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n940), .A3(new_n934), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT43), .B1(new_n941), .B2(new_n933), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT44), .B1(new_n936), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(new_n941), .B2(new_n933), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n933), .A2(new_n944), .A3(new_n935), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n945), .B2(new_n946), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n943), .B1(new_n950), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g526(.A(new_n478), .ZN(new_n952));
  OAI211_X1 g527(.A(G40), .B(new_n468), .C1(new_n952), .C2(new_n476), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n881), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT109), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n955), .B1(new_n884), .B2(G1384), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(new_n953), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n828), .A2(G2067), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n828), .A2(G2067), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n959), .B(new_n963), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1996), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n961), .A2(new_n967), .A3(new_n764), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n959), .A2(new_n963), .A3(G1996), .A4(new_n763), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n970), .A2(KEYINPUT110), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(KEYINPUT110), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n959), .A2(new_n963), .ZN(new_n974));
  INV_X1    g549(.A(new_n740), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n738), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(G290), .B(G1986), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n961), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT119), .ZN(new_n981));
  INV_X1    g556(.A(new_n598), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(G1981), .ZN(new_n983));
  INV_X1    g558(.A(G1981), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT116), .B1(new_n598), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G61), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n593), .B1(new_n568), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G651), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n988), .A2(new_n984), .A3(new_n595), .A4(new_n596), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n983), .B1(new_n985), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n989), .A2(new_n990), .ZN(new_n996));
  INV_X1    g571(.A(new_n597), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n997), .A2(KEYINPUT116), .A3(new_n984), .A4(new_n988), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n996), .A2(new_n998), .B1(new_n982), .B2(G1981), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT49), .B1(new_n999), .B2(KEYINPUT117), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n957), .A2(new_n953), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n995), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(new_n897), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n495), .B2(new_n880), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n954), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n712), .A2(new_n714), .A3(KEYINPUT115), .A4(G1976), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1007), .A2(new_n1009), .A3(G8), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT52), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1013), .A2(new_n1003), .A3(new_n1010), .A4(new_n1007), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1004), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n530), .A2(G8), .A3(new_n531), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(KEYINPUT112), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n1021));
  NAND4_X1  g596(.A1(new_n530), .A2(G8), .A3(new_n531), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT113), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1008), .A2(KEYINPUT45), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n954), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT45), .B1(new_n503), .B2(new_n956), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n726), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n503), .B2(new_n956), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n953), .B1(new_n1029), .B2(new_n1008), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT111), .B(G2090), .Z(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1002), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1020), .A2(new_n1036), .A3(new_n1022), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1024), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT114), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1024), .A2(new_n1037), .A3(new_n1040), .A4(new_n1035), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1027), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n953), .B1(KEYINPUT45), .B2(new_n1008), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1971), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n503), .A2(new_n1029), .A3(new_n956), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT50), .B1(new_n884), .B2(G1384), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1046), .A2(new_n954), .A3(new_n1047), .A4(new_n1033), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT118), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G8), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1045), .A2(new_n1049), .A3(KEYINPUT118), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1037), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1036), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1051), .A2(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n956), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n954), .A3(new_n960), .ZN(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1031), .A2(new_n1032), .A3(new_n808), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(G8), .A3(new_n629), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(KEYINPUT63), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1055), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1015), .B1(new_n1042), .B2(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n1002), .B(G286), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(new_n1004), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1035), .B1(new_n1024), .B2(new_n1037), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT63), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1003), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n995), .A2(new_n1000), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(new_n1006), .A3(new_n590), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n985), .A2(new_n991), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1071), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1070), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n981), .B1(new_n1065), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1015), .A2(new_n1062), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1035), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1076), .B1(new_n1083), .B2(KEYINPUT63), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1039), .A2(new_n1041), .B1(new_n1055), .B2(new_n1063), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1084), .B(KEYINPUT119), .C1(new_n1085), .C2(new_n1015), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1079), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1042), .A2(new_n1004), .A3(new_n1066), .A4(new_n1055), .ZN(new_n1088));
  INV_X1    g663(.A(G1348), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1008), .A2(new_n1029), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n954), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1089), .B1(new_n1091), .B2(new_n1030), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1001), .A2(new_n833), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n624), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n625), .A2(new_n1092), .A3(KEYINPUT60), .A4(new_n1093), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1026), .A2(new_n1027), .A3(G1996), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT58), .B(G1341), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1001), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n558), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT59), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1105), .B(new_n558), .C1(new_n1100), .C2(new_n1102), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n1108));
  XNOR2_X1  g683(.A(G299), .B(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1046), .A2(new_n954), .A3(new_n1047), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1043), .A2(new_n1044), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1109), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(new_n1114), .A3(new_n1109), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(KEYINPUT61), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1117), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(new_n1115), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1099), .A2(new_n1107), .A3(new_n1118), .A4(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n624), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1117), .B1(new_n1115), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G2078), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1043), .A2(new_n1044), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(KEYINPUT122), .B2(new_n1126), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(KEYINPUT122), .B2(new_n1126), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n957), .B2(new_n955), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n953), .A2(KEYINPUT121), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n953), .A2(KEYINPUT121), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1025), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G1961), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1091), .B2(new_n1030), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(G171), .B1(new_n1129), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1128), .A2(G2078), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1057), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1140), .A2(new_n1143), .A3(G301), .A4(new_n1137), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(KEYINPUT54), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT123), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1139), .A2(new_n1147), .A3(new_n1144), .A4(KEYINPUT54), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1059), .A2(new_n1060), .A3(G168), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1002), .B1(KEYINPUT120), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(KEYINPUT120), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1150), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1061), .A2(G8), .A3(new_n576), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1154), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1143), .A2(new_n1137), .ZN(new_n1160));
  OAI21_X1  g735(.A(G171), .B1(new_n1160), .B2(new_n1129), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1140), .A2(G301), .A3(new_n1137), .A4(new_n1135), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT54), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1125), .A2(new_n1149), .A3(new_n1164), .ZN(new_n1165));
  OR3_X1    g740(.A1(new_n1157), .A2(KEYINPUT62), .A3(new_n1158), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1161), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT62), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1088), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n980), .B1(new_n1087), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n978), .A2(KEYINPUT125), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n973), .A2(new_n1173), .A3(new_n977), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n958), .A2(G290), .A3(G1986), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT48), .Z(new_n1176));
  AND3_X1   g751(.A1(new_n1172), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n961), .A2(new_n967), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT46), .ZN(new_n1179));
  INV_X1    g754(.A(new_n974), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1179), .B(new_n966), .C1(new_n1180), .C2(new_n764), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT47), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n738), .A2(new_n975), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT124), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n965), .B1(new_n973), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1182), .B1(new_n1185), .B2(new_n1180), .ZN(new_n1186));
  OAI21_X1  g761(.A(KEYINPUT126), .B1(new_n1177), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1172), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1185), .A2(new_n1180), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1182), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1171), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1171), .A2(new_n1192), .A3(KEYINPUT127), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g772(.A(G319), .ZN(new_n1199));
  NOR4_X1   g773(.A1(G229), .A2(new_n1199), .A3(G401), .A4(G227), .ZN(new_n1200));
  OAI211_X1 g774(.A(new_n894), .B(new_n1200), .C1(new_n947), .C2(new_n949), .ZN(G225));
  INV_X1    g775(.A(G225), .ZN(G308));
endmodule


